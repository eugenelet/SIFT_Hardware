module Gaussian_Blur_3x3(
  clk,
  rst_n,
  buffer_data_0,
  buffer_data_1,
  buffer_data_2,
  current_col,
  blur_out
);

input                 clk;
input                 rst_n;
input         [5:0]   current_col;
input       [175:0]   buffer_data_0;
input       [175:0]   buffer_data_1;
input       [175:0]   buffer_data_2;
output reg  [127:0]   blur_out; // wire

always @(posedge clk) begin
  if (!rst_n) begin
    G_Kernel_3x3[0][31:0]  <= 32'h17BC5428; //18'b00_0101_1110_1111_0001;//'d092717;
    G_Kernel_3x3[0][63:32] <= 32'h1E7ABFF3; //18'b00_0111_1001_1110_1010;//'d119061;
    G_Kernel_3x3[0][95:64] <= 32'h17BC5428; //18'b00_0101_1110_1111_0001;//'d092717;
    G_Kernel_3x3[1][31:0]  <= 32'h1E7ABFF3; //18'b00_0111_1001_1110_1010;//'d119061;
    G_Kernel_3x3[1][63:32] <= 32'h2723AF8E; //18'b00_1001_1100_1000_1110;//'d152888;
    G_Kernel_3x3[1][95:64] <= 32'h1E7ABFF3; //18'b00_0111_1001_1110_1011;//'d119061;
  end
end

reg    [23:0]    layer0[0:15]; //wire
reg    [23:0]    layer1[0:15]; //wire
reg    [23:0]    layer2[0:15]; //wire
always @(*) begin
  case(current_col)
    'd0: begin
        layer0[0][7:0] = 0;
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = 0;
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = 0;
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd1: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd2: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd3: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd4: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd5: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd6: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd7: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd8: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd9: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd10: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd11: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd12: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd13: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd14: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd15: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd16: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd17: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd18: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd19: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd20: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd21: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd22: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd23: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd24: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd25: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd26: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd27: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd28: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd29: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd30: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd31: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd32: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd33: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd34: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd35: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd36: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd37: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd38: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = buffer_data_2[159:152];
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = buffer_data_1[159:152];
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = buffer_data_0[159:152];
    end
    'd39: begin
        layer0[0][7:0] = buffer_data_2[23:16];
        layer0[0][15:8] = buffer_data_2[31:24];
        layer0[0][23:16] = buffer_data_2[39:32];
        layer1[0][7:0] = buffer_data_1[23:16];
        layer1[0][15:8] = buffer_data_1[31:24];
        layer1[0][23:16] = buffer_data_1[39:32];
        layer2[0][7:0] = buffer_data_0[23:16];
        layer2[0][15:8] = buffer_data_0[31:24];
        layer2[0][23:16] = buffer_data_0[39:32];
        layer0[1][7:0] = buffer_data_2[31:24];
        layer0[1][15:8] = buffer_data_2[39:32];
        layer0[1][23:16] = buffer_data_2[47:40];
        layer1[1][7:0] = buffer_data_1[31:24];
        layer1[1][15:8] = buffer_data_1[39:32];
        layer1[1][23:16] = buffer_data_1[47:40];
        layer2[1][7:0] = buffer_data_0[31:24];
        layer2[1][15:8] = buffer_data_0[39:32];
        layer2[1][23:16] = buffer_data_0[47:40];
        layer0[2][7:0] = buffer_data_2[39:32];
        layer0[2][15:8] = buffer_data_2[47:40];
        layer0[2][23:16] = buffer_data_2[55:48];
        layer1[2][7:0] = buffer_data_1[39:32];
        layer1[2][15:8] = buffer_data_1[47:40];
        layer1[2][23:16] = buffer_data_1[55:48];
        layer2[2][7:0] = buffer_data_0[39:32];
        layer2[2][15:8] = buffer_data_0[47:40];
        layer2[2][23:16] = buffer_data_0[55:48];
        layer0[3][7:0] = buffer_data_2[47:40];
        layer0[3][15:8] = buffer_data_2[55:48];
        layer0[3][23:16] = buffer_data_2[63:56];
        layer1[3][7:0] = buffer_data_1[47:40];
        layer1[3][15:8] = buffer_data_1[55:48];
        layer1[3][23:16] = buffer_data_1[63:56];
        layer2[3][7:0] = buffer_data_0[47:40];
        layer2[3][15:8] = buffer_data_0[55:48];
        layer2[3][23:16] = buffer_data_0[63:56];
        layer0[4][7:0] = buffer_data_2[55:48];
        layer0[4][15:8] = buffer_data_2[63:56];
        layer0[4][23:16] = buffer_data_2[71:64];
        layer1[4][7:0] = buffer_data_1[55:48];
        layer1[4][15:8] = buffer_data_1[63:56];
        layer1[4][23:16] = buffer_data_1[71:64];
        layer2[4][7:0] = buffer_data_0[55:48];
        layer2[4][15:8] = buffer_data_0[63:56];
        layer2[4][23:16] = buffer_data_0[71:64];
        layer0[5][7:0] = buffer_data_2[63:56];
        layer0[5][15:8] = buffer_data_2[71:64];
        layer0[5][23:16] = buffer_data_2[79:72];
        layer1[5][7:0] = buffer_data_1[63:56];
        layer1[5][15:8] = buffer_data_1[71:64];
        layer1[5][23:16] = buffer_data_1[79:72];
        layer2[5][7:0] = buffer_data_0[63:56];
        layer2[5][15:8] = buffer_data_0[71:64];
        layer2[5][23:16] = buffer_data_0[79:72];
        layer0[6][7:0] = buffer_data_2[71:64];
        layer0[6][15:8] = buffer_data_2[79:72];
        layer0[6][23:16] = buffer_data_2[87:80];
        layer1[6][7:0] = buffer_data_1[71:64];
        layer1[6][15:8] = buffer_data_1[79:72];
        layer1[6][23:16] = buffer_data_1[87:80];
        layer2[6][7:0] = buffer_data_0[71:64];
        layer2[6][15:8] = buffer_data_0[79:72];
        layer2[6][23:16] = buffer_data_0[87:80];
        layer0[7][7:0] = buffer_data_2[79:72];
        layer0[7][15:8] = buffer_data_2[87:80];
        layer0[7][23:16] = buffer_data_2[95:88];
        layer1[7][7:0] = buffer_data_1[79:72];
        layer1[7][15:8] = buffer_data_1[87:80];
        layer1[7][23:16] = buffer_data_1[95:88];
        layer2[7][7:0] = buffer_data_0[79:72];
        layer2[7][15:8] = buffer_data_0[87:80];
        layer2[7][23:16] = buffer_data_0[95:88];
        layer0[8][7:0] = buffer_data_2[87:80];
        layer0[8][15:8] = buffer_data_2[95:88];
        layer0[8][23:16] = buffer_data_2[103:96];
        layer1[8][7:0] = buffer_data_1[87:80];
        layer1[8][15:8] = buffer_data_1[95:88];
        layer1[8][23:16] = buffer_data_1[103:96];
        layer2[8][7:0] = buffer_data_0[87:80];
        layer2[8][15:8] = buffer_data_0[95:88];
        layer2[8][23:16] = buffer_data_0[103:96];
        layer0[9][7:0] = buffer_data_2[95:88];
        layer0[9][15:8] = buffer_data_2[103:96];
        layer0[9][23:16] = buffer_data_2[111:104];
        layer1[9][7:0] = buffer_data_1[95:88];
        layer1[9][15:8] = buffer_data_1[103:96];
        layer1[9][23:16] = buffer_data_1[111:104];
        layer2[9][7:0] = buffer_data_0[95:88];
        layer2[9][15:8] = buffer_data_0[103:96];
        layer2[9][23:16] = buffer_data_0[111:104];
        layer0[10][7:0] = buffer_data_2[103:96];
        layer0[10][15:8] = buffer_data_2[111:104];
        layer0[10][23:16] = buffer_data_2[119:112];
        layer1[10][7:0] = buffer_data_1[103:96];
        layer1[10][15:8] = buffer_data_1[111:104];
        layer1[10][23:16] = buffer_data_1[119:112];
        layer2[10][7:0] = buffer_data_0[103:96];
        layer2[10][15:8] = buffer_data_0[111:104];
        layer2[10][23:16] = buffer_data_0[119:112];
        layer0[11][7:0] = buffer_data_2[111:104];
        layer0[11][15:8] = buffer_data_2[119:112];
        layer0[11][23:16] = buffer_data_2[127:120];
        layer1[11][7:0] = buffer_data_1[111:104];
        layer1[11][15:8] = buffer_data_1[119:112];
        layer1[11][23:16] = buffer_data_1[127:120];
        layer2[11][7:0] = buffer_data_0[111:104];
        layer2[11][15:8] = buffer_data_0[119:112];
        layer2[11][23:16] = buffer_data_0[127:120];
        layer0[12][7:0] = buffer_data_2[119:112];
        layer0[12][15:8] = buffer_data_2[127:120];
        layer0[12][23:16] = buffer_data_2[135:128];
        layer1[12][7:0] = buffer_data_1[119:112];
        layer1[12][15:8] = buffer_data_1[127:120];
        layer1[12][23:16] = buffer_data_1[135:128];
        layer2[12][7:0] = buffer_data_0[119:112];
        layer2[12][15:8] = buffer_data_0[127:120];
        layer2[12][23:16] = buffer_data_0[135:128];
        layer0[13][7:0] = buffer_data_2[127:120];
        layer0[13][15:8] = buffer_data_2[135:128];
        layer0[13][23:16] = buffer_data_2[143:136];
        layer1[13][7:0] = buffer_data_1[127:120];
        layer1[13][15:8] = buffer_data_1[135:128];
        layer1[13][23:16] = buffer_data_1[143:136];
        layer2[13][7:0] = buffer_data_0[127:120];
        layer2[13][15:8] = buffer_data_0[135:128];
        layer2[13][23:16] = buffer_data_0[143:136];
        layer0[14][7:0] = buffer_data_2[135:128];
        layer0[14][15:8] = buffer_data_2[143:136];
        layer0[14][23:16] = buffer_data_2[151:144];
        layer1[14][7:0] = buffer_data_1[135:128];
        layer1[14][15:8] = buffer_data_1[143:136];
        layer1[14][23:16] = buffer_data_1[151:144];
        layer2[14][7:0] = buffer_data_0[135:128];
        layer2[14][15:8] = buffer_data_0[143:136];
        layer2[14][23:16] = buffer_data_0[151:144];
        layer0[15][7:0] = buffer_data_2[143:136];
        layer0[15][15:8] = buffer_data_2[151:144];
        layer0[15][23:16] = 0;
        layer1[15][7:0] = buffer_data_1[143:136];
        layer1[15][15:8] = buffer_data_1[151:144];
        layer1[15][23:16] = 0;
        layer2[15][7:0] = buffer_data_0[143:136];
        layer2[15][15:8] = buffer_data_0[151:144];
        layer2[15][23:16] = 0;
    end
    default: begin
        layer0[0][7:0] = 'd0;
        layer0[0][15:8] = 'd0;
        layer0[0][23:16] = 'd0;
        layer1[0][7:0] = 'd0;
        layer1[0][15:8] = 'd0;
        layer1[0][23:16] = 'd0;
        layer2[0][7:0] = 'd0;
        layer2[0][15:8] = 'd0;
        layer2[0][23:16] = 'd0;
        layer0[1][7:0] = 'd0;
        layer0[1][15:8] = 'd0;
        layer0[1][23:16] = 'd0;
        layer1[1][7:0] = 'd0;
        layer1[1][15:8] = 'd0;
        layer1[1][23:16] = 'd0;
        layer2[1][7:0] = 'd0;
        layer2[1][15:8] = 'd0;
        layer2[1][23:16] = 'd0;
        layer0[2][7:0] = 'd0;
        layer0[2][15:8] = 'd0;
        layer0[2][23:16] = 'd0;
        layer1[2][7:0] = 'd0;
        layer1[2][15:8] = 'd0;
        layer1[2][23:16] = 'd0;
        layer2[2][7:0] = 'd0;
        layer2[2][15:8] = 'd0;
        layer2[2][23:16] = 'd0;
        layer0[3][7:0] = 'd0;
        layer0[3][15:8] = 'd0;
        layer0[3][23:16] = 'd0;
        layer1[3][7:0] = 'd0;
        layer1[3][15:8] = 'd0;
        layer1[3][23:16] = 'd0;
        layer2[3][7:0] = 'd0;
        layer2[3][15:8] = 'd0;
        layer2[3][23:16] = 'd0;
        layer0[4][7:0] = 'd0;
        layer0[4][15:8] = 'd0;
        layer0[4][23:16] = 'd0;
        layer1[4][7:0] = 'd0;
        layer1[4][15:8] = 'd0;
        layer1[4][23:16] = 'd0;
        layer2[4][7:0] = 'd0;
        layer2[4][15:8] = 'd0;
        layer2[4][23:16] = 'd0;
        layer0[5][7:0] = 'd0;
        layer0[5][15:8] = 'd0;
        layer0[5][23:16] = 'd0;
        layer1[5][7:0] = 'd0;
        layer1[5][15:8] = 'd0;
        layer1[5][23:16] = 'd0;
        layer2[5][7:0] = 'd0;
        layer2[5][15:8] = 'd0;
        layer2[5][23:16] = 'd0;
        layer0[6][7:0] = 'd0;
        layer0[6][15:8] = 'd0;
        layer0[6][23:16] = 'd0;
        layer1[6][7:0] = 'd0;
        layer1[6][15:8] = 'd0;
        layer1[6][23:16] = 'd0;
        layer2[6][7:0] = 'd0;
        layer2[6][15:8] = 'd0;
        layer2[6][23:16] = 'd0;
        layer0[7][7:0] = 'd0;
        layer0[7][15:8] = 'd0;
        layer0[7][23:16] = 'd0;
        layer1[7][7:0] = 'd0;
        layer1[7][15:8] = 'd0;
        layer1[7][23:16] = 'd0;
        layer2[7][7:0] = 'd0;
        layer2[7][15:8] = 'd0;
        layer2[7][23:16] = 'd0;
        layer0[8][7:0] = 'd0;
        layer0[8][15:8] = 'd0;
        layer0[8][23:16] = 'd0;
        layer1[8][7:0] = 'd0;
        layer1[8][15:8] = 'd0;
        layer1[8][23:16] = 'd0;
        layer2[8][7:0] = 'd0;
        layer2[8][15:8] = 'd0;
        layer2[8][23:16] = 'd0;
        layer0[9][7:0] = 'd0;
        layer0[9][15:8] = 'd0;
        layer0[9][23:16] = 'd0;
        layer1[9][7:0] = 'd0;
        layer1[9][15:8] = 'd0;
        layer1[9][23:16] = 'd0;
        layer2[9][7:0] = 'd0;
        layer2[9][15:8] = 'd0;
        layer2[9][23:16] = 'd0;
        layer0[10][7:0] = 'd0;
        layer0[10][15:8] = 'd0;
        layer0[10][23:16] = 'd0;
        layer1[10][7:0] = 'd0;
        layer1[10][15:8] = 'd0;
        layer1[10][23:16] = 'd0;
        layer2[10][7:0] = 'd0;
        layer2[10][15:8] = 'd0;
        layer2[10][23:16] = 'd0;
        layer0[11][7:0] = 'd0;
        layer0[11][15:8] = 'd0;
        layer0[11][23:16] = 'd0;
        layer1[11][7:0] = 'd0;
        layer1[11][15:8] = 'd0;
        layer1[11][23:16] = 'd0;
        layer2[11][7:0] = 'd0;
        layer2[11][15:8] = 'd0;
        layer2[11][23:16] = 'd0;
        layer0[12][7:0] = 'd0;
        layer0[12][15:8] = 'd0;
        layer0[12][23:16] = 'd0;
        layer1[12][7:0] = 'd0;
        layer1[12][15:8] = 'd0;
        layer1[12][23:16] = 'd0;
        layer2[12][7:0] = 'd0;
        layer2[12][15:8] = 'd0;
        layer2[12][23:16] = 'd0;
        layer0[13][7:0] = 'd0;
        layer0[13][15:8] = 'd0;
        layer0[13][23:16] = 'd0;
        layer1[13][7:0] = 'd0;
        layer1[13][15:8] = 'd0;
        layer1[13][23:16] = 'd0;
        layer2[13][7:0] = 'd0;
        layer2[13][15:8] = 'd0;
        layer2[13][23:16] = 'd0;
        layer0[14][7:0] = 'd0;
        layer0[14][15:8] = 'd0;
        layer0[14][23:16] = 'd0;
        layer1[14][7:0] = 'd0;
        layer1[14][15:8] = 'd0;
        layer1[14][23:16] = 'd0;
        layer2[14][7:0] = 'd0;
        layer2[14][15:8] = 'd0;
        layer2[14][23:16] = 'd0;
        layer0[15][7:0] = 'd0;
        layer0[15][15:8] = 'd0;
        layer0[15][23:16] = 'd0;
        layer1[15][7:0] = 'd0;
        layer1[15][15:8] = 'd0;
        layer1[15][23:16] = 'd0;
        layer2[15][7:0] = 'd0;
        layer2[15][15:8] = 'd0;
        layer2[15][23:16] = 'd0;
    end
  endcase
end

wire  [39:0]  kernel_img_mul_0[0:8];
assign kernel_img_mul_0[0] = layer0[0][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_0[1] = layer0[0][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_0[2] = layer0[0][23:16] *  G_Kernel_3x3[0][95:64];
assign kernel_img_mul_0[3] = layer1[0][7:0] *  G_Kernel_3x3[1][31:0];
assign kernel_img_mul_0[4] = layer1[0][15:8] *  G_Kernel_3x3[1][63:32];
assign kernel_img_mul_0[5] = layer1[0][23:16] *  G_Kernel_3x3[1][95:64];
assign kernel_img_mul_0[6] = layer2[0][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_0[7] = layer2[0][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_0[8] = layer2[0][23:16] *  G_Kernel_3x3[0][95:64];
wire  [39:0]  kernel_img_sum_0 = kernel_img_mul_0[0] + kernel_img_mul_0[1] + kernel_img_mul_0[2] + 
                kernel_img_mul_0[3] + kernel_img_mul_0[4] + kernel_img_mul_0[5] + 
                kernel_img_mul_0[6] + kernel_img_mul_0[7] + kernel_img_mul_0[8];
wire  [39:0]  kernel_img_mul_1[0:8];
assign kernel_img_mul_1[0] = layer0[1][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_1[1] = layer0[1][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_1[2] = layer0[1][23:16] *  G_Kernel_3x3[0][95:64];
assign kernel_img_mul_1[3] = layer1[1][7:0] *  G_Kernel_3x3[1][31:0];
assign kernel_img_mul_1[4] = layer1[1][15:8] *  G_Kernel_3x3[1][63:32];
assign kernel_img_mul_1[5] = layer1[1][23:16] *  G_Kernel_3x3[1][95:64];
assign kernel_img_mul_1[6] = layer2[1][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_1[7] = layer2[1][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_1[8] = layer2[1][23:16] *  G_Kernel_3x3[0][95:64];
wire  [39:0]  kernel_img_sum_1 = kernel_img_mul_1[0] + kernel_img_mul_1[1] + kernel_img_mul_1[2] + 
                kernel_img_mul_1[3] + kernel_img_mul_1[4] + kernel_img_mul_1[5] + 
                kernel_img_mul_1[6] + kernel_img_mul_1[7] + kernel_img_mul_1[8];
wire  [39:0]  kernel_img_mul_2[0:8];
assign kernel_img_mul_2[0] = layer0[2][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_2[1] = layer0[2][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_2[2] = layer0[2][23:16] *  G_Kernel_3x3[0][95:64];
assign kernel_img_mul_2[3] = layer1[2][7:0] *  G_Kernel_3x3[1][31:0];
assign kernel_img_mul_2[4] = layer1[2][15:8] *  G_Kernel_3x3[1][63:32];
assign kernel_img_mul_2[5] = layer1[2][23:16] *  G_Kernel_3x3[1][95:64];
assign kernel_img_mul_2[6] = layer2[2][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_2[7] = layer2[2][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_2[8] = layer2[2][23:16] *  G_Kernel_3x3[0][95:64];
wire  [39:0]  kernel_img_sum_2 = kernel_img_mul_2[0] + kernel_img_mul_2[1] + kernel_img_mul_2[2] + 
                kernel_img_mul_2[3] + kernel_img_mul_2[4] + kernel_img_mul_2[5] + 
                kernel_img_mul_2[6] + kernel_img_mul_2[7] + kernel_img_mul_2[8];
wire  [39:0]  kernel_img_mul_3[0:8];
assign kernel_img_mul_3[0] = layer0[3][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_3[1] = layer0[3][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_3[2] = layer0[3][23:16] *  G_Kernel_3x3[0][95:64];
assign kernel_img_mul_3[3] = layer1[3][7:0] *  G_Kernel_3x3[1][31:0];
assign kernel_img_mul_3[4] = layer1[3][15:8] *  G_Kernel_3x3[1][63:32];
assign kernel_img_mul_3[5] = layer1[3][23:16] *  G_Kernel_3x3[1][95:64];
assign kernel_img_mul_3[6] = layer2[3][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_3[7] = layer2[3][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_3[8] = layer2[3][23:16] *  G_Kernel_3x3[0][95:64];
wire  [39:0]  kernel_img_sum_3 = kernel_img_mul_3[0] + kernel_img_mul_3[1] + kernel_img_mul_3[2] + 
                kernel_img_mul_3[3] + kernel_img_mul_3[4] + kernel_img_mul_3[5] + 
                kernel_img_mul_3[6] + kernel_img_mul_3[7] + kernel_img_mul_3[8];
wire  [39:0]  kernel_img_mul_4[0:8];
assign kernel_img_mul_4[0] = layer0[4][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_4[1] = layer0[4][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_4[2] = layer0[4][23:16] *  G_Kernel_3x3[0][95:64];
assign kernel_img_mul_4[3] = layer1[4][7:0] *  G_Kernel_3x3[1][31:0];
assign kernel_img_mul_4[4] = layer1[4][15:8] *  G_Kernel_3x3[1][63:32];
assign kernel_img_mul_4[5] = layer1[4][23:16] *  G_Kernel_3x3[1][95:64];
assign kernel_img_mul_4[6] = layer2[4][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_4[7] = layer2[4][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_4[8] = layer2[4][23:16] *  G_Kernel_3x3[0][95:64];
wire  [39:0]  kernel_img_sum_4 = kernel_img_mul_4[0] + kernel_img_mul_4[1] + kernel_img_mul_4[2] + 
                kernel_img_mul_4[3] + kernel_img_mul_4[4] + kernel_img_mul_4[5] + 
                kernel_img_mul_4[6] + kernel_img_mul_4[7] + kernel_img_mul_4[8];
wire  [39:0]  kernel_img_mul_5[0:8];
assign kernel_img_mul_5[0] = layer0[5][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_5[1] = layer0[5][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_5[2] = layer0[5][23:16] *  G_Kernel_3x3[0][95:64];
assign kernel_img_mul_5[3] = layer1[5][7:0] *  G_Kernel_3x3[1][31:0];
assign kernel_img_mul_5[4] = layer1[5][15:8] *  G_Kernel_3x3[1][63:32];
assign kernel_img_mul_5[5] = layer1[5][23:16] *  G_Kernel_3x3[1][95:64];
assign kernel_img_mul_5[6] = layer2[5][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_5[7] = layer2[5][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_5[8] = layer2[5][23:16] *  G_Kernel_3x3[0][95:64];
wire  [39:0]  kernel_img_sum_5 = kernel_img_mul_5[0] + kernel_img_mul_5[1] + kernel_img_mul_5[2] + 
                kernel_img_mul_5[3] + kernel_img_mul_5[4] + kernel_img_mul_5[5] + 
                kernel_img_mul_5[6] + kernel_img_mul_5[7] + kernel_img_mul_5[8];
wire  [39:0]  kernel_img_mul_6[0:8];
assign kernel_img_mul_6[0] = layer0[6][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_6[1] = layer0[6][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_6[2] = layer0[6][23:16] *  G_Kernel_3x3[0][95:64];
assign kernel_img_mul_6[3] = layer1[6][7:0] *  G_Kernel_3x3[1][31:0];
assign kernel_img_mul_6[4] = layer1[6][15:8] *  G_Kernel_3x3[1][63:32];
assign kernel_img_mul_6[5] = layer1[6][23:16] *  G_Kernel_3x3[1][95:64];
assign kernel_img_mul_6[6] = layer2[6][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_6[7] = layer2[6][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_6[8] = layer2[6][23:16] *  G_Kernel_3x3[0][95:64];
wire  [39:0]  kernel_img_sum_6 = kernel_img_mul_6[0] + kernel_img_mul_6[1] + kernel_img_mul_6[2] + 
                kernel_img_mul_6[3] + kernel_img_mul_6[4] + kernel_img_mul_6[5] + 
                kernel_img_mul_6[6] + kernel_img_mul_6[7] + kernel_img_mul_6[8];
wire  [39:0]  kernel_img_mul_7[0:8];
assign kernel_img_mul_7[0] = layer0[7][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_7[1] = layer0[7][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_7[2] = layer0[7][23:16] *  G_Kernel_3x3[0][95:64];
assign kernel_img_mul_7[3] = layer1[7][7:0] *  G_Kernel_3x3[1][31:0];
assign kernel_img_mul_7[4] = layer1[7][15:8] *  G_Kernel_3x3[1][63:32];
assign kernel_img_mul_7[5] = layer1[7][23:16] *  G_Kernel_3x3[1][95:64];
assign kernel_img_mul_7[6] = layer2[7][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_7[7] = layer2[7][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_7[8] = layer2[7][23:16] *  G_Kernel_3x3[0][95:64];
wire  [39:0]  kernel_img_sum_7 = kernel_img_mul_7[0] + kernel_img_mul_7[1] + kernel_img_mul_7[2] + 
                kernel_img_mul_7[3] + kernel_img_mul_7[4] + kernel_img_mul_7[5] + 
                kernel_img_mul_7[6] + kernel_img_mul_7[7] + kernel_img_mul_7[8];
wire  [39:0]  kernel_img_mul_8[0:8];
assign kernel_img_mul_8[0] = layer0[8][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_8[1] = layer0[8][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_8[2] = layer0[8][23:16] *  G_Kernel_3x3[0][95:64];
assign kernel_img_mul_8[3] = layer1[8][7:0] *  G_Kernel_3x3[1][31:0];
assign kernel_img_mul_8[4] = layer1[8][15:8] *  G_Kernel_3x3[1][63:32];
assign kernel_img_mul_8[5] = layer1[8][23:16] *  G_Kernel_3x3[1][95:64];
assign kernel_img_mul_8[6] = layer2[8][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_8[7] = layer2[8][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_8[8] = layer2[8][23:16] *  G_Kernel_3x3[0][95:64];
wire  [39:0]  kernel_img_sum_8 = kernel_img_mul_8[0] + kernel_img_mul_8[1] + kernel_img_mul_8[2] + 
                kernel_img_mul_8[3] + kernel_img_mul_8[4] + kernel_img_mul_8[5] + 
                kernel_img_mul_8[6] + kernel_img_mul_8[7] + kernel_img_mul_8[8];
wire  [39:0]  kernel_img_mul_9[0:8];
assign kernel_img_mul_9[0] = layer0[9][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_9[1] = layer0[9][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_9[2] = layer0[9][23:16] *  G_Kernel_3x3[0][95:64];
assign kernel_img_mul_9[3] = layer1[9][7:0] *  G_Kernel_3x3[1][31:0];
assign kernel_img_mul_9[4] = layer1[9][15:8] *  G_Kernel_3x3[1][63:32];
assign kernel_img_mul_9[5] = layer1[9][23:16] *  G_Kernel_3x3[1][95:64];
assign kernel_img_mul_9[6] = layer2[9][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_9[7] = layer2[9][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_9[8] = layer2[9][23:16] *  G_Kernel_3x3[0][95:64];
wire  [39:0]  kernel_img_sum_9 = kernel_img_mul_9[0] + kernel_img_mul_9[1] + kernel_img_mul_9[2] + 
                kernel_img_mul_9[3] + kernel_img_mul_9[4] + kernel_img_mul_9[5] + 
                kernel_img_mul_9[6] + kernel_img_mul_9[7] + kernel_img_mul_9[8];
wire  [39:0]  kernel_img_mul_10[0:8];
assign kernel_img_mul_10[0] = layer0[10][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_10[1] = layer0[10][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_10[2] = layer0[10][23:16] *  G_Kernel_3x3[0][95:64];
assign kernel_img_mul_10[3] = layer1[10][7:0] *  G_Kernel_3x3[1][31:0];
assign kernel_img_mul_10[4] = layer1[10][15:8] *  G_Kernel_3x3[1][63:32];
assign kernel_img_mul_10[5] = layer1[10][23:16] *  G_Kernel_3x3[1][95:64];
assign kernel_img_mul_10[6] = layer2[10][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_10[7] = layer2[10][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_10[8] = layer2[10][23:16] *  G_Kernel_3x3[0][95:64];
wire  [39:0]  kernel_img_sum_10 = kernel_img_mul_10[0] + kernel_img_mul_10[1] + kernel_img_mul_10[2] + 
                kernel_img_mul_10[3] + kernel_img_mul_10[4] + kernel_img_mul_10[5] + 
                kernel_img_mul_10[6] + kernel_img_mul_10[7] + kernel_img_mul_10[8];
wire  [39:0]  kernel_img_mul_11[0:8];
assign kernel_img_mul_11[0] = layer0[11][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_11[1] = layer0[11][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_11[2] = layer0[11][23:16] *  G_Kernel_3x3[0][95:64];
assign kernel_img_mul_11[3] = layer1[11][7:0] *  G_Kernel_3x3[1][31:0];
assign kernel_img_mul_11[4] = layer1[11][15:8] *  G_Kernel_3x3[1][63:32];
assign kernel_img_mul_11[5] = layer1[11][23:16] *  G_Kernel_3x3[1][95:64];
assign kernel_img_mul_11[6] = layer2[11][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_11[7] = layer2[11][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_11[8] = layer2[11][23:16] *  G_Kernel_3x3[0][95:64];
wire  [39:0]  kernel_img_sum_11 = kernel_img_mul_11[0] + kernel_img_mul_11[1] + kernel_img_mul_11[2] + 
                kernel_img_mul_11[3] + kernel_img_mul_11[4] + kernel_img_mul_11[5] + 
                kernel_img_mul_11[6] + kernel_img_mul_11[7] + kernel_img_mul_11[8];
wire  [39:0]  kernel_img_mul_12[0:8];
assign kernel_img_mul_12[0] = layer0[12][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_12[1] = layer0[12][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_12[2] = layer0[12][23:16] *  G_Kernel_3x3[0][95:64];
assign kernel_img_mul_12[3] = layer1[12][7:0] *  G_Kernel_3x3[1][31:0];
assign kernel_img_mul_12[4] = layer1[12][15:8] *  G_Kernel_3x3[1][63:32];
assign kernel_img_mul_12[5] = layer1[12][23:16] *  G_Kernel_3x3[1][95:64];
assign kernel_img_mul_12[6] = layer2[12][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_12[7] = layer2[12][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_12[8] = layer2[12][23:16] *  G_Kernel_3x3[0][95:64];
wire  [39:0]  kernel_img_sum_12 = kernel_img_mul_12[0] + kernel_img_mul_12[1] + kernel_img_mul_12[2] + 
                kernel_img_mul_12[3] + kernel_img_mul_12[4] + kernel_img_mul_12[5] + 
                kernel_img_mul_12[6] + kernel_img_mul_12[7] + kernel_img_mul_12[8];
wire  [39:0]  kernel_img_mul_13[0:8];
assign kernel_img_mul_13[0] = layer0[13][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_13[1] = layer0[13][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_13[2] = layer0[13][23:16] *  G_Kernel_3x3[0][95:64];
assign kernel_img_mul_13[3] = layer1[13][7:0] *  G_Kernel_3x3[1][31:0];
assign kernel_img_mul_13[4] = layer1[13][15:8] *  G_Kernel_3x3[1][63:32];
assign kernel_img_mul_13[5] = layer1[13][23:16] *  G_Kernel_3x3[1][95:64];
assign kernel_img_mul_13[6] = layer2[13][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_13[7] = layer2[13][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_13[8] = layer2[13][23:16] *  G_Kernel_3x3[0][95:64];
wire  [39:0]  kernel_img_sum_13 = kernel_img_mul_13[0] + kernel_img_mul_13[1] + kernel_img_mul_13[2] + 
                kernel_img_mul_13[3] + kernel_img_mul_13[4] + kernel_img_mul_13[5] + 
                kernel_img_mul_13[6] + kernel_img_mul_13[7] + kernel_img_mul_13[8];
wire  [39:0]  kernel_img_mul_14[0:8];
assign kernel_img_mul_14[0] = layer0[14][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_14[1] = layer0[14][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_14[2] = layer0[14][23:16] *  G_Kernel_3x3[0][95:64];
assign kernel_img_mul_14[3] = layer1[14][7:0] *  G_Kernel_3x3[1][31:0];
assign kernel_img_mul_14[4] = layer1[14][15:8] *  G_Kernel_3x3[1][63:32];
assign kernel_img_mul_14[5] = layer1[14][23:16] *  G_Kernel_3x3[1][95:64];
assign kernel_img_mul_14[6] = layer2[14][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_14[7] = layer2[14][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_14[8] = layer2[14][23:16] *  G_Kernel_3x3[0][95:64];
wire  [39:0]  kernel_img_sum_14 = kernel_img_mul_14[0] + kernel_img_mul_14[1] + kernel_img_mul_14[2] + 
                kernel_img_mul_14[3] + kernel_img_mul_14[4] + kernel_img_mul_14[5] + 
                kernel_img_mul_14[6] + kernel_img_mul_14[7] + kernel_img_mul_14[8];
wire  [39:0]  kernel_img_mul_15[0:8];
assign kernel_img_mul_15[0] = layer0[15][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_15[1] = layer0[15][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_15[2] = layer0[15][23:16] *  G_Kernel_3x3[0][95:64];
assign kernel_img_mul_15[3] = layer1[15][7:0] *  G_Kernel_3x3[1][31:0];
assign kernel_img_mul_15[4] = layer1[15][15:8] *  G_Kernel_3x3[1][63:32];
assign kernel_img_mul_15[5] = layer1[15][23:16] *  G_Kernel_3x3[1][95:64];
assign kernel_img_mul_15[6] = layer2[15][7:0] *  G_Kernel_3x3[0][31:0];
assign kernel_img_mul_15[7] = layer2[15][15:8] *  G_Kernel_3x3[0][63:32];
assign kernel_img_mul_15[8] = layer2[15][23:16] *  G_Kernel_3x3[0][95:64];
wire  [39:0]  kernel_img_sum_15 = kernel_img_mul_15[0] + kernel_img_mul_15[1] + kernel_img_mul_15[2] + 
                kernel_img_mul_15[3] + kernel_img_mul_15[4] + kernel_img_mul_15[5] + 
                kernel_img_mul_15[6] + kernel_img_mul_15[7] + kernel_img_mul_15[8];
always @(*) begin
    blur_out[7:0] = kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
    blur_out[15:8] = kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
    blur_out[23:16] = kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
    blur_out[31:24] = kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
    blur_out[39:32] = kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
    blur_out[47:40] = kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
    blur_out[55:48] = kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
    blur_out[63:56] = kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
    blur_out[71:64] = kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
    blur_out[79:72] = kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
    blur_out[87:80] = kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
    blur_out[95:88] = kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
    blur_out[103:96] = kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
    blur_out[111:104] = kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
    blur_out[119:112] = kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
    blur_out[127:120] = kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
end


endmodule