module Gaussian_Blur_5x5_0(
  clk,
  rst_n,
  buffer_data_0,
  buffer_data_1,
  buffer_data_2,
  buffer_data_3,
  buffer_data_4,
  current_col,
  blur_out,
  start,
  done
);

input                 clk;
input                 rst_n;
input                 start;
output                done;
input         [5:0]   current_col;
input       [175:0]   buffer_data_0;
input       [175:0]   buffer_data_1;
input       [175:0]   buffer_data_2;
input       [175:0]   buffer_data_3;
input       [175:0]   buffer_data_4;
output reg  [127:0]   blur_out; // wire

parameter  ST_MUX         = 0,
           ST_MUL         = 1,
           ST_ADD         = 2,
           ST_UPDATE      = 3;
reg     [2:0] current_state,
              next_state;
assign done = (current_state==ST_UPDATE) ? 1 : 0;

wire       [39:0]  G_Kernel_5x5_0;
wire       [39:0]  G_Kernel_5x5_1;
wire       [39:0]  G_Kernel_5x5_2;
assign  G_Kernel_5x5_0[7:0]   = 8'h05; //F2F79A;  // 18'b000001011111001011;//'d023238;
assign  G_Kernel_5x5_0[15:8]  = 8'h08; //A86809;  // 18'b000010001010100001;//d033819;
assign  G_Kernel_5x5_0[23:16] = 8'h09; //CFB50A;  // 18'b000010011100111110;//d038325;
assign  G_Kernel_5x5_0[31:24] = 8'h08; //A86809;  // 18'b000010001010100001;//d033819;
assign  G_Kernel_5x5_0[39:32] = 8'h05; //F2F79A;  // 18'b000001011111001011;//'d023238;
assign  G_Kernel_5x5_1[7:0]   = 8'h08; //A86809;  // 18'b000010001010100001;//d033819;
assign  G_Kernel_5x5_1[15:8]  = 8'h0C; //999546;  // 18'b000011001001100110;//d049218;
assign  G_Kernel_5x5_1[23:16] = 8'h0E; //475732;  // 18'b000011100100011101;//d055776;
assign  G_Kernel_5x5_1[31:24] = 8'h0C; //999546;  // 18'b000011001001100110;//d049218;
assign  G_Kernel_5x5_1[39:32] = 8'h08; //A86809;  // 18'b000010001010100001;//d033819;
assign  G_Kernel_5x5_2[7:0]   = 8'h09; //CFB50A;  // 18'b000010011100111110;//d038325;
assign  G_Kernel_5x5_2[15:8]  = 8'h0E; //475732;  // 18'b000011100100011101;//d055776;
assign  G_Kernel_5x5_2[23:16] = 8'h10; //2E5B3F;  // 18'b000100000010111001;//d063207;
assign  G_Kernel_5x5_2[31:24] = 8'h0E; //475732;  // 18'b000011100100011101;//d055776;
assign  G_Kernel_5x5_2[39:32] = 8'h09; //CFB50A;  // 18'b000010011100111110;//d038325;

reg    [39:0]    layer0[0:15]; //wire
reg    [39:0]    layer1[0:15]; //wire
reg    [39:0]    layer2[0:15]; //wire
reg    [39:0]    layer3[0:15]; //wire
reg    [39:0]    layer4[0:15]; //wire
always @(posedge clk) begin
  if(!rst_n) begin
    layer0[0] <= 'd0;
    layer0[1] <= 'd0;
    layer0[2] <= 'd0;
    layer0[3] <= 'd0;
    layer0[4] <= 'd0;
    layer0[5] <= 'd0;
    layer0[6] <= 'd0;
    layer0[7] <= 'd0;
    layer0[8] <= 'd0;
    layer0[9] <= 'd0;
    layer0[10] <= 'd0;
    layer0[11] <= 'd0;
    layer0[12] <= 'd0;
    layer0[13] <= 'd0;
    layer0[14] <= 'd0;
    layer0[15] <= 'd0;
    layer1[0] <= 'd0;
    layer1[1] <= 'd0;
    layer1[2] <= 'd0;
    layer1[3] <= 'd0;
    layer1[4] <= 'd0;
    layer1[5] <= 'd0;
    layer1[6] <= 'd0;
    layer1[7] <= 'd0;
    layer1[8] <= 'd0;
    layer1[9] <= 'd0;
    layer1[10] <= 'd0;
    layer1[11] <= 'd0;
    layer1[12] <= 'd0;
    layer1[13] <= 'd0;
    layer1[14] <= 'd0;
    layer1[15] <= 'd0;
    layer2[0] <= 'd0;
    layer2[1] <= 'd0;
    layer2[2] <= 'd0;
    layer2[3] <= 'd0;
    layer2[4] <= 'd0;
    layer2[5] <= 'd0;
    layer2[6] <= 'd0;
    layer2[7] <= 'd0;
    layer2[8] <= 'd0;
    layer2[9] <= 'd0;
    layer2[10] <= 'd0;
    layer2[11] <= 'd0;
    layer2[12] <= 'd0;
    layer2[13] <= 'd0;
    layer2[14] <= 'd0;
    layer2[15] <= 'd0;
    layer3[0] <= 'd0;
    layer3[1] <= 'd0;
    layer3[2] <= 'd0;
    layer3[3] <= 'd0;
    layer3[4] <= 'd0;
    layer3[5] <= 'd0;
    layer3[6] <= 'd0;
    layer3[7] <= 'd0;
    layer3[8] <= 'd0;
    layer3[9] <= 'd0;
    layer3[10] <= 'd0;
    layer3[11] <= 'd0;
    layer3[12] <= 'd0;
    layer3[13] <= 'd0;
    layer3[14] <= 'd0;
    layer3[15] <= 'd0;
    layer4[0] <= 'd0;
    layer4[1] <= 'd0;
    layer4[2] <= 'd0;
    layer4[3] <= 'd0;
    layer4[4] <= 'd0;
    layer4[5] <= 'd0;
    layer4[6] <= 'd0;
    layer4[7] <= 'd0;
    layer4[8] <= 'd0;
    layer4[9] <= 'd0;
    layer4[10] <= 'd0;
    layer4[11] <= 'd0;
    layer4[12] <= 'd0;
    layer4[13] <= 'd0;
    layer4[14] <= 'd0;
    layer4[15] <= 'd0;
  end
  else if(current_state==ST_MUX) begin
    case(current_col)
      'd0: begin
        layer0[0][7:0] <= 0;
        layer0[0][15:8] <= 0;
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= 0;
        layer1[0][15:8] <= 0;
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= 0;
        layer2[0][15:8] <= 0;
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= 0;
        layer3[0][15:8] <= 0;
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= 0;
        layer4[0][15:8] <= 0;
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= 0;
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= 0;
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= 0;
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= 0;
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= 0;
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd1: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd2: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd3: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd4: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd5: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd6: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd7: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd8: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd9: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd10: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd11: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd12: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd13: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd14: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd15: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd16: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd17: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd18: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd19: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd20: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd21: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd22: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd23: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd24: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd25: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd26: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd27: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd28: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd29: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd30: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd31: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd32: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd33: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd34: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd35: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd36: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd37: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd38: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= buffer_data_4[159:152];
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= buffer_data_3[159:152];
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= buffer_data_2[159:152];
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= buffer_data_1[159:152];
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= buffer_data_0[159:152];
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= buffer_data_4[159:152];
        layer0[15][39:32] <= buffer_data_4[167:160];
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= buffer_data_3[159:152];
        layer1[15][39:32] <= buffer_data_3[167:160];
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= buffer_data_2[159:152];
        layer2[15][39:32] <= buffer_data_2[167:160];
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= buffer_data_1[159:152];
        layer3[15][39:32] <= buffer_data_1[167:160];
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= buffer_data_0[159:152];
        layer4[15][39:32] <= buffer_data_0[167:160];
    end
      'd39: begin
        layer0[0][7:0] <= buffer_data_4[15:8];
        layer0[0][15:8] <= buffer_data_4[23:16];
        layer0[0][23:16] <= buffer_data_4[31:24];
        layer0[0][31:24] <= buffer_data_4[39:32];
        layer0[0][39:32] <= buffer_data_4[47:40];
        layer1[0][7:0] <= buffer_data_3[15:8];
        layer1[0][15:8] <= buffer_data_3[23:16];
        layer1[0][23:16] <= buffer_data_3[31:24];
        layer1[0][31:24] <= buffer_data_3[39:32];
        layer1[0][39:32] <= buffer_data_3[47:40];
        layer2[0][7:0] <= buffer_data_2[15:8];
        layer2[0][15:8] <= buffer_data_2[23:16];
        layer2[0][23:16] <= buffer_data_2[31:24];
        layer2[0][31:24] <= buffer_data_2[39:32];
        layer2[0][39:32] <= buffer_data_2[47:40];
        layer3[0][7:0] <= buffer_data_1[15:8];
        layer3[0][15:8] <= buffer_data_1[23:16];
        layer3[0][23:16] <= buffer_data_1[31:24];
        layer3[0][31:24] <= buffer_data_1[39:32];
        layer3[0][39:32] <= buffer_data_1[47:40];
        layer4[0][7:0] <= buffer_data_0[15:8];
        layer4[0][15:8] <= buffer_data_0[23:16];
        layer4[0][23:16] <= buffer_data_0[31:24];
        layer4[0][31:24] <= buffer_data_0[39:32];
        layer4[0][39:32] <= buffer_data_0[47:40];
        layer0[1][7:0] <= buffer_data_4[23:16];
        layer0[1][15:8] <= buffer_data_4[31:24];
        layer0[1][23:16] <= buffer_data_4[39:32];
        layer0[1][31:24] <= buffer_data_4[47:40];
        layer0[1][39:32] <= buffer_data_4[55:48];
        layer1[1][7:0] <= buffer_data_3[23:16];
        layer1[1][15:8] <= buffer_data_3[31:24];
        layer1[1][23:16] <= buffer_data_3[39:32];
        layer1[1][31:24] <= buffer_data_3[47:40];
        layer1[1][39:32] <= buffer_data_3[55:48];
        layer2[1][7:0] <= buffer_data_2[23:16];
        layer2[1][15:8] <= buffer_data_2[31:24];
        layer2[1][23:16] <= buffer_data_2[39:32];
        layer2[1][31:24] <= buffer_data_2[47:40];
        layer2[1][39:32] <= buffer_data_2[55:48];
        layer3[1][7:0] <= buffer_data_1[23:16];
        layer3[1][15:8] <= buffer_data_1[31:24];
        layer3[1][23:16] <= buffer_data_1[39:32];
        layer3[1][31:24] <= buffer_data_1[47:40];
        layer3[1][39:32] <= buffer_data_1[55:48];
        layer4[1][7:0] <= buffer_data_0[23:16];
        layer4[1][15:8] <= buffer_data_0[31:24];
        layer4[1][23:16] <= buffer_data_0[39:32];
        layer4[1][31:24] <= buffer_data_0[47:40];
        layer4[1][39:32] <= buffer_data_0[55:48];
        layer0[2][7:0] <= buffer_data_4[31:24];
        layer0[2][15:8] <= buffer_data_4[39:32];
        layer0[2][23:16] <= buffer_data_4[47:40];
        layer0[2][31:24] <= buffer_data_4[55:48];
        layer0[2][39:32] <= buffer_data_4[63:56];
        layer1[2][7:0] <= buffer_data_3[31:24];
        layer1[2][15:8] <= buffer_data_3[39:32];
        layer1[2][23:16] <= buffer_data_3[47:40];
        layer1[2][31:24] <= buffer_data_3[55:48];
        layer1[2][39:32] <= buffer_data_3[63:56];
        layer2[2][7:0] <= buffer_data_2[31:24];
        layer2[2][15:8] <= buffer_data_2[39:32];
        layer2[2][23:16] <= buffer_data_2[47:40];
        layer2[2][31:24] <= buffer_data_2[55:48];
        layer2[2][39:32] <= buffer_data_2[63:56];
        layer3[2][7:0] <= buffer_data_1[31:24];
        layer3[2][15:8] <= buffer_data_1[39:32];
        layer3[2][23:16] <= buffer_data_1[47:40];
        layer3[2][31:24] <= buffer_data_1[55:48];
        layer3[2][39:32] <= buffer_data_1[63:56];
        layer4[2][7:0] <= buffer_data_0[31:24];
        layer4[2][15:8] <= buffer_data_0[39:32];
        layer4[2][23:16] <= buffer_data_0[47:40];
        layer4[2][31:24] <= buffer_data_0[55:48];
        layer4[2][39:32] <= buffer_data_0[63:56];
        layer0[3][7:0] <= buffer_data_4[39:32];
        layer0[3][15:8] <= buffer_data_4[47:40];
        layer0[3][23:16] <= buffer_data_4[55:48];
        layer0[3][31:24] <= buffer_data_4[63:56];
        layer0[3][39:32] <= buffer_data_4[71:64];
        layer1[3][7:0] <= buffer_data_3[39:32];
        layer1[3][15:8] <= buffer_data_3[47:40];
        layer1[3][23:16] <= buffer_data_3[55:48];
        layer1[3][31:24] <= buffer_data_3[63:56];
        layer1[3][39:32] <= buffer_data_3[71:64];
        layer2[3][7:0] <= buffer_data_2[39:32];
        layer2[3][15:8] <= buffer_data_2[47:40];
        layer2[3][23:16] <= buffer_data_2[55:48];
        layer2[3][31:24] <= buffer_data_2[63:56];
        layer2[3][39:32] <= buffer_data_2[71:64];
        layer3[3][7:0] <= buffer_data_1[39:32];
        layer3[3][15:8] <= buffer_data_1[47:40];
        layer3[3][23:16] <= buffer_data_1[55:48];
        layer3[3][31:24] <= buffer_data_1[63:56];
        layer3[3][39:32] <= buffer_data_1[71:64];
        layer4[3][7:0] <= buffer_data_0[39:32];
        layer4[3][15:8] <= buffer_data_0[47:40];
        layer4[3][23:16] <= buffer_data_0[55:48];
        layer4[3][31:24] <= buffer_data_0[63:56];
        layer4[3][39:32] <= buffer_data_0[71:64];
        layer0[4][7:0] <= buffer_data_4[47:40];
        layer0[4][15:8] <= buffer_data_4[55:48];
        layer0[4][23:16] <= buffer_data_4[63:56];
        layer0[4][31:24] <= buffer_data_4[71:64];
        layer0[4][39:32] <= buffer_data_4[79:72];
        layer1[4][7:0] <= buffer_data_3[47:40];
        layer1[4][15:8] <= buffer_data_3[55:48];
        layer1[4][23:16] <= buffer_data_3[63:56];
        layer1[4][31:24] <= buffer_data_3[71:64];
        layer1[4][39:32] <= buffer_data_3[79:72];
        layer2[4][7:0] <= buffer_data_2[47:40];
        layer2[4][15:8] <= buffer_data_2[55:48];
        layer2[4][23:16] <= buffer_data_2[63:56];
        layer2[4][31:24] <= buffer_data_2[71:64];
        layer2[4][39:32] <= buffer_data_2[79:72];
        layer3[4][7:0] <= buffer_data_1[47:40];
        layer3[4][15:8] <= buffer_data_1[55:48];
        layer3[4][23:16] <= buffer_data_1[63:56];
        layer3[4][31:24] <= buffer_data_1[71:64];
        layer3[4][39:32] <= buffer_data_1[79:72];
        layer4[4][7:0] <= buffer_data_0[47:40];
        layer4[4][15:8] <= buffer_data_0[55:48];
        layer4[4][23:16] <= buffer_data_0[63:56];
        layer4[4][31:24] <= buffer_data_0[71:64];
        layer4[4][39:32] <= buffer_data_0[79:72];
        layer0[5][7:0] <= buffer_data_4[55:48];
        layer0[5][15:8] <= buffer_data_4[63:56];
        layer0[5][23:16] <= buffer_data_4[71:64];
        layer0[5][31:24] <= buffer_data_4[79:72];
        layer0[5][39:32] <= buffer_data_4[87:80];
        layer1[5][7:0] <= buffer_data_3[55:48];
        layer1[5][15:8] <= buffer_data_3[63:56];
        layer1[5][23:16] <= buffer_data_3[71:64];
        layer1[5][31:24] <= buffer_data_3[79:72];
        layer1[5][39:32] <= buffer_data_3[87:80];
        layer2[5][7:0] <= buffer_data_2[55:48];
        layer2[5][15:8] <= buffer_data_2[63:56];
        layer2[5][23:16] <= buffer_data_2[71:64];
        layer2[5][31:24] <= buffer_data_2[79:72];
        layer2[5][39:32] <= buffer_data_2[87:80];
        layer3[5][7:0] <= buffer_data_1[55:48];
        layer3[5][15:8] <= buffer_data_1[63:56];
        layer3[5][23:16] <= buffer_data_1[71:64];
        layer3[5][31:24] <= buffer_data_1[79:72];
        layer3[5][39:32] <= buffer_data_1[87:80];
        layer4[5][7:0] <= buffer_data_0[55:48];
        layer4[5][15:8] <= buffer_data_0[63:56];
        layer4[5][23:16] <= buffer_data_0[71:64];
        layer4[5][31:24] <= buffer_data_0[79:72];
        layer4[5][39:32] <= buffer_data_0[87:80];
        layer0[6][7:0] <= buffer_data_4[63:56];
        layer0[6][15:8] <= buffer_data_4[71:64];
        layer0[6][23:16] <= buffer_data_4[79:72];
        layer0[6][31:24] <= buffer_data_4[87:80];
        layer0[6][39:32] <= buffer_data_4[95:88];
        layer1[6][7:0] <= buffer_data_3[63:56];
        layer1[6][15:8] <= buffer_data_3[71:64];
        layer1[6][23:16] <= buffer_data_3[79:72];
        layer1[6][31:24] <= buffer_data_3[87:80];
        layer1[6][39:32] <= buffer_data_3[95:88];
        layer2[6][7:0] <= buffer_data_2[63:56];
        layer2[6][15:8] <= buffer_data_2[71:64];
        layer2[6][23:16] <= buffer_data_2[79:72];
        layer2[6][31:24] <= buffer_data_2[87:80];
        layer2[6][39:32] <= buffer_data_2[95:88];
        layer3[6][7:0] <= buffer_data_1[63:56];
        layer3[6][15:8] <= buffer_data_1[71:64];
        layer3[6][23:16] <= buffer_data_1[79:72];
        layer3[6][31:24] <= buffer_data_1[87:80];
        layer3[6][39:32] <= buffer_data_1[95:88];
        layer4[6][7:0] <= buffer_data_0[63:56];
        layer4[6][15:8] <= buffer_data_0[71:64];
        layer4[6][23:16] <= buffer_data_0[79:72];
        layer4[6][31:24] <= buffer_data_0[87:80];
        layer4[6][39:32] <= buffer_data_0[95:88];
        layer0[7][7:0] <= buffer_data_4[71:64];
        layer0[7][15:8] <= buffer_data_4[79:72];
        layer0[7][23:16] <= buffer_data_4[87:80];
        layer0[7][31:24] <= buffer_data_4[95:88];
        layer0[7][39:32] <= buffer_data_4[103:96];
        layer1[7][7:0] <= buffer_data_3[71:64];
        layer1[7][15:8] <= buffer_data_3[79:72];
        layer1[7][23:16] <= buffer_data_3[87:80];
        layer1[7][31:24] <= buffer_data_3[95:88];
        layer1[7][39:32] <= buffer_data_3[103:96];
        layer2[7][7:0] <= buffer_data_2[71:64];
        layer2[7][15:8] <= buffer_data_2[79:72];
        layer2[7][23:16] <= buffer_data_2[87:80];
        layer2[7][31:24] <= buffer_data_2[95:88];
        layer2[7][39:32] <= buffer_data_2[103:96];
        layer3[7][7:0] <= buffer_data_1[71:64];
        layer3[7][15:8] <= buffer_data_1[79:72];
        layer3[7][23:16] <= buffer_data_1[87:80];
        layer3[7][31:24] <= buffer_data_1[95:88];
        layer3[7][39:32] <= buffer_data_1[103:96];
        layer4[7][7:0] <= buffer_data_0[71:64];
        layer4[7][15:8] <= buffer_data_0[79:72];
        layer4[7][23:16] <= buffer_data_0[87:80];
        layer4[7][31:24] <= buffer_data_0[95:88];
        layer4[7][39:32] <= buffer_data_0[103:96];
        layer0[8][7:0] <= buffer_data_4[79:72];
        layer0[8][15:8] <= buffer_data_4[87:80];
        layer0[8][23:16] <= buffer_data_4[95:88];
        layer0[8][31:24] <= buffer_data_4[103:96];
        layer0[8][39:32] <= buffer_data_4[111:104];
        layer1[8][7:0] <= buffer_data_3[79:72];
        layer1[8][15:8] <= buffer_data_3[87:80];
        layer1[8][23:16] <= buffer_data_3[95:88];
        layer1[8][31:24] <= buffer_data_3[103:96];
        layer1[8][39:32] <= buffer_data_3[111:104];
        layer2[8][7:0] <= buffer_data_2[79:72];
        layer2[8][15:8] <= buffer_data_2[87:80];
        layer2[8][23:16] <= buffer_data_2[95:88];
        layer2[8][31:24] <= buffer_data_2[103:96];
        layer2[8][39:32] <= buffer_data_2[111:104];
        layer3[8][7:0] <= buffer_data_1[79:72];
        layer3[8][15:8] <= buffer_data_1[87:80];
        layer3[8][23:16] <= buffer_data_1[95:88];
        layer3[8][31:24] <= buffer_data_1[103:96];
        layer3[8][39:32] <= buffer_data_1[111:104];
        layer4[8][7:0] <= buffer_data_0[79:72];
        layer4[8][15:8] <= buffer_data_0[87:80];
        layer4[8][23:16] <= buffer_data_0[95:88];
        layer4[8][31:24] <= buffer_data_0[103:96];
        layer4[8][39:32] <= buffer_data_0[111:104];
        layer0[9][7:0] <= buffer_data_4[87:80];
        layer0[9][15:8] <= buffer_data_4[95:88];
        layer0[9][23:16] <= buffer_data_4[103:96];
        layer0[9][31:24] <= buffer_data_4[111:104];
        layer0[9][39:32] <= buffer_data_4[119:112];
        layer1[9][7:0] <= buffer_data_3[87:80];
        layer1[9][15:8] <= buffer_data_3[95:88];
        layer1[9][23:16] <= buffer_data_3[103:96];
        layer1[9][31:24] <= buffer_data_3[111:104];
        layer1[9][39:32] <= buffer_data_3[119:112];
        layer2[9][7:0] <= buffer_data_2[87:80];
        layer2[9][15:8] <= buffer_data_2[95:88];
        layer2[9][23:16] <= buffer_data_2[103:96];
        layer2[9][31:24] <= buffer_data_2[111:104];
        layer2[9][39:32] <= buffer_data_2[119:112];
        layer3[9][7:0] <= buffer_data_1[87:80];
        layer3[9][15:8] <= buffer_data_1[95:88];
        layer3[9][23:16] <= buffer_data_1[103:96];
        layer3[9][31:24] <= buffer_data_1[111:104];
        layer3[9][39:32] <= buffer_data_1[119:112];
        layer4[9][7:0] <= buffer_data_0[87:80];
        layer4[9][15:8] <= buffer_data_0[95:88];
        layer4[9][23:16] <= buffer_data_0[103:96];
        layer4[9][31:24] <= buffer_data_0[111:104];
        layer4[9][39:32] <= buffer_data_0[119:112];
        layer0[10][7:0] <= buffer_data_4[95:88];
        layer0[10][15:8] <= buffer_data_4[103:96];
        layer0[10][23:16] <= buffer_data_4[111:104];
        layer0[10][31:24] <= buffer_data_4[119:112];
        layer0[10][39:32] <= buffer_data_4[127:120];
        layer1[10][7:0] <= buffer_data_3[95:88];
        layer1[10][15:8] <= buffer_data_3[103:96];
        layer1[10][23:16] <= buffer_data_3[111:104];
        layer1[10][31:24] <= buffer_data_3[119:112];
        layer1[10][39:32] <= buffer_data_3[127:120];
        layer2[10][7:0] <= buffer_data_2[95:88];
        layer2[10][15:8] <= buffer_data_2[103:96];
        layer2[10][23:16] <= buffer_data_2[111:104];
        layer2[10][31:24] <= buffer_data_2[119:112];
        layer2[10][39:32] <= buffer_data_2[127:120];
        layer3[10][7:0] <= buffer_data_1[95:88];
        layer3[10][15:8] <= buffer_data_1[103:96];
        layer3[10][23:16] <= buffer_data_1[111:104];
        layer3[10][31:24] <= buffer_data_1[119:112];
        layer3[10][39:32] <= buffer_data_1[127:120];
        layer4[10][7:0] <= buffer_data_0[95:88];
        layer4[10][15:8] <= buffer_data_0[103:96];
        layer4[10][23:16] <= buffer_data_0[111:104];
        layer4[10][31:24] <= buffer_data_0[119:112];
        layer4[10][39:32] <= buffer_data_0[127:120];
        layer0[11][7:0] <= buffer_data_4[103:96];
        layer0[11][15:8] <= buffer_data_4[111:104];
        layer0[11][23:16] <= buffer_data_4[119:112];
        layer0[11][31:24] <= buffer_data_4[127:120];
        layer0[11][39:32] <= buffer_data_4[135:128];
        layer1[11][7:0] <= buffer_data_3[103:96];
        layer1[11][15:8] <= buffer_data_3[111:104];
        layer1[11][23:16] <= buffer_data_3[119:112];
        layer1[11][31:24] <= buffer_data_3[127:120];
        layer1[11][39:32] <= buffer_data_3[135:128];
        layer2[11][7:0] <= buffer_data_2[103:96];
        layer2[11][15:8] <= buffer_data_2[111:104];
        layer2[11][23:16] <= buffer_data_2[119:112];
        layer2[11][31:24] <= buffer_data_2[127:120];
        layer2[11][39:32] <= buffer_data_2[135:128];
        layer3[11][7:0] <= buffer_data_1[103:96];
        layer3[11][15:8] <= buffer_data_1[111:104];
        layer3[11][23:16] <= buffer_data_1[119:112];
        layer3[11][31:24] <= buffer_data_1[127:120];
        layer3[11][39:32] <= buffer_data_1[135:128];
        layer4[11][7:0] <= buffer_data_0[103:96];
        layer4[11][15:8] <= buffer_data_0[111:104];
        layer4[11][23:16] <= buffer_data_0[119:112];
        layer4[11][31:24] <= buffer_data_0[127:120];
        layer4[11][39:32] <= buffer_data_0[135:128];
        layer0[12][7:0] <= buffer_data_4[111:104];
        layer0[12][15:8] <= buffer_data_4[119:112];
        layer0[12][23:16] <= buffer_data_4[127:120];
        layer0[12][31:24] <= buffer_data_4[135:128];
        layer0[12][39:32] <= buffer_data_4[143:136];
        layer1[12][7:0] <= buffer_data_3[111:104];
        layer1[12][15:8] <= buffer_data_3[119:112];
        layer1[12][23:16] <= buffer_data_3[127:120];
        layer1[12][31:24] <= buffer_data_3[135:128];
        layer1[12][39:32] <= buffer_data_3[143:136];
        layer2[12][7:0] <= buffer_data_2[111:104];
        layer2[12][15:8] <= buffer_data_2[119:112];
        layer2[12][23:16] <= buffer_data_2[127:120];
        layer2[12][31:24] <= buffer_data_2[135:128];
        layer2[12][39:32] <= buffer_data_2[143:136];
        layer3[12][7:0] <= buffer_data_1[111:104];
        layer3[12][15:8] <= buffer_data_1[119:112];
        layer3[12][23:16] <= buffer_data_1[127:120];
        layer3[12][31:24] <= buffer_data_1[135:128];
        layer3[12][39:32] <= buffer_data_1[143:136];
        layer4[12][7:0] <= buffer_data_0[111:104];
        layer4[12][15:8] <= buffer_data_0[119:112];
        layer4[12][23:16] <= buffer_data_0[127:120];
        layer4[12][31:24] <= buffer_data_0[135:128];
        layer4[12][39:32] <= buffer_data_0[143:136];
        layer0[13][7:0] <= buffer_data_4[119:112];
        layer0[13][15:8] <= buffer_data_4[127:120];
        layer0[13][23:16] <= buffer_data_4[135:128];
        layer0[13][31:24] <= buffer_data_4[143:136];
        layer0[13][39:32] <= buffer_data_4[151:144];
        layer1[13][7:0] <= buffer_data_3[119:112];
        layer1[13][15:8] <= buffer_data_3[127:120];
        layer1[13][23:16] <= buffer_data_3[135:128];
        layer1[13][31:24] <= buffer_data_3[143:136];
        layer1[13][39:32] <= buffer_data_3[151:144];
        layer2[13][7:0] <= buffer_data_2[119:112];
        layer2[13][15:8] <= buffer_data_2[127:120];
        layer2[13][23:16] <= buffer_data_2[135:128];
        layer2[13][31:24] <= buffer_data_2[143:136];
        layer2[13][39:32] <= buffer_data_2[151:144];
        layer3[13][7:0] <= buffer_data_1[119:112];
        layer3[13][15:8] <= buffer_data_1[127:120];
        layer3[13][23:16] <= buffer_data_1[135:128];
        layer3[13][31:24] <= buffer_data_1[143:136];
        layer3[13][39:32] <= buffer_data_1[151:144];
        layer4[13][7:0] <= buffer_data_0[119:112];
        layer4[13][15:8] <= buffer_data_0[127:120];
        layer4[13][23:16] <= buffer_data_0[135:128];
        layer4[13][31:24] <= buffer_data_0[143:136];
        layer4[13][39:32] <= buffer_data_0[151:144];
        layer0[14][7:0] <= buffer_data_4[127:120];
        layer0[14][15:8] <= buffer_data_4[135:128];
        layer0[14][23:16] <= buffer_data_4[143:136];
        layer0[14][31:24] <= buffer_data_4[151:144];
        layer0[14][39:32] <= 0;
        layer1[14][7:0] <= buffer_data_3[127:120];
        layer1[14][15:8] <= buffer_data_3[135:128];
        layer1[14][23:16] <= buffer_data_3[143:136];
        layer1[14][31:24] <= buffer_data_3[151:144];
        layer1[14][39:32] <= 0;
        layer2[14][7:0] <= buffer_data_2[127:120];
        layer2[14][15:8] <= buffer_data_2[135:128];
        layer2[14][23:16] <= buffer_data_2[143:136];
        layer2[14][31:24] <= buffer_data_2[151:144];
        layer2[14][39:32] <= 0;
        layer3[14][7:0] <= buffer_data_1[127:120];
        layer3[14][15:8] <= buffer_data_1[135:128];
        layer3[14][23:16] <= buffer_data_1[143:136];
        layer3[14][31:24] <= buffer_data_1[151:144];
        layer3[14][39:32] <= 0;
        layer4[14][7:0] <= buffer_data_0[127:120];
        layer4[14][15:8] <= buffer_data_0[135:128];
        layer4[14][23:16] <= buffer_data_0[143:136];
        layer4[14][31:24] <= buffer_data_0[151:144];
        layer4[14][39:32] <= 0;
        layer0[15][7:0] <= buffer_data_4[135:128];
        layer0[15][15:8] <= buffer_data_4[143:136];
        layer0[15][23:16] <= buffer_data_4[151:144];
        layer0[15][31:24] <= 0;
        layer0[15][39:32] <= 0;
        layer1[15][7:0] <= buffer_data_3[135:128];
        layer1[15][15:8] <= buffer_data_3[143:136];
        layer1[15][23:16] <= buffer_data_3[151:144];
        layer1[15][31:24] <= 0;
        layer1[15][39:32] <= 0;
        layer2[15][7:0] <= buffer_data_2[135:128];
        layer2[15][15:8] <= buffer_data_2[143:136];
        layer2[15][23:16] <= buffer_data_2[151:144];
        layer2[15][31:24] <= 0;
        layer2[15][39:32] <= 0;
        layer3[15][7:0] <= buffer_data_1[135:128];
        layer3[15][15:8] <= buffer_data_1[143:136];
        layer3[15][23:16] <= buffer_data_1[151:144];
        layer3[15][31:24] <= 0;
        layer3[15][39:32] <= 0;
        layer4[15][7:0] <= buffer_data_0[135:128];
        layer4[15][15:8] <= buffer_data_0[143:136];
        layer4[15][23:16] <= buffer_data_0[151:144];
        layer4[15][31:24] <= 0;
        layer4[15][39:32] <= 0;
    end
      default: begin
        layer0[0][7:0] <= 'd0;
        layer0[0][15:8] <= 'd0;
        layer0[0][23:16] <= 'd0;
        layer0[0][31:24] <= 'd0;
        layer0[0][39:32] <= 'd0;
        layer1[0][7:0] <= 'd0;
        layer1[0][15:8] <= 'd0;
        layer1[0][23:16] <= 'd0;
        layer1[0][31:24] <= 'd0;
        layer1[0][39:32] <= 'd0;
        layer2[0][7:0] <= 'd0;
        layer2[0][15:8] <= 'd0;
        layer2[0][23:16] <= 'd0;
        layer2[0][31:24] <= 'd0;
        layer2[0][39:32] <= 'd0;
        layer3[0][7:0] <= 'd0;
        layer3[0][15:8] <= 'd0;
        layer3[0][23:16] <= 'd0;
        layer3[0][31:24] <= 'd0;
        layer3[0][39:32] <= 'd0;
        layer4[0][7:0] <= 'd0;
        layer4[0][15:8] <= 'd0;
        layer4[0][23:16] <= 'd0;
        layer4[0][31:24] <= 'd0;
        layer4[0][39:32] <= 'd0;
        layer0[1][7:0] <= 'd0;
        layer0[1][15:8] <= 'd0;
        layer0[1][23:16] <= 'd0;
        layer0[1][31:24] <= 'd0;
        layer0[1][39:32] <= 'd0;
        layer1[1][7:0] <= 'd0;
        layer1[1][15:8] <= 'd0;
        layer1[1][23:16] <= 'd0;
        layer1[1][31:24] <= 'd0;
        layer1[1][39:32] <= 'd0;
        layer2[1][7:0] <= 'd0;
        layer2[1][15:8] <= 'd0;
        layer2[1][23:16] <= 'd0;
        layer2[1][31:24] <= 'd0;
        layer2[1][39:32] <= 'd0;
        layer3[1][7:0] <= 'd0;
        layer3[1][15:8] <= 'd0;
        layer3[1][23:16] <= 'd0;
        layer3[1][31:24] <= 'd0;
        layer3[1][39:32] <= 'd0;
        layer4[1][7:0] <= 'd0;
        layer4[1][15:8] <= 'd0;
        layer4[1][23:16] <= 'd0;
        layer4[1][31:24] <= 'd0;
        layer4[1][39:32] <= 'd0;
        layer0[2][7:0] <= 'd0;
        layer0[2][15:8] <= 'd0;
        layer0[2][23:16] <= 'd0;
        layer0[2][31:24] <= 'd0;
        layer0[2][39:32] <= 'd0;
        layer1[2][7:0] <= 'd0;
        layer1[2][15:8] <= 'd0;
        layer1[2][23:16] <= 'd0;
        layer1[2][31:24] <= 'd0;
        layer1[2][39:32] <= 'd0;
        layer2[2][7:0] <= 'd0;
        layer2[2][15:8] <= 'd0;
        layer2[2][23:16] <= 'd0;
        layer2[2][31:24] <= 'd0;
        layer2[2][39:32] <= 'd0;
        layer3[2][7:0] <= 'd0;
        layer3[2][15:8] <= 'd0;
        layer3[2][23:16] <= 'd0;
        layer3[2][31:24] <= 'd0;
        layer3[2][39:32] <= 'd0;
        layer4[2][7:0] <= 'd0;
        layer4[2][15:8] <= 'd0;
        layer4[2][23:16] <= 'd0;
        layer4[2][31:24] <= 'd0;
        layer4[2][39:32] <= 'd0;
        layer0[3][7:0] <= 'd0;
        layer0[3][15:8] <= 'd0;
        layer0[3][23:16] <= 'd0;
        layer0[3][31:24] <= 'd0;
        layer0[3][39:32] <= 'd0;
        layer1[3][7:0] <= 'd0;
        layer1[3][15:8] <= 'd0;
        layer1[3][23:16] <= 'd0;
        layer1[3][31:24] <= 'd0;
        layer1[3][39:32] <= 'd0;
        layer2[3][7:0] <= 'd0;
        layer2[3][15:8] <= 'd0;
        layer2[3][23:16] <= 'd0;
        layer2[3][31:24] <= 'd0;
        layer2[3][39:32] <= 'd0;
        layer3[3][7:0] <= 'd0;
        layer3[3][15:8] <= 'd0;
        layer3[3][23:16] <= 'd0;
        layer3[3][31:24] <= 'd0;
        layer3[3][39:32] <= 'd0;
        layer4[3][7:0] <= 'd0;
        layer4[3][15:8] <= 'd0;
        layer4[3][23:16] <= 'd0;
        layer4[3][31:24] <= 'd0;
        layer4[3][39:32] <= 'd0;
        layer0[4][7:0] <= 'd0;
        layer0[4][15:8] <= 'd0;
        layer0[4][23:16] <= 'd0;
        layer0[4][31:24] <= 'd0;
        layer0[4][39:32] <= 'd0;
        layer1[4][7:0] <= 'd0;
        layer1[4][15:8] <= 'd0;
        layer1[4][23:16] <= 'd0;
        layer1[4][31:24] <= 'd0;
        layer1[4][39:32] <= 'd0;
        layer2[4][7:0] <= 'd0;
        layer2[4][15:8] <= 'd0;
        layer2[4][23:16] <= 'd0;
        layer2[4][31:24] <= 'd0;
        layer2[4][39:32] <= 'd0;
        layer3[4][7:0] <= 'd0;
        layer3[4][15:8] <= 'd0;
        layer3[4][23:16] <= 'd0;
        layer3[4][31:24] <= 'd0;
        layer3[4][39:32] <= 'd0;
        layer4[4][7:0] <= 'd0;
        layer4[4][15:8] <= 'd0;
        layer4[4][23:16] <= 'd0;
        layer4[4][31:24] <= 'd0;
        layer4[4][39:32] <= 'd0;
        layer0[5][7:0] <= 'd0;
        layer0[5][15:8] <= 'd0;
        layer0[5][23:16] <= 'd0;
        layer0[5][31:24] <= 'd0;
        layer0[5][39:32] <= 'd0;
        layer1[5][7:0] <= 'd0;
        layer1[5][15:8] <= 'd0;
        layer1[5][23:16] <= 'd0;
        layer1[5][31:24] <= 'd0;
        layer1[5][39:32] <= 'd0;
        layer2[5][7:0] <= 'd0;
        layer2[5][15:8] <= 'd0;
        layer2[5][23:16] <= 'd0;
        layer2[5][31:24] <= 'd0;
        layer2[5][39:32] <= 'd0;
        layer3[5][7:0] <= 'd0;
        layer3[5][15:8] <= 'd0;
        layer3[5][23:16] <= 'd0;
        layer3[5][31:24] <= 'd0;
        layer3[5][39:32] <= 'd0;
        layer4[5][7:0] <= 'd0;
        layer4[5][15:8] <= 'd0;
        layer4[5][23:16] <= 'd0;
        layer4[5][31:24] <= 'd0;
        layer4[5][39:32] <= 'd0;
        layer0[6][7:0] <= 'd0;
        layer0[6][15:8] <= 'd0;
        layer0[6][23:16] <= 'd0;
        layer0[6][31:24] <= 'd0;
        layer0[6][39:32] <= 'd0;
        layer1[6][7:0] <= 'd0;
        layer1[6][15:8] <= 'd0;
        layer1[6][23:16] <= 'd0;
        layer1[6][31:24] <= 'd0;
        layer1[6][39:32] <= 'd0;
        layer2[6][7:0] <= 'd0;
        layer2[6][15:8] <= 'd0;
        layer2[6][23:16] <= 'd0;
        layer2[6][31:24] <= 'd0;
        layer2[6][39:32] <= 'd0;
        layer3[6][7:0] <= 'd0;
        layer3[6][15:8] <= 'd0;
        layer3[6][23:16] <= 'd0;
        layer3[6][31:24] <= 'd0;
        layer3[6][39:32] <= 'd0;
        layer4[6][7:0] <= 'd0;
        layer4[6][15:8] <= 'd0;
        layer4[6][23:16] <= 'd0;
        layer4[6][31:24] <= 'd0;
        layer4[6][39:32] <= 'd0;
        layer0[7][7:0] <= 'd0;
        layer0[7][15:8] <= 'd0;
        layer0[7][23:16] <= 'd0;
        layer0[7][31:24] <= 'd0;
        layer0[7][39:32] <= 'd0;
        layer1[7][7:0] <= 'd0;
        layer1[7][15:8] <= 'd0;
        layer1[7][23:16] <= 'd0;
        layer1[7][31:24] <= 'd0;
        layer1[7][39:32] <= 'd0;
        layer2[7][7:0] <= 'd0;
        layer2[7][15:8] <= 'd0;
        layer2[7][23:16] <= 'd0;
        layer2[7][31:24] <= 'd0;
        layer2[7][39:32] <= 'd0;
        layer3[7][7:0] <= 'd0;
        layer3[7][15:8] <= 'd0;
        layer3[7][23:16] <= 'd0;
        layer3[7][31:24] <= 'd0;
        layer3[7][39:32] <= 'd0;
        layer4[7][7:0] <= 'd0;
        layer4[7][15:8] <= 'd0;
        layer4[7][23:16] <= 'd0;
        layer4[7][31:24] <= 'd0;
        layer4[7][39:32] <= 'd0;
        layer0[8][7:0] <= 'd0;
        layer0[8][15:8] <= 'd0;
        layer0[8][23:16] <= 'd0;
        layer0[8][31:24] <= 'd0;
        layer0[8][39:32] <= 'd0;
        layer1[8][7:0] <= 'd0;
        layer1[8][15:8] <= 'd0;
        layer1[8][23:16] <= 'd0;
        layer1[8][31:24] <= 'd0;
        layer1[8][39:32] <= 'd0;
        layer2[8][7:0] <= 'd0;
        layer2[8][15:8] <= 'd0;
        layer2[8][23:16] <= 'd0;
        layer2[8][31:24] <= 'd0;
        layer2[8][39:32] <= 'd0;
        layer3[8][7:0] <= 'd0;
        layer3[8][15:8] <= 'd0;
        layer3[8][23:16] <= 'd0;
        layer3[8][31:24] <= 'd0;
        layer3[8][39:32] <= 'd0;
        layer4[8][7:0] <= 'd0;
        layer4[8][15:8] <= 'd0;
        layer4[8][23:16] <= 'd0;
        layer4[8][31:24] <= 'd0;
        layer4[8][39:32] <= 'd0;
        layer0[9][7:0] <= 'd0;
        layer0[9][15:8] <= 'd0;
        layer0[9][23:16] <= 'd0;
        layer0[9][31:24] <= 'd0;
        layer0[9][39:32] <= 'd0;
        layer1[9][7:0] <= 'd0;
        layer1[9][15:8] <= 'd0;
        layer1[9][23:16] <= 'd0;
        layer1[9][31:24] <= 'd0;
        layer1[9][39:32] <= 'd0;
        layer2[9][7:0] <= 'd0;
        layer2[9][15:8] <= 'd0;
        layer2[9][23:16] <= 'd0;
        layer2[9][31:24] <= 'd0;
        layer2[9][39:32] <= 'd0;
        layer3[9][7:0] <= 'd0;
        layer3[9][15:8] <= 'd0;
        layer3[9][23:16] <= 'd0;
        layer3[9][31:24] <= 'd0;
        layer3[9][39:32] <= 'd0;
        layer4[9][7:0] <= 'd0;
        layer4[9][15:8] <= 'd0;
        layer4[9][23:16] <= 'd0;
        layer4[9][31:24] <= 'd0;
        layer4[9][39:32] <= 'd0;
        layer0[10][7:0] <= 'd0;
        layer0[10][15:8] <= 'd0;
        layer0[10][23:16] <= 'd0;
        layer0[10][31:24] <= 'd0;
        layer0[10][39:32] <= 'd0;
        layer1[10][7:0] <= 'd0;
        layer1[10][15:8] <= 'd0;
        layer1[10][23:16] <= 'd0;
        layer1[10][31:24] <= 'd0;
        layer1[10][39:32] <= 'd0;
        layer2[10][7:0] <= 'd0;
        layer2[10][15:8] <= 'd0;
        layer2[10][23:16] <= 'd0;
        layer2[10][31:24] <= 'd0;
        layer2[10][39:32] <= 'd0;
        layer3[10][7:0] <= 'd0;
        layer3[10][15:8] <= 'd0;
        layer3[10][23:16] <= 'd0;
        layer3[10][31:24] <= 'd0;
        layer3[10][39:32] <= 'd0;
        layer4[10][7:0] <= 'd0;
        layer4[10][15:8] <= 'd0;
        layer4[10][23:16] <= 'd0;
        layer4[10][31:24] <= 'd0;
        layer4[10][39:32] <= 'd0;
        layer0[11][7:0] <= 'd0;
        layer0[11][15:8] <= 'd0;
        layer0[11][23:16] <= 'd0;
        layer0[11][31:24] <= 'd0;
        layer0[11][39:32] <= 'd0;
        layer1[11][7:0] <= 'd0;
        layer1[11][15:8] <= 'd0;
        layer1[11][23:16] <= 'd0;
        layer1[11][31:24] <= 'd0;
        layer1[11][39:32] <= 'd0;
        layer2[11][7:0] <= 'd0;
        layer2[11][15:8] <= 'd0;
        layer2[11][23:16] <= 'd0;
        layer2[11][31:24] <= 'd0;
        layer2[11][39:32] <= 'd0;
        layer3[11][7:0] <= 'd0;
        layer3[11][15:8] <= 'd0;
        layer3[11][23:16] <= 'd0;
        layer3[11][31:24] <= 'd0;
        layer3[11][39:32] <= 'd0;
        layer4[11][7:0] <= 'd0;
        layer4[11][15:8] <= 'd0;
        layer4[11][23:16] <= 'd0;
        layer4[11][31:24] <= 'd0;
        layer4[11][39:32] <= 'd0;
        layer0[12][7:0] <= 'd0;
        layer0[12][15:8] <= 'd0;
        layer0[12][23:16] <= 'd0;
        layer0[12][31:24] <= 'd0;
        layer0[12][39:32] <= 'd0;
        layer1[12][7:0] <= 'd0;
        layer1[12][15:8] <= 'd0;
        layer1[12][23:16] <= 'd0;
        layer1[12][31:24] <= 'd0;
        layer1[12][39:32] <= 'd0;
        layer2[12][7:0] <= 'd0;
        layer2[12][15:8] <= 'd0;
        layer2[12][23:16] <= 'd0;
        layer2[12][31:24] <= 'd0;
        layer2[12][39:32] <= 'd0;
        layer3[12][7:0] <= 'd0;
        layer3[12][15:8] <= 'd0;
        layer3[12][23:16] <= 'd0;
        layer3[12][31:24] <= 'd0;
        layer3[12][39:32] <= 'd0;
        layer4[12][7:0] <= 'd0;
        layer4[12][15:8] <= 'd0;
        layer4[12][23:16] <= 'd0;
        layer4[12][31:24] <= 'd0;
        layer4[12][39:32] <= 'd0;
        layer0[13][7:0] <= 'd0;
        layer0[13][15:8] <= 'd0;
        layer0[13][23:16] <= 'd0;
        layer0[13][31:24] <= 'd0;
        layer0[13][39:32] <= 'd0;
        layer1[13][7:0] <= 'd0;
        layer1[13][15:8] <= 'd0;
        layer1[13][23:16] <= 'd0;
        layer1[13][31:24] <= 'd0;
        layer1[13][39:32] <= 'd0;
        layer2[13][7:0] <= 'd0;
        layer2[13][15:8] <= 'd0;
        layer2[13][23:16] <= 'd0;
        layer2[13][31:24] <= 'd0;
        layer2[13][39:32] <= 'd0;
        layer3[13][7:0] <= 'd0;
        layer3[13][15:8] <= 'd0;
        layer3[13][23:16] <= 'd0;
        layer3[13][31:24] <= 'd0;
        layer3[13][39:32] <= 'd0;
        layer4[13][7:0] <= 'd0;
        layer4[13][15:8] <= 'd0;
        layer4[13][23:16] <= 'd0;
        layer4[13][31:24] <= 'd0;
        layer4[13][39:32] <= 'd0;
        layer0[14][7:0] <= 'd0;
        layer0[14][15:8] <= 'd0;
        layer0[14][23:16] <= 'd0;
        layer0[14][31:24] <= 'd0;
        layer0[14][39:32] <= 'd0;
        layer1[14][7:0] <= 'd0;
        layer1[14][15:8] <= 'd0;
        layer1[14][23:16] <= 'd0;
        layer1[14][31:24] <= 'd0;
        layer1[14][39:32] <= 'd0;
        layer2[14][7:0] <= 'd0;
        layer2[14][15:8] <= 'd0;
        layer2[14][23:16] <= 'd0;
        layer2[14][31:24] <= 'd0;
        layer2[14][39:32] <= 'd0;
        layer3[14][7:0] <= 'd0;
        layer3[14][15:8] <= 'd0;
        layer3[14][23:16] <= 'd0;
        layer3[14][31:24] <= 'd0;
        layer3[14][39:32] <= 'd0;
        layer4[14][7:0] <= 'd0;
        layer4[14][15:8] <= 'd0;
        layer4[14][23:16] <= 'd0;
        layer4[14][31:24] <= 'd0;
        layer4[14][39:32] <= 'd0;
        layer0[15][7:0] <= 'd0;
        layer0[15][15:8] <= 'd0;
        layer0[15][23:16] <= 'd0;
        layer0[15][31:24] <= 'd0;
        layer0[15][39:32] <= 'd0;
        layer1[15][7:0] <= 'd0;
        layer1[15][15:8] <= 'd0;
        layer1[15][23:16] <= 'd0;
        layer1[15][31:24] <= 'd0;
        layer1[15][39:32] <= 'd0;
        layer2[15][7:0] <= 'd0;
        layer2[15][15:8] <= 'd0;
        layer2[15][23:16] <= 'd0;
        layer2[15][31:24] <= 'd0;
        layer2[15][39:32] <= 'd0;
        layer3[15][7:0] <= 'd0;
        layer3[15][15:8] <= 'd0;
        layer3[15][23:16] <= 'd0;
        layer3[15][31:24] <= 'd0;
        layer3[15][39:32] <= 'd0;
        layer4[15][7:0] <= 'd0;
        layer4[15][15:8] <= 'd0;
        layer4[15][23:16] <= 'd0;
        layer4[15][31:24] <= 'd0;
        layer4[15][39:32] <= 'd0;
      end
    endcase
  end
end

reg  [15:0]  kernel_img_mul_0[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_0[0] <= 'd0;
    kernel_img_mul_0[1] <= 'd0;
    kernel_img_mul_0[2] <= 'd0;
    kernel_img_mul_0[3] <= 'd0;
    kernel_img_mul_0[4] <= 'd0;
    kernel_img_mul_0[5] <= 'd0;
    kernel_img_mul_0[6] <= 'd0;
    kernel_img_mul_0[7] <= 'd0;
    kernel_img_mul_0[8] <= 'd0;
    kernel_img_mul_0[9] <= 'd0;
    kernel_img_mul_0[10] <= 'd0;
    kernel_img_mul_0[11] <= 'd0;
    kernel_img_mul_0[12] <= 'd0;
    kernel_img_mul_0[13] <= 'd0;
    kernel_img_mul_0[14] <= 'd0;
    kernel_img_mul_0[15] <= 'd0;
    kernel_img_mul_0[16] <= 'd0;
    kernel_img_mul_0[17] <= 'd0;
    kernel_img_mul_0[18] <= 'd0;
    kernel_img_mul_0[19] <= 'd0;
    kernel_img_mul_0[20] <= 'd0;
    kernel_img_mul_0[21] <= 'd0;
    kernel_img_mul_0[22] <= 'd0;
    kernel_img_mul_0[23] <= 'd0;
    kernel_img_mul_0[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_0[0] <= { {8{1'b0}},layer0[0][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_0[1] <= { {8{1'b0}},layer0[0][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_0[2] <= { {8{1'b0}},layer0[0][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_0[3] <= { {8{1'b0}},layer0[0][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_0[4] <= { {8{1'b0}},layer0[0][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_0[5] <= { {8{1'b0}},layer1[0][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_0[6] <= { {8{1'b0}},layer1[0][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_0[7] <= { {8{1'b0}},layer1[0][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_0[8] <= { {8{1'b0}},layer1[0][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_0[9] <= { {8{1'b0}},layer1[0][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_0[10] <= { {8{1'b0}},layer2[0][7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_0[11] <= { {8{1'b0}},layer2[0][15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_0[12] <= { {8{1'b0}},layer2[0][23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_0[13] <= { {8{1'b0}},layer2[0][31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_0[14] <= { {8{1'b0}},layer2[0][39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_0[15] <= { {8{1'b0}},layer3[0][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_0[16] <= { {8{1'b0}},layer3[0][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_0[17] <= { {8{1'b0}},layer3[0][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_0[18] <= { {8{1'b0}},layer3[0][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_0[19] <= { {8{1'b0}},layer3[0][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_0[20] <= { {8{1'b0}},layer4[0][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_0[21] <= { {8{1'b0}},layer4[0][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_0[22] <= { {8{1'b0}},layer4[0][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_0[23] <= { {8{1'b0}},layer4[0][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_0[24] <= { {8{1'b0}},layer4[0][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_0;
reg  [15:0]  kernel_img_sum_2_0;
reg  [15:0]  kernel_img_sum_3_0;
reg  [15:0]  kernel_img_sum_4_0;
reg  [15:0]  kernel_img_sum_5_0;
reg  [15:0]  kernel_img_sum_6_0;
reg  [15:0]  kernel_img_sum_7_0;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_0 <= kernel_img_mul_0[0] + kernel_img_mul_0[1] + kernel_img_mul_0[2] + kernel_img_mul_0[3] + kernel_img_mul_0[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_0 <= kernel_img_mul_0[5] + kernel_img_mul_0[6] + kernel_img_mul_0[7] + kernel_img_mul_0[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_0 <= kernel_img_mul_0[9] + kernel_img_mul_0[10] + kernel_img_mul_0[11] + kernel_img_mul_0[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_0 <= kernel_img_mul_0[13] + kernel_img_mul_0[14] + kernel_img_mul_0[15] + kernel_img_mul_0[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_0 <= kernel_img_mul_0[17] + kernel_img_mul_0[18] + kernel_img_mul_0[19] + kernel_img_mul_0[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_0 <= kernel_img_mul_0[21] + kernel_img_mul_0[22] + kernel_img_mul_0[23] + kernel_img_mul_0[24];
  end
end
always@(*) begin
  kernel_img_sum_7_0 = kernel_img_sum_1_0 + kernel_img_sum_2_0 + kernel_img_sum_3_0 + kernel_img_sum_4_0 + kernel_img_sum_5_0 + kernel_img_sum_6_0;
end
reg  [15:0]  kernel_img_mul_1[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_1[0] <= 'd0;
    kernel_img_mul_1[1] <= 'd0;
    kernel_img_mul_1[2] <= 'd0;
    kernel_img_mul_1[3] <= 'd0;
    kernel_img_mul_1[4] <= 'd0;
    kernel_img_mul_1[5] <= 'd0;
    kernel_img_mul_1[6] <= 'd0;
    kernel_img_mul_1[7] <= 'd0;
    kernel_img_mul_1[8] <= 'd0;
    kernel_img_mul_1[9] <= 'd0;
    kernel_img_mul_1[10] <= 'd0;
    kernel_img_mul_1[11] <= 'd0;
    kernel_img_mul_1[12] <= 'd0;
    kernel_img_mul_1[13] <= 'd0;
    kernel_img_mul_1[14] <= 'd0;
    kernel_img_mul_1[15] <= 'd0;
    kernel_img_mul_1[16] <= 'd0;
    kernel_img_mul_1[17] <= 'd0;
    kernel_img_mul_1[18] <= 'd0;
    kernel_img_mul_1[19] <= 'd0;
    kernel_img_mul_1[20] <= 'd0;
    kernel_img_mul_1[21] <= 'd0;
    kernel_img_mul_1[22] <= 'd0;
    kernel_img_mul_1[23] <= 'd0;
    kernel_img_mul_1[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_1[0] <= { {8{1'b0}},layer0[1][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_1[1] <= { {8{1'b0}},layer0[1][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_1[2] <= { {8{1'b0}},layer0[1][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_1[3] <= { {8{1'b0}},layer0[1][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_1[4] <= { {8{1'b0}},layer0[1][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_1[5] <= { {8{1'b0}},layer1[1][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_1[6] <= { {8{1'b0}},layer1[1][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_1[7] <= { {8{1'b0}},layer1[1][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_1[8] <= { {8{1'b0}},layer1[1][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_1[9] <= { {8{1'b0}},layer1[1][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_1[10] <= { {8{1'b0}},layer2[1][7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_1[11] <= { {8{1'b0}},layer2[1][15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_1[12] <= { {8{1'b0}},layer2[1][23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_1[13] <= { {8{1'b0}},layer2[1][31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_1[14] <= { {8{1'b0}},layer2[1][39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_1[15] <= { {8{1'b0}},layer3[1][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_1[16] <= { {8{1'b0}},layer3[1][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_1[17] <= { {8{1'b0}},layer3[1][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_1[18] <= { {8{1'b0}},layer3[1][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_1[19] <= { {8{1'b0}},layer3[1][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_1[20] <= { {8{1'b0}},layer4[1][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_1[21] <= { {8{1'b0}},layer4[1][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_1[22] <= { {8{1'b0}},layer4[1][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_1[23] <= { {8{1'b0}},layer4[1][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_1[24] <= { {8{1'b0}},layer4[1][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_1;
reg  [15:0]  kernel_img_sum_2_1;
reg  [15:0]  kernel_img_sum_3_1;
reg  [15:0]  kernel_img_sum_4_1;
reg  [15:0]  kernel_img_sum_5_1;
reg  [15:0]  kernel_img_sum_6_1;
reg  [15:0]  kernel_img_sum_7_1;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_1 <= kernel_img_mul_1[0] + kernel_img_mul_1[1] + kernel_img_mul_1[2] + kernel_img_mul_1[3] + kernel_img_mul_1[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_1 <= kernel_img_mul_1[5] + kernel_img_mul_1[6] + kernel_img_mul_1[7] + kernel_img_mul_1[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_1 <= kernel_img_mul_1[9] + kernel_img_mul_1[10] + kernel_img_mul_1[11] + kernel_img_mul_1[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_1 <= kernel_img_mul_1[13] + kernel_img_mul_1[14] + kernel_img_mul_1[15] + kernel_img_mul_1[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_1 <= kernel_img_mul_1[17] + kernel_img_mul_1[18] + kernel_img_mul_1[19] + kernel_img_mul_1[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_1 <= kernel_img_mul_1[21] + kernel_img_mul_1[22] + kernel_img_mul_1[23] + kernel_img_mul_1[24];
  end
end
always@(*) begin
  kernel_img_sum_7_1 = kernel_img_sum_1_1 + kernel_img_sum_2_1 + kernel_img_sum_3_1 + kernel_img_sum_4_1 + kernel_img_sum_5_1 + kernel_img_sum_6_1;
end
reg  [15:0]  kernel_img_mul_2[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_2[0] <= 'd0;
    kernel_img_mul_2[1] <= 'd0;
    kernel_img_mul_2[2] <= 'd0;
    kernel_img_mul_2[3] <= 'd0;
    kernel_img_mul_2[4] <= 'd0;
    kernel_img_mul_2[5] <= 'd0;
    kernel_img_mul_2[6] <= 'd0;
    kernel_img_mul_2[7] <= 'd0;
    kernel_img_mul_2[8] <= 'd0;
    kernel_img_mul_2[9] <= 'd0;
    kernel_img_mul_2[10] <= 'd0;
    kernel_img_mul_2[11] <= 'd0;
    kernel_img_mul_2[12] <= 'd0;
    kernel_img_mul_2[13] <= 'd0;
    kernel_img_mul_2[14] <= 'd0;
    kernel_img_mul_2[15] <= 'd0;
    kernel_img_mul_2[16] <= 'd0;
    kernel_img_mul_2[17] <= 'd0;
    kernel_img_mul_2[18] <= 'd0;
    kernel_img_mul_2[19] <= 'd0;
    kernel_img_mul_2[20] <= 'd0;
    kernel_img_mul_2[21] <= 'd0;
    kernel_img_mul_2[22] <= 'd0;
    kernel_img_mul_2[23] <= 'd0;
    kernel_img_mul_2[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_2[0] <= { {8{1'b0}},layer0[2][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_2[1] <= { {8{1'b0}},layer0[2][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_2[2] <= { {8{1'b0}},layer0[2][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_2[3] <= { {8{1'b0}},layer0[2][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_2[4] <= { {8{1'b0}},layer0[2][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_2[5] <= { {8{1'b0}},layer1[2][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_2[6] <= { {8{1'b0}},layer1[2][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_2[7] <= { {8{1'b0}},layer1[2][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_2[8] <= { {8{1'b0}},layer1[2][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_2[9] <= { {8{1'b0}},layer1[2][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_2[10] <= { {8{1'b0}},layer2[2][7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_2[11] <= { {8{1'b0}},layer2[2][15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_2[12] <= { {8{1'b0}},layer2[2][23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_2[13] <= { {8{1'b0}},layer2[2][31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_2[14] <= { {8{1'b0}},layer2[2][39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_2[15] <= { {8{1'b0}},layer3[2][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_2[16] <= { {8{1'b0}},layer3[2][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_2[17] <= { {8{1'b0}},layer3[2][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_2[18] <= { {8{1'b0}},layer3[2][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_2[19] <= { {8{1'b0}},layer3[2][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_2[20] <= { {8{1'b0}},layer4[2][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_2[21] <= { {8{1'b0}},layer4[2][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_2[22] <= { {8{1'b0}},layer4[2][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_2[23] <= { {8{1'b0}},layer4[2][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_2[24] <= { {8{1'b0}},layer4[2][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_2;
reg  [15:0]  kernel_img_sum_2_2;
reg  [15:0]  kernel_img_sum_3_2;
reg  [15:0]  kernel_img_sum_4_2;
reg  [15:0]  kernel_img_sum_5_2;
reg  [15:0]  kernel_img_sum_6_2;
reg  [15:0]  kernel_img_sum_7_2;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_2 <= kernel_img_mul_2[0] + kernel_img_mul_2[1] + kernel_img_mul_2[2] + kernel_img_mul_2[3] + kernel_img_mul_2[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_2 <= kernel_img_mul_2[5] + kernel_img_mul_2[6] + kernel_img_mul_2[7] + kernel_img_mul_2[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_2 <= kernel_img_mul_2[9] + kernel_img_mul_2[10] + kernel_img_mul_2[11] + kernel_img_mul_2[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_2 <= kernel_img_mul_2[13] + kernel_img_mul_2[14] + kernel_img_mul_2[15] + kernel_img_mul_2[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_2 <= kernel_img_mul_2[17] + kernel_img_mul_2[18] + kernel_img_mul_2[19] + kernel_img_mul_2[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_2 <= kernel_img_mul_2[21] + kernel_img_mul_2[22] + kernel_img_mul_2[23] + kernel_img_mul_2[24];
  end
end
always@(*) begin
  kernel_img_sum_7_2 = kernel_img_sum_1_2 + kernel_img_sum_2_2 + kernel_img_sum_3_2 + kernel_img_sum_4_2 + kernel_img_sum_5_2 + kernel_img_sum_6_2;
end
reg  [15:0]  kernel_img_mul_3[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_3[0] <= 'd0;
    kernel_img_mul_3[1] <= 'd0;
    kernel_img_mul_3[2] <= 'd0;
    kernel_img_mul_3[3] <= 'd0;
    kernel_img_mul_3[4] <= 'd0;
    kernel_img_mul_3[5] <= 'd0;
    kernel_img_mul_3[6] <= 'd0;
    kernel_img_mul_3[7] <= 'd0;
    kernel_img_mul_3[8] <= 'd0;
    kernel_img_mul_3[9] <= 'd0;
    kernel_img_mul_3[10] <= 'd0;
    kernel_img_mul_3[11] <= 'd0;
    kernel_img_mul_3[12] <= 'd0;
    kernel_img_mul_3[13] <= 'd0;
    kernel_img_mul_3[14] <= 'd0;
    kernel_img_mul_3[15] <= 'd0;
    kernel_img_mul_3[16] <= 'd0;
    kernel_img_mul_3[17] <= 'd0;
    kernel_img_mul_3[18] <= 'd0;
    kernel_img_mul_3[19] <= 'd0;
    kernel_img_mul_3[20] <= 'd0;
    kernel_img_mul_3[21] <= 'd0;
    kernel_img_mul_3[22] <= 'd0;
    kernel_img_mul_3[23] <= 'd0;
    kernel_img_mul_3[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_3[0] <= { {8{1'b0}},layer0[3][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_3[1] <= { {8{1'b0}},layer0[3][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_3[2] <= { {8{1'b0}},layer0[3][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_3[3] <= { {8{1'b0}},layer0[3][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_3[4] <= { {8{1'b0}},layer0[3][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_3[5] <= { {8{1'b0}},layer1[3][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_3[6] <= { {8{1'b0}},layer1[3][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_3[7] <= { {8{1'b0}},layer1[3][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_3[8] <= { {8{1'b0}},layer1[3][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_3[9] <= { {8{1'b0}},layer1[3][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_3[10] <= { {8{1'b0}},layer2[3][7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_3[11] <= { {8{1'b0}},layer2[3][15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_3[12] <= { {8{1'b0}},layer2[3][23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_3[13] <= { {8{1'b0}},layer2[3][31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_3[14] <= { {8{1'b0}},layer2[3][39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_3[15] <= { {8{1'b0}},layer3[3][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_3[16] <= { {8{1'b0}},layer3[3][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_3[17] <= { {8{1'b0}},layer3[3][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_3[18] <= { {8{1'b0}},layer3[3][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_3[19] <= { {8{1'b0}},layer3[3][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_3[20] <= { {8{1'b0}},layer4[3][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_3[21] <= { {8{1'b0}},layer4[3][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_3[22] <= { {8{1'b0}},layer4[3][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_3[23] <= { {8{1'b0}},layer4[3][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_3[24] <= { {8{1'b0}},layer4[3][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_3;
reg  [15:0]  kernel_img_sum_2_3;
reg  [15:0]  kernel_img_sum_3_3;
reg  [15:0]  kernel_img_sum_4_3;
reg  [15:0]  kernel_img_sum_5_3;
reg  [15:0]  kernel_img_sum_6_3;
reg  [15:0]  kernel_img_sum_7_3;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_3 <= kernel_img_mul_3[0] + kernel_img_mul_3[1] + kernel_img_mul_3[2] + kernel_img_mul_3[3] + kernel_img_mul_3[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_3 <= kernel_img_mul_3[5] + kernel_img_mul_3[6] + kernel_img_mul_3[7] + kernel_img_mul_3[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_3 <= kernel_img_mul_3[9] + kernel_img_mul_3[10] + kernel_img_mul_3[11] + kernel_img_mul_3[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_3 <= kernel_img_mul_3[13] + kernel_img_mul_3[14] + kernel_img_mul_3[15] + kernel_img_mul_3[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_3 <= kernel_img_mul_3[17] + kernel_img_mul_3[18] + kernel_img_mul_3[19] + kernel_img_mul_3[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_3 <= kernel_img_mul_3[21] + kernel_img_mul_3[22] + kernel_img_mul_3[23] + kernel_img_mul_3[24];
  end
end
always@(*) begin
  kernel_img_sum_7_3 = kernel_img_sum_1_3 + kernel_img_sum_2_3 + kernel_img_sum_3_3 + kernel_img_sum_4_3 + kernel_img_sum_5_3 + kernel_img_sum_6_3;
end
reg  [15:0]  kernel_img_mul_4[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_4[0] <= 'd0;
    kernel_img_mul_4[1] <= 'd0;
    kernel_img_mul_4[2] <= 'd0;
    kernel_img_mul_4[3] <= 'd0;
    kernel_img_mul_4[4] <= 'd0;
    kernel_img_mul_4[5] <= 'd0;
    kernel_img_mul_4[6] <= 'd0;
    kernel_img_mul_4[7] <= 'd0;
    kernel_img_mul_4[8] <= 'd0;
    kernel_img_mul_4[9] <= 'd0;
    kernel_img_mul_4[10] <= 'd0;
    kernel_img_mul_4[11] <= 'd0;
    kernel_img_mul_4[12] <= 'd0;
    kernel_img_mul_4[13] <= 'd0;
    kernel_img_mul_4[14] <= 'd0;
    kernel_img_mul_4[15] <= 'd0;
    kernel_img_mul_4[16] <= 'd0;
    kernel_img_mul_4[17] <= 'd0;
    kernel_img_mul_4[18] <= 'd0;
    kernel_img_mul_4[19] <= 'd0;
    kernel_img_mul_4[20] <= 'd0;
    kernel_img_mul_4[21] <= 'd0;
    kernel_img_mul_4[22] <= 'd0;
    kernel_img_mul_4[23] <= 'd0;
    kernel_img_mul_4[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_4[0] <= { {8{1'b0}},layer0[4][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_4[1] <= { {8{1'b0}},layer0[4][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_4[2] <= { {8{1'b0}},layer0[4][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_4[3] <= { {8{1'b0}},layer0[4][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_4[4] <= { {8{1'b0}},layer0[4][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_4[5] <= { {8{1'b0}},layer1[4][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_4[6] <= { {8{1'b0}},layer1[4][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_4[7] <= { {8{1'b0}},layer1[4][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_4[8] <= { {8{1'b0}},layer1[4][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_4[9] <= { {8{1'b0}},layer1[4][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_4[10] <= { {8{1'b0}},layer2[4][7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_4[11] <= { {8{1'b0}},layer2[4][15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_4[12] <= { {8{1'b0}},layer2[4][23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_4[13] <= { {8{1'b0}},layer2[4][31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_4[14] <= { {8{1'b0}},layer2[4][39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_4[15] <= { {8{1'b0}},layer3[4][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_4[16] <= { {8{1'b0}},layer3[4][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_4[17] <= { {8{1'b0}},layer3[4][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_4[18] <= { {8{1'b0}},layer3[4][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_4[19] <= { {8{1'b0}},layer3[4][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_4[20] <= { {8{1'b0}},layer4[4][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_4[21] <= { {8{1'b0}},layer4[4][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_4[22] <= { {8{1'b0}},layer4[4][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_4[23] <= { {8{1'b0}},layer4[4][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_4[24] <= { {8{1'b0}},layer4[4][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_4;
reg  [15:0]  kernel_img_sum_2_4;
reg  [15:0]  kernel_img_sum_3_4;
reg  [15:0]  kernel_img_sum_4_4;
reg  [15:0]  kernel_img_sum_5_4;
reg  [15:0]  kernel_img_sum_6_4;
reg  [15:0]  kernel_img_sum_7_4;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_4 <= kernel_img_mul_4[0] + kernel_img_mul_4[1] + kernel_img_mul_4[2] + kernel_img_mul_4[3] + kernel_img_mul_4[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_4 <= kernel_img_mul_4[5] + kernel_img_mul_4[6] + kernel_img_mul_4[7] + kernel_img_mul_4[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_4 <= kernel_img_mul_4[9] + kernel_img_mul_4[10] + kernel_img_mul_4[11] + kernel_img_mul_4[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_4 <= kernel_img_mul_4[13] + kernel_img_mul_4[14] + kernel_img_mul_4[15] + kernel_img_mul_4[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_4 <= kernel_img_mul_4[17] + kernel_img_mul_4[18] + kernel_img_mul_4[19] + kernel_img_mul_4[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_4 <= kernel_img_mul_4[21] + kernel_img_mul_4[22] + kernel_img_mul_4[23] + kernel_img_mul_4[24];
  end
end
always@(*) begin
  kernel_img_sum_7_4 = kernel_img_sum_1_4 + kernel_img_sum_2_4 + kernel_img_sum_3_4 + kernel_img_sum_4_4 + kernel_img_sum_5_4 + kernel_img_sum_6_4;
end
reg  [15:0]  kernel_img_mul_5[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_5[0] <= 'd0;
    kernel_img_mul_5[1] <= 'd0;
    kernel_img_mul_5[2] <= 'd0;
    kernel_img_mul_5[3] <= 'd0;
    kernel_img_mul_5[4] <= 'd0;
    kernel_img_mul_5[5] <= 'd0;
    kernel_img_mul_5[6] <= 'd0;
    kernel_img_mul_5[7] <= 'd0;
    kernel_img_mul_5[8] <= 'd0;
    kernel_img_mul_5[9] <= 'd0;
    kernel_img_mul_5[10] <= 'd0;
    kernel_img_mul_5[11] <= 'd0;
    kernel_img_mul_5[12] <= 'd0;
    kernel_img_mul_5[13] <= 'd0;
    kernel_img_mul_5[14] <= 'd0;
    kernel_img_mul_5[15] <= 'd0;
    kernel_img_mul_5[16] <= 'd0;
    kernel_img_mul_5[17] <= 'd0;
    kernel_img_mul_5[18] <= 'd0;
    kernel_img_mul_5[19] <= 'd0;
    kernel_img_mul_5[20] <= 'd0;
    kernel_img_mul_5[21] <= 'd0;
    kernel_img_mul_5[22] <= 'd0;
    kernel_img_mul_5[23] <= 'd0;
    kernel_img_mul_5[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_5[0] <= { {8{1'b0}},layer0[5][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_5[1] <= { {8{1'b0}},layer0[5][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_5[2] <= { {8{1'b0}},layer0[5][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_5[3] <= { {8{1'b0}},layer0[5][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_5[4] <= { {8{1'b0}},layer0[5][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_5[5] <= { {8{1'b0}},layer1[5][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_5[6] <= { {8{1'b0}},layer1[5][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_5[7] <= { {8{1'b0}},layer1[5][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_5[8] <= { {8{1'b0}},layer1[5][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_5[9] <= { {8{1'b0}},layer1[5][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_5[10] <= { {8{1'b0}},layer2[5][7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_5[11] <= { {8{1'b0}},layer2[5][15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_5[12] <= { {8{1'b0}},layer2[5][23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_5[13] <= { {8{1'b0}},layer2[5][31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_5[14] <= { {8{1'b0}},layer2[5][39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_5[15] <= { {8{1'b0}},layer3[5][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_5[16] <= { {8{1'b0}},layer3[5][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_5[17] <= { {8{1'b0}},layer3[5][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_5[18] <= { {8{1'b0}},layer3[5][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_5[19] <= { {8{1'b0}},layer3[5][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_5[20] <= { {8{1'b0}},layer4[5][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_5[21] <= { {8{1'b0}},layer4[5][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_5[22] <= { {8{1'b0}},layer4[5][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_5[23] <= { {8{1'b0}},layer4[5][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_5[24] <= { {8{1'b0}},layer4[5][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_5;
reg  [15:0]  kernel_img_sum_2_5;
reg  [15:0]  kernel_img_sum_3_5;
reg  [15:0]  kernel_img_sum_4_5;
reg  [15:0]  kernel_img_sum_5_5;
reg  [15:0]  kernel_img_sum_6_5;
reg  [15:0]  kernel_img_sum_7_5;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_5 <= kernel_img_mul_5[0] + kernel_img_mul_5[1] + kernel_img_mul_5[2] + kernel_img_mul_5[3] + kernel_img_mul_5[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_5 <= kernel_img_mul_5[5] + kernel_img_mul_5[6] + kernel_img_mul_5[7] + kernel_img_mul_5[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_5 <= kernel_img_mul_5[9] + kernel_img_mul_5[10] + kernel_img_mul_5[11] + kernel_img_mul_5[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_5 <= kernel_img_mul_5[13] + kernel_img_mul_5[14] + kernel_img_mul_5[15] + kernel_img_mul_5[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_5 <= kernel_img_mul_5[17] + kernel_img_mul_5[18] + kernel_img_mul_5[19] + kernel_img_mul_5[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_5 <= kernel_img_mul_5[21] + kernel_img_mul_5[22] + kernel_img_mul_5[23] + kernel_img_mul_5[24];
  end
end
always@(*) begin
  kernel_img_sum_7_5 = kernel_img_sum_1_5 + kernel_img_sum_2_5 + kernel_img_sum_3_5 + kernel_img_sum_4_5 + kernel_img_sum_5_5 + kernel_img_sum_6_5;
end
reg  [15:0]  kernel_img_mul_6[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_6[0] <= 'd0;
    kernel_img_mul_6[1] <= 'd0;
    kernel_img_mul_6[2] <= 'd0;
    kernel_img_mul_6[3] <= 'd0;
    kernel_img_mul_6[4] <= 'd0;
    kernel_img_mul_6[5] <= 'd0;
    kernel_img_mul_6[6] <= 'd0;
    kernel_img_mul_6[7] <= 'd0;
    kernel_img_mul_6[8] <= 'd0;
    kernel_img_mul_6[9] <= 'd0;
    kernel_img_mul_6[10] <= 'd0;
    kernel_img_mul_6[11] <= 'd0;
    kernel_img_mul_6[12] <= 'd0;
    kernel_img_mul_6[13] <= 'd0;
    kernel_img_mul_6[14] <= 'd0;
    kernel_img_mul_6[15] <= 'd0;
    kernel_img_mul_6[16] <= 'd0;
    kernel_img_mul_6[17] <= 'd0;
    kernel_img_mul_6[18] <= 'd0;
    kernel_img_mul_6[19] <= 'd0;
    kernel_img_mul_6[20] <= 'd0;
    kernel_img_mul_6[21] <= 'd0;
    kernel_img_mul_6[22] <= 'd0;
    kernel_img_mul_6[23] <= 'd0;
    kernel_img_mul_6[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_6[0] <= { {8{1'b0}},layer0[6][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_6[1] <= { {8{1'b0}},layer0[6][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_6[2] <= { {8{1'b0}},layer0[6][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_6[3] <= { {8{1'b0}},layer0[6][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_6[4] <= { {8{1'b0}},layer0[6][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_6[5] <= { {8{1'b0}},layer1[6][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_6[6] <= { {8{1'b0}},layer1[6][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_6[7] <= { {8{1'b0}},layer1[6][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_6[8] <= { {8{1'b0}},layer1[6][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_6[9] <= { {8{1'b0}},layer1[6][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_6[10] <= { {8{1'b0}},layer2[6][7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_6[11] <= { {8{1'b0}},layer2[6][15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_6[12] <= { {8{1'b0}},layer2[6][23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_6[13] <= { {8{1'b0}},layer2[6][31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_6[14] <= { {8{1'b0}},layer2[6][39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_6[15] <= { {8{1'b0}},layer3[6][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_6[16] <= { {8{1'b0}},layer3[6][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_6[17] <= { {8{1'b0}},layer3[6][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_6[18] <= { {8{1'b0}},layer3[6][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_6[19] <= { {8{1'b0}},layer3[6][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_6[20] <= { {8{1'b0}},layer4[6][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_6[21] <= { {8{1'b0}},layer4[6][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_6[22] <= { {8{1'b0}},layer4[6][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_6[23] <= { {8{1'b0}},layer4[6][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_6[24] <= { {8{1'b0}},layer4[6][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_6;
reg  [15:0]  kernel_img_sum_2_6;
reg  [15:0]  kernel_img_sum_3_6;
reg  [15:0]  kernel_img_sum_4_6;
reg  [15:0]  kernel_img_sum_5_6;
reg  [15:0]  kernel_img_sum_6_6;
reg  [15:0]  kernel_img_sum_7_6;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_6 <= kernel_img_mul_6[0] + kernel_img_mul_6[1] + kernel_img_mul_6[2] + kernel_img_mul_6[3] + kernel_img_mul_6[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_6 <= kernel_img_mul_6[5] + kernel_img_mul_6[6] + kernel_img_mul_6[7] + kernel_img_mul_6[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_6 <= kernel_img_mul_6[9] + kernel_img_mul_6[10] + kernel_img_mul_6[11] + kernel_img_mul_6[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_6 <= kernel_img_mul_6[13] + kernel_img_mul_6[14] + kernel_img_mul_6[15] + kernel_img_mul_6[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_6 <= kernel_img_mul_6[17] + kernel_img_mul_6[18] + kernel_img_mul_6[19] + kernel_img_mul_6[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_6 <= kernel_img_mul_6[21] + kernel_img_mul_6[22] + kernel_img_mul_6[23] + kernel_img_mul_6[24];
  end
end
always@(*) begin
  kernel_img_sum_7_6 = kernel_img_sum_1_6 + kernel_img_sum_2_6 + kernel_img_sum_3_6 + kernel_img_sum_4_6 + kernel_img_sum_5_6 + kernel_img_sum_6_6;
end
reg  [15:0]  kernel_img_mul_7[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_7[0] <= 'd0;
    kernel_img_mul_7[1] <= 'd0;
    kernel_img_mul_7[2] <= 'd0;
    kernel_img_mul_7[3] <= 'd0;
    kernel_img_mul_7[4] <= 'd0;
    kernel_img_mul_7[5] <= 'd0;
    kernel_img_mul_7[6] <= 'd0;
    kernel_img_mul_7[7] <= 'd0;
    kernel_img_mul_7[8] <= 'd0;
    kernel_img_mul_7[9] <= 'd0;
    kernel_img_mul_7[10] <= 'd0;
    kernel_img_mul_7[11] <= 'd0;
    kernel_img_mul_7[12] <= 'd0;
    kernel_img_mul_7[13] <= 'd0;
    kernel_img_mul_7[14] <= 'd0;
    kernel_img_mul_7[15] <= 'd0;
    kernel_img_mul_7[16] <= 'd0;
    kernel_img_mul_7[17] <= 'd0;
    kernel_img_mul_7[18] <= 'd0;
    kernel_img_mul_7[19] <= 'd0;
    kernel_img_mul_7[20] <= 'd0;
    kernel_img_mul_7[21] <= 'd0;
    kernel_img_mul_7[22] <= 'd0;
    kernel_img_mul_7[23] <= 'd0;
    kernel_img_mul_7[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_7[0] <= { {8{1'b0}},layer0[7][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_7[1] <= { {8{1'b0}},layer0[7][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_7[2] <= { {8{1'b0}},layer0[7][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_7[3] <= { {8{1'b0}},layer0[7][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_7[4] <= { {8{1'b0}},layer0[7][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_7[5] <= { {8{1'b0}},layer1[7][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_7[6] <= { {8{1'b0}},layer1[7][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_7[7] <= { {8{1'b0}},layer1[7][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_7[8] <= { {8{1'b0}},layer1[7][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_7[9] <= { {8{1'b0}},layer1[7][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_7[10] <= { {8{1'b0}},layer2[7][7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_7[11] <= { {8{1'b0}},layer2[7][15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_7[12] <= { {8{1'b0}},layer2[7][23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_7[13] <= { {8{1'b0}},layer2[7][31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_7[14] <= { {8{1'b0}},layer2[7][39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_7[15] <= { {8{1'b0}},layer3[7][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_7[16] <= { {8{1'b0}},layer3[7][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_7[17] <= { {8{1'b0}},layer3[7][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_7[18] <= { {8{1'b0}},layer3[7][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_7[19] <= { {8{1'b0}},layer3[7][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_7[20] <= { {8{1'b0}},layer4[7][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_7[21] <= { {8{1'b0}},layer4[7][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_7[22] <= { {8{1'b0}},layer4[7][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_7[23] <= { {8{1'b0}},layer4[7][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_7[24] <= { {8{1'b0}},layer4[7][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_7;
reg  [15:0]  kernel_img_sum_2_7;
reg  [15:0]  kernel_img_sum_3_7;
reg  [15:0]  kernel_img_sum_4_7;
reg  [15:0]  kernel_img_sum_5_7;
reg  [15:0]  kernel_img_sum_6_7;
reg  [15:0]  kernel_img_sum_7_7;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_7 <= kernel_img_mul_7[0] + kernel_img_mul_7[1] + kernel_img_mul_7[2] + kernel_img_mul_7[3] + kernel_img_mul_7[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_7 <= kernel_img_mul_7[5] + kernel_img_mul_7[6] + kernel_img_mul_7[7] + kernel_img_mul_7[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_7 <= kernel_img_mul_7[9] + kernel_img_mul_7[10] + kernel_img_mul_7[11] + kernel_img_mul_7[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_7 <= kernel_img_mul_7[13] + kernel_img_mul_7[14] + kernel_img_mul_7[15] + kernel_img_mul_7[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_7 <= kernel_img_mul_7[17] + kernel_img_mul_7[18] + kernel_img_mul_7[19] + kernel_img_mul_7[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_7 <= kernel_img_mul_7[21] + kernel_img_mul_7[22] + kernel_img_mul_7[23] + kernel_img_mul_7[24];
  end
end
always@(*) begin
  kernel_img_sum_7_7 = kernel_img_sum_1_7 + kernel_img_sum_2_7 + kernel_img_sum_3_7 + kernel_img_sum_4_7 + kernel_img_sum_5_7 + kernel_img_sum_6_7;
end
reg  [15:0]  kernel_img_mul_8[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_8[0] <= 'd0;
    kernel_img_mul_8[1] <= 'd0;
    kernel_img_mul_8[2] <= 'd0;
    kernel_img_mul_8[3] <= 'd0;
    kernel_img_mul_8[4] <= 'd0;
    kernel_img_mul_8[5] <= 'd0;
    kernel_img_mul_8[6] <= 'd0;
    kernel_img_mul_8[7] <= 'd0;
    kernel_img_mul_8[8] <= 'd0;
    kernel_img_mul_8[9] <= 'd0;
    kernel_img_mul_8[10] <= 'd0;
    kernel_img_mul_8[11] <= 'd0;
    kernel_img_mul_8[12] <= 'd0;
    kernel_img_mul_8[13] <= 'd0;
    kernel_img_mul_8[14] <= 'd0;
    kernel_img_mul_8[15] <= 'd0;
    kernel_img_mul_8[16] <= 'd0;
    kernel_img_mul_8[17] <= 'd0;
    kernel_img_mul_8[18] <= 'd0;
    kernel_img_mul_8[19] <= 'd0;
    kernel_img_mul_8[20] <= 'd0;
    kernel_img_mul_8[21] <= 'd0;
    kernel_img_mul_8[22] <= 'd0;
    kernel_img_mul_8[23] <= 'd0;
    kernel_img_mul_8[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_8[0] <= { {8{1'b0}},layer0[8][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_8[1] <= { {8{1'b0}},layer0[8][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_8[2] <= { {8{1'b0}},layer0[8][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_8[3] <= { {8{1'b0}},layer0[8][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_8[4] <= { {8{1'b0}},layer0[8][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_8[5] <= { {8{1'b0}},layer1[8][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_8[6] <= { {8{1'b0}},layer1[8][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_8[7] <= { {8{1'b0}},layer1[8][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_8[8] <= { {8{1'b0}},layer1[8][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_8[9] <= { {8{1'b0}},layer1[8][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_8[10] <= { {8{1'b0}},layer2[8][7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_8[11] <= { {8{1'b0}},layer2[8][15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_8[12] <= { {8{1'b0}},layer2[8][23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_8[13] <= { {8{1'b0}},layer2[8][31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_8[14] <= { {8{1'b0}},layer2[8][39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_8[15] <= { {8{1'b0}},layer3[8][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_8[16] <= { {8{1'b0}},layer3[8][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_8[17] <= { {8{1'b0}},layer3[8][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_8[18] <= { {8{1'b0}},layer3[8][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_8[19] <= { {8{1'b0}},layer3[8][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_8[20] <= { {8{1'b0}},layer4[8][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_8[21] <= { {8{1'b0}},layer4[8][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_8[22] <= { {8{1'b0}},layer4[8][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_8[23] <= { {8{1'b0}},layer4[8][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_8[24] <= { {8{1'b0}},layer4[8][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_8;
reg  [15:0]  kernel_img_sum_2_8;
reg  [15:0]  kernel_img_sum_3_8;
reg  [15:0]  kernel_img_sum_4_8;
reg  [15:0]  kernel_img_sum_5_8;
reg  [15:0]  kernel_img_sum_6_8;
reg  [15:0]  kernel_img_sum_7_8;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_8 <= kernel_img_mul_8[0] + kernel_img_mul_8[1] + kernel_img_mul_8[2] + kernel_img_mul_8[3] + kernel_img_mul_8[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_8 <= kernel_img_mul_8[5] + kernel_img_mul_8[6] + kernel_img_mul_8[7] + kernel_img_mul_8[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_8 <= kernel_img_mul_8[9] + kernel_img_mul_8[10] + kernel_img_mul_8[11] + kernel_img_mul_8[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_8 <= kernel_img_mul_8[13] + kernel_img_mul_8[14] + kernel_img_mul_8[15] + kernel_img_mul_8[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_8 <= kernel_img_mul_8[17] + kernel_img_mul_8[18] + kernel_img_mul_8[19] + kernel_img_mul_8[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_8 <= kernel_img_mul_8[21] + kernel_img_mul_8[22] + kernel_img_mul_8[23] + kernel_img_mul_8[24];
  end
end
always@(*) begin
  kernel_img_sum_7_8 = kernel_img_sum_1_8 + kernel_img_sum_2_8 + kernel_img_sum_3_8 + kernel_img_sum_4_8 + kernel_img_sum_5_8 + kernel_img_sum_6_8;
end
reg  [15:0]  kernel_img_mul_9[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_9[0] <= 'd0;
    kernel_img_mul_9[1] <= 'd0;
    kernel_img_mul_9[2] <= 'd0;
    kernel_img_mul_9[3] <= 'd0;
    kernel_img_mul_9[4] <= 'd0;
    kernel_img_mul_9[5] <= 'd0;
    kernel_img_mul_9[6] <= 'd0;
    kernel_img_mul_9[7] <= 'd0;
    kernel_img_mul_9[8] <= 'd0;
    kernel_img_mul_9[9] <= 'd0;
    kernel_img_mul_9[10] <= 'd0;
    kernel_img_mul_9[11] <= 'd0;
    kernel_img_mul_9[12] <= 'd0;
    kernel_img_mul_9[13] <= 'd0;
    kernel_img_mul_9[14] <= 'd0;
    kernel_img_mul_9[15] <= 'd0;
    kernel_img_mul_9[16] <= 'd0;
    kernel_img_mul_9[17] <= 'd0;
    kernel_img_mul_9[18] <= 'd0;
    kernel_img_mul_9[19] <= 'd0;
    kernel_img_mul_9[20] <= 'd0;
    kernel_img_mul_9[21] <= 'd0;
    kernel_img_mul_9[22] <= 'd0;
    kernel_img_mul_9[23] <= 'd0;
    kernel_img_mul_9[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_9[0] <= { {8{1'b0}},layer0[9][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_9[1] <= { {8{1'b0}},layer0[9][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_9[2] <= { {8{1'b0}},layer0[9][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_9[3] <= { {8{1'b0}},layer0[9][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_9[4] <= { {8{1'b0}},layer0[9][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_9[5] <= { {8{1'b0}},layer1[9][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_9[6] <= { {8{1'b0}},layer1[9][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_9[7] <= { {8{1'b0}},layer1[9][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_9[8] <= { {8{1'b0}},layer1[9][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_9[9] <= { {8{1'b0}},layer1[9][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_9[10] <= { {8{1'b0}},layer2[9][7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_9[11] <= { {8{1'b0}},layer2[9][15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_9[12] <= { {8{1'b0}},layer2[9][23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_9[13] <= { {8{1'b0}},layer2[9][31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_9[14] <= { {8{1'b0}},layer2[9][39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_9[15] <= { {8{1'b0}},layer3[9][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_9[16] <= { {8{1'b0}},layer3[9][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_9[17] <= { {8{1'b0}},layer3[9][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_9[18] <= { {8{1'b0}},layer3[9][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_9[19] <= { {8{1'b0}},layer3[9][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_9[20] <= { {8{1'b0}},layer4[9][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_9[21] <= { {8{1'b0}},layer4[9][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_9[22] <= { {8{1'b0}},layer4[9][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_9[23] <= { {8{1'b0}},layer4[9][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_9[24] <= { {8{1'b0}},layer4[9][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_9;
reg  [15:0]  kernel_img_sum_2_9;
reg  [15:0]  kernel_img_sum_3_9;
reg  [15:0]  kernel_img_sum_4_9;
reg  [15:0]  kernel_img_sum_5_9;
reg  [15:0]  kernel_img_sum_6_9;
reg  [15:0]  kernel_img_sum_7_9;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_9 <= kernel_img_mul_9[0] + kernel_img_mul_9[1] + kernel_img_mul_9[2] + kernel_img_mul_9[3] + kernel_img_mul_9[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_9 <= kernel_img_mul_9[5] + kernel_img_mul_9[6] + kernel_img_mul_9[7] + kernel_img_mul_9[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_9 <= kernel_img_mul_9[9] + kernel_img_mul_9[10] + kernel_img_mul_9[11] + kernel_img_mul_9[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_9 <= kernel_img_mul_9[13] + kernel_img_mul_9[14] + kernel_img_mul_9[15] + kernel_img_mul_9[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_9 <= kernel_img_mul_9[17] + kernel_img_mul_9[18] + kernel_img_mul_9[19] + kernel_img_mul_9[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_9 <= kernel_img_mul_9[21] + kernel_img_mul_9[22] + kernel_img_mul_9[23] + kernel_img_mul_9[24];
  end
end
always@(*) begin
  kernel_img_sum_7_9 = kernel_img_sum_1_9 + kernel_img_sum_2_9 + kernel_img_sum_3_9 + kernel_img_sum_4_9 + kernel_img_sum_5_9 + kernel_img_sum_6_9;
end
reg  [15:0]  kernel_img_mul_10[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_10[0] <= 'd0;
    kernel_img_mul_10[1] <= 'd0;
    kernel_img_mul_10[2] <= 'd0;
    kernel_img_mul_10[3] <= 'd0;
    kernel_img_mul_10[4] <= 'd0;
    kernel_img_mul_10[5] <= 'd0;
    kernel_img_mul_10[6] <= 'd0;
    kernel_img_mul_10[7] <= 'd0;
    kernel_img_mul_10[8] <= 'd0;
    kernel_img_mul_10[9] <= 'd0;
    kernel_img_mul_10[10] <= 'd0;
    kernel_img_mul_10[11] <= 'd0;
    kernel_img_mul_10[12] <= 'd0;
    kernel_img_mul_10[13] <= 'd0;
    kernel_img_mul_10[14] <= 'd0;
    kernel_img_mul_10[15] <= 'd0;
    kernel_img_mul_10[16] <= 'd0;
    kernel_img_mul_10[17] <= 'd0;
    kernel_img_mul_10[18] <= 'd0;
    kernel_img_mul_10[19] <= 'd0;
    kernel_img_mul_10[20] <= 'd0;
    kernel_img_mul_10[21] <= 'd0;
    kernel_img_mul_10[22] <= 'd0;
    kernel_img_mul_10[23] <= 'd0;
    kernel_img_mul_10[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_10[0] <= { {8{1'b0}},layer0[10][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_10[1] <= { {8{1'b0}},layer0[10][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_10[2] <= { {8{1'b0}},layer0[10][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_10[3] <= { {8{1'b0}},layer0[10][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_10[4] <= { {8{1'b0}},layer0[10][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_10[5] <= { {8{1'b0}},layer1[10][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_10[6] <= { {8{1'b0}},layer1[10][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_10[7] <= { {8{1'b0}},layer1[10][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_10[8] <= { {8{1'b0}},layer1[10][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_10[9] <= { {8{1'b0}},layer1[10][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_10[10] <= { {8{1'b0}},layer2[10][7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_10[11] <= { {8{1'b0}},layer2[10][15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_10[12] <= { {8{1'b0}},layer2[10][23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_10[13] <= { {8{1'b0}},layer2[10][31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_10[14] <= { {8{1'b0}},layer2[10][39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_10[15] <= { {8{1'b0}},layer3[10][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_10[16] <= { {8{1'b0}},layer3[10][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_10[17] <= { {8{1'b0}},layer3[10][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_10[18] <= { {8{1'b0}},layer3[10][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_10[19] <= { {8{1'b0}},layer3[10][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_10[20] <= { {8{1'b0}},layer4[10][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_10[21] <= { {8{1'b0}},layer4[10][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_10[22] <= { {8{1'b0}},layer4[10][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_10[23] <= { {8{1'b0}},layer4[10][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_10[24] <= { {8{1'b0}},layer4[10][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_10;
reg  [15:0]  kernel_img_sum_2_10;
reg  [15:0]  kernel_img_sum_3_10;
reg  [15:0]  kernel_img_sum_4_10;
reg  [15:0]  kernel_img_sum_5_10;
reg  [15:0]  kernel_img_sum_6_10;
reg  [15:0]  kernel_img_sum_7_10;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_10 <= kernel_img_mul_10[0] + kernel_img_mul_10[1] + kernel_img_mul_10[2] + kernel_img_mul_10[3] + kernel_img_mul_10[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_10 <= kernel_img_mul_10[5] + kernel_img_mul_10[6] + kernel_img_mul_10[7] + kernel_img_mul_10[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_10 <= kernel_img_mul_10[9] + kernel_img_mul_10[10] + kernel_img_mul_10[11] + kernel_img_mul_10[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_10 <= kernel_img_mul_10[13] + kernel_img_mul_10[14] + kernel_img_mul_10[15] + kernel_img_mul_10[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_10 <= kernel_img_mul_10[17] + kernel_img_mul_10[18] + kernel_img_mul_10[19] + kernel_img_mul_10[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_10 <= kernel_img_mul_10[21] + kernel_img_mul_10[22] + kernel_img_mul_10[23] + kernel_img_mul_10[24];
  end
end
always@(*) begin
  kernel_img_sum_7_10 = kernel_img_sum_1_10 + kernel_img_sum_2_10 + kernel_img_sum_3_10 + kernel_img_sum_4_10 + kernel_img_sum_5_10 + kernel_img_sum_6_10;
end
reg  [15:0]  kernel_img_mul_11[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_11[0] <= 'd0;
    kernel_img_mul_11[1] <= 'd0;
    kernel_img_mul_11[2] <= 'd0;
    kernel_img_mul_11[3] <= 'd0;
    kernel_img_mul_11[4] <= 'd0;
    kernel_img_mul_11[5] <= 'd0;
    kernel_img_mul_11[6] <= 'd0;
    kernel_img_mul_11[7] <= 'd0;
    kernel_img_mul_11[8] <= 'd0;
    kernel_img_mul_11[9] <= 'd0;
    kernel_img_mul_11[10] <= 'd0;
    kernel_img_mul_11[11] <= 'd0;
    kernel_img_mul_11[12] <= 'd0;
    kernel_img_mul_11[13] <= 'd0;
    kernel_img_mul_11[14] <= 'd0;
    kernel_img_mul_11[15] <= 'd0;
    kernel_img_mul_11[16] <= 'd0;
    kernel_img_mul_11[17] <= 'd0;
    kernel_img_mul_11[18] <= 'd0;
    kernel_img_mul_11[19] <= 'd0;
    kernel_img_mul_11[20] <= 'd0;
    kernel_img_mul_11[21] <= 'd0;
    kernel_img_mul_11[22] <= 'd0;
    kernel_img_mul_11[23] <= 'd0;
    kernel_img_mul_11[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_11[0] <= { {8{1'b0}},layer0[11][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_11[1] <= { {8{1'b0}},layer0[11][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_11[2] <= { {8{1'b0}},layer0[11][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_11[3] <= { {8{1'b0}},layer0[11][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_11[4] <= { {8{1'b0}},layer0[11][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_11[5] <= { {8{1'b0}},layer1[11][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_11[6] <= { {8{1'b0}},layer1[11][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_11[7] <= { {8{1'b0}},layer1[11][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_11[8] <= { {8{1'b0}},layer1[11][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_11[9] <= { {8{1'b0}},layer1[11][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_11[10] <= { {8{1'b0}},layer2[11][7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_11[11] <= { {8{1'b0}},layer2[11][15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_11[12] <= { {8{1'b0}},layer2[11][23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_11[13] <= { {8{1'b0}},layer2[11][31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_11[14] <= { {8{1'b0}},layer2[11][39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_11[15] <= { {8{1'b0}},layer3[11][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_11[16] <= { {8{1'b0}},layer3[11][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_11[17] <= { {8{1'b0}},layer3[11][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_11[18] <= { {8{1'b0}},layer3[11][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_11[19] <= { {8{1'b0}},layer3[11][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_11[20] <= { {8{1'b0}},layer4[11][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_11[21] <= { {8{1'b0}},layer4[11][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_11[22] <= { {8{1'b0}},layer4[11][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_11[23] <= { {8{1'b0}},layer4[11][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_11[24] <= { {8{1'b0}},layer4[11][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_11;
reg  [15:0]  kernel_img_sum_2_11;
reg  [15:0]  kernel_img_sum_3_11;
reg  [15:0]  kernel_img_sum_4_11;
reg  [15:0]  kernel_img_sum_5_11;
reg  [15:0]  kernel_img_sum_6_11;
reg  [15:0]  kernel_img_sum_7_11;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_11 <= kernel_img_mul_11[0] + kernel_img_mul_11[1] + kernel_img_mul_11[2] + kernel_img_mul_11[3] + kernel_img_mul_11[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_11 <= kernel_img_mul_11[5] + kernel_img_mul_11[6] + kernel_img_mul_11[7] + kernel_img_mul_11[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_11 <= kernel_img_mul_11[9] + kernel_img_mul_11[10] + kernel_img_mul_11[11] + kernel_img_mul_11[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_11 <= kernel_img_mul_11[13] + kernel_img_mul_11[14] + kernel_img_mul_11[15] + kernel_img_mul_11[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_11 <= kernel_img_mul_11[17] + kernel_img_mul_11[18] + kernel_img_mul_11[19] + kernel_img_mul_11[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_11 <= kernel_img_mul_11[21] + kernel_img_mul_11[22] + kernel_img_mul_11[23] + kernel_img_mul_11[24];
  end
end
always@(*) begin
  kernel_img_sum_7_11 = kernel_img_sum_1_11 + kernel_img_sum_2_11 + kernel_img_sum_3_11 + kernel_img_sum_4_11 + kernel_img_sum_5_11 + kernel_img_sum_6_11;
end
reg  [15:0]  kernel_img_mul_12[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_12[0] <= 'd0;
    kernel_img_mul_12[1] <= 'd0;
    kernel_img_mul_12[2] <= 'd0;
    kernel_img_mul_12[3] <= 'd0;
    kernel_img_mul_12[4] <= 'd0;
    kernel_img_mul_12[5] <= 'd0;
    kernel_img_mul_12[6] <= 'd0;
    kernel_img_mul_12[7] <= 'd0;
    kernel_img_mul_12[8] <= 'd0;
    kernel_img_mul_12[9] <= 'd0;
    kernel_img_mul_12[10] <= 'd0;
    kernel_img_mul_12[11] <= 'd0;
    kernel_img_mul_12[12] <= 'd0;
    kernel_img_mul_12[13] <= 'd0;
    kernel_img_mul_12[14] <= 'd0;
    kernel_img_mul_12[15] <= 'd0;
    kernel_img_mul_12[16] <= 'd0;
    kernel_img_mul_12[17] <= 'd0;
    kernel_img_mul_12[18] <= 'd0;
    kernel_img_mul_12[19] <= 'd0;
    kernel_img_mul_12[20] <= 'd0;
    kernel_img_mul_12[21] <= 'd0;
    kernel_img_mul_12[22] <= 'd0;
    kernel_img_mul_12[23] <= 'd0;
    kernel_img_mul_12[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_12[0] <= { {8{1'b0}},layer0[12][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_12[1] <= { {8{1'b0}},layer0[12][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_12[2] <= { {8{1'b0}},layer0[12][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_12[3] <= { {8{1'b0}},layer0[12][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_12[4] <= { {8{1'b0}},layer0[12][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_12[5] <= { {8{1'b0}},layer1[12][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_12[6] <= { {8{1'b0}},layer1[12][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_12[7] <= { {8{1'b0}},layer1[12][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_12[8] <= { {8{1'b0}},layer1[12][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_12[9] <= { {8{1'b0}},layer1[12][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_12[10] <= { {8{1'b0}},layer2[12][7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_12[11] <= { {8{1'b0}},layer2[12][15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_12[12] <= { {8{1'b0}},layer2[12][23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_12[13] <= { {8{1'b0}},layer2[12][31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_12[14] <= { {8{1'b0}},layer2[12][39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_12[15] <= { {8{1'b0}},layer3[12][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_12[16] <= { {8{1'b0}},layer3[12][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_12[17] <= { {8{1'b0}},layer3[12][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_12[18] <= { {8{1'b0}},layer3[12][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_12[19] <= { {8{1'b0}},layer3[12][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_12[20] <= { {8{1'b0}},layer4[12][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_12[21] <= { {8{1'b0}},layer4[12][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_12[22] <= { {8{1'b0}},layer4[12][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_12[23] <= { {8{1'b0}},layer4[12][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_12[24] <= { {8{1'b0}},layer4[12][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_12;
reg  [15:0]  kernel_img_sum_2_12;
reg  [15:0]  kernel_img_sum_3_12;
reg  [15:0]  kernel_img_sum_4_12;
reg  [15:0]  kernel_img_sum_5_12;
reg  [15:0]  kernel_img_sum_6_12;
reg  [15:0]  kernel_img_sum_7_12;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_12 <= kernel_img_mul_12[0] + kernel_img_mul_12[1] + kernel_img_mul_12[2] + kernel_img_mul_12[3] + kernel_img_mul_12[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_12 <= kernel_img_mul_12[5] + kernel_img_mul_12[6] + kernel_img_mul_12[7] + kernel_img_mul_12[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_12 <= kernel_img_mul_12[9] + kernel_img_mul_12[10] + kernel_img_mul_12[11] + kernel_img_mul_12[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_12 <= kernel_img_mul_12[13] + kernel_img_mul_12[14] + kernel_img_mul_12[15] + kernel_img_mul_12[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_12 <= kernel_img_mul_12[17] + kernel_img_mul_12[18] + kernel_img_mul_12[19] + kernel_img_mul_12[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_12 <= kernel_img_mul_12[21] + kernel_img_mul_12[22] + kernel_img_mul_12[23] + kernel_img_mul_12[24];
  end
end
always@(*) begin
  kernel_img_sum_7_12 = kernel_img_sum_1_12 + kernel_img_sum_2_12 + kernel_img_sum_3_12 + kernel_img_sum_4_12 + kernel_img_sum_5_12 + kernel_img_sum_6_12;
end
reg  [15:0]  kernel_img_mul_13[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_13[0] <= 'd0;
    kernel_img_mul_13[1] <= 'd0;
    kernel_img_mul_13[2] <= 'd0;
    kernel_img_mul_13[3] <= 'd0;
    kernel_img_mul_13[4] <= 'd0;
    kernel_img_mul_13[5] <= 'd0;
    kernel_img_mul_13[6] <= 'd0;
    kernel_img_mul_13[7] <= 'd0;
    kernel_img_mul_13[8] <= 'd0;
    kernel_img_mul_13[9] <= 'd0;
    kernel_img_mul_13[10] <= 'd0;
    kernel_img_mul_13[11] <= 'd0;
    kernel_img_mul_13[12] <= 'd0;
    kernel_img_mul_13[13] <= 'd0;
    kernel_img_mul_13[14] <= 'd0;
    kernel_img_mul_13[15] <= 'd0;
    kernel_img_mul_13[16] <= 'd0;
    kernel_img_mul_13[17] <= 'd0;
    kernel_img_mul_13[18] <= 'd0;
    kernel_img_mul_13[19] <= 'd0;
    kernel_img_mul_13[20] <= 'd0;
    kernel_img_mul_13[21] <= 'd0;
    kernel_img_mul_13[22] <= 'd0;
    kernel_img_mul_13[23] <= 'd0;
    kernel_img_mul_13[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_13[0] <= { {8{1'b0}},layer0[13][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_13[1] <= { {8{1'b0}},layer0[13][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_13[2] <= { {8{1'b0}},layer0[13][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_13[3] <= { {8{1'b0}},layer0[13][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_13[4] <= { {8{1'b0}},layer0[13][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_13[5] <= { {8{1'b0}},layer1[13][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_13[6] <= { {8{1'b0}},layer1[13][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_13[7] <= { {8{1'b0}},layer1[13][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_13[8] <= { {8{1'b0}},layer1[13][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_13[9] <= { {8{1'b0}},layer1[13][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_13[10] <= { {8{1'b0}},layer2[13][7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_13[11] <= { {8{1'b0}},layer2[13][15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_13[12] <= { {8{1'b0}},layer2[13][23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_13[13] <= { {8{1'b0}},layer2[13][31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_13[14] <= { {8{1'b0}},layer2[13][39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_13[15] <= { {8{1'b0}},layer3[13][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_13[16] <= { {8{1'b0}},layer3[13][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_13[17] <= { {8{1'b0}},layer3[13][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_13[18] <= { {8{1'b0}},layer3[13][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_13[19] <= { {8{1'b0}},layer3[13][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_13[20] <= { {8{1'b0}},layer4[13][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_13[21] <= { {8{1'b0}},layer4[13][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_13[22] <= { {8{1'b0}},layer4[13][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_13[23] <= { {8{1'b0}},layer4[13][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_13[24] <= { {8{1'b0}},layer4[13][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_13;
reg  [15:0]  kernel_img_sum_2_13;
reg  [15:0]  kernel_img_sum_3_13;
reg  [15:0]  kernel_img_sum_4_13;
reg  [15:0]  kernel_img_sum_5_13;
reg  [15:0]  kernel_img_sum_6_13;
reg  [15:0]  kernel_img_sum_7_13;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_13 <= kernel_img_mul_13[0] + kernel_img_mul_13[1] + kernel_img_mul_13[2] + kernel_img_mul_13[3] + kernel_img_mul_13[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_13 <= kernel_img_mul_13[5] + kernel_img_mul_13[6] + kernel_img_mul_13[7] + kernel_img_mul_13[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_13 <= kernel_img_mul_13[9] + kernel_img_mul_13[10] + kernel_img_mul_13[11] + kernel_img_mul_13[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_13 <= kernel_img_mul_13[13] + kernel_img_mul_13[14] + kernel_img_mul_13[15] + kernel_img_mul_13[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_13 <= kernel_img_mul_13[17] + kernel_img_mul_13[18] + kernel_img_mul_13[19] + kernel_img_mul_13[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_13 <= kernel_img_mul_13[21] + kernel_img_mul_13[22] + kernel_img_mul_13[23] + kernel_img_mul_13[24];
  end
end
always@(*) begin
  kernel_img_sum_7_13 = kernel_img_sum_1_13 + kernel_img_sum_2_13 + kernel_img_sum_3_13 + kernel_img_sum_4_13 + kernel_img_sum_5_13 + kernel_img_sum_6_13;
end
reg  [15:0]  kernel_img_mul_14[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_14[0] <= 'd0;
    kernel_img_mul_14[1] <= 'd0;
    kernel_img_mul_14[2] <= 'd0;
    kernel_img_mul_14[3] <= 'd0;
    kernel_img_mul_14[4] <= 'd0;
    kernel_img_mul_14[5] <= 'd0;
    kernel_img_mul_14[6] <= 'd0;
    kernel_img_mul_14[7] <= 'd0;
    kernel_img_mul_14[8] <= 'd0;
    kernel_img_mul_14[9] <= 'd0;
    kernel_img_mul_14[10] <= 'd0;
    kernel_img_mul_14[11] <= 'd0;
    kernel_img_mul_14[12] <= 'd0;
    kernel_img_mul_14[13] <= 'd0;
    kernel_img_mul_14[14] <= 'd0;
    kernel_img_mul_14[15] <= 'd0;
    kernel_img_mul_14[16] <= 'd0;
    kernel_img_mul_14[17] <= 'd0;
    kernel_img_mul_14[18] <= 'd0;
    kernel_img_mul_14[19] <= 'd0;
    kernel_img_mul_14[20] <= 'd0;
    kernel_img_mul_14[21] <= 'd0;
    kernel_img_mul_14[22] <= 'd0;
    kernel_img_mul_14[23] <= 'd0;
    kernel_img_mul_14[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_14[0] <= { {8{1'b0}},layer0[14][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_14[1] <= { {8{1'b0}},layer0[14][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_14[2] <= { {8{1'b0}},layer0[14][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_14[3] <= { {8{1'b0}},layer0[14][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_14[4] <= { {8{1'b0}},layer0[14][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_14[5] <= { {8{1'b0}},layer1[14][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_14[6] <= { {8{1'b0}},layer1[14][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_14[7] <= { {8{1'b0}},layer1[14][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_14[8] <= { {8{1'b0}},layer1[14][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_14[9] <= { {8{1'b0}},layer1[14][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_14[10] <= { {8{1'b0}},layer2[14][7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_14[11] <= { {8{1'b0}},layer2[14][15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_14[12] <= { {8{1'b0}},layer2[14][23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_14[13] <= { {8{1'b0}},layer2[14][31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_14[14] <= { {8{1'b0}},layer2[14][39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_14[15] <= { {8{1'b0}},layer3[14][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_14[16] <= { {8{1'b0}},layer3[14][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_14[17] <= { {8{1'b0}},layer3[14][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_14[18] <= { {8{1'b0}},layer3[14][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_14[19] <= { {8{1'b0}},layer3[14][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_14[20] <= { {8{1'b0}},layer4[14][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_14[21] <= { {8{1'b0}},layer4[14][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_14[22] <= { {8{1'b0}},layer4[14][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_14[23] <= { {8{1'b0}},layer4[14][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_14[24] <= { {8{1'b0}},layer4[14][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_14;
reg  [15:0]  kernel_img_sum_2_14;
reg  [15:0]  kernel_img_sum_3_14;
reg  [15:0]  kernel_img_sum_4_14;
reg  [15:0]  kernel_img_sum_5_14;
reg  [15:0]  kernel_img_sum_6_14;
reg  [15:0]  kernel_img_sum_7_14;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_14 <= kernel_img_mul_14[0] + kernel_img_mul_14[1] + kernel_img_mul_14[2] + kernel_img_mul_14[3] + kernel_img_mul_14[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_14 <= kernel_img_mul_14[5] + kernel_img_mul_14[6] + kernel_img_mul_14[7] + kernel_img_mul_14[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_14 <= kernel_img_mul_14[9] + kernel_img_mul_14[10] + kernel_img_mul_14[11] + kernel_img_mul_14[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_14 <= kernel_img_mul_14[13] + kernel_img_mul_14[14] + kernel_img_mul_14[15] + kernel_img_mul_14[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_14 <= kernel_img_mul_14[17] + kernel_img_mul_14[18] + kernel_img_mul_14[19] + kernel_img_mul_14[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_14 <= kernel_img_mul_14[21] + kernel_img_mul_14[22] + kernel_img_mul_14[23] + kernel_img_mul_14[24];
  end
end
always@(*) begin
  kernel_img_sum_7_14 = kernel_img_sum_1_14 + kernel_img_sum_2_14 + kernel_img_sum_3_14 + kernel_img_sum_4_14 + kernel_img_sum_5_14 + kernel_img_sum_6_14;
end
reg  [15:0]  kernel_img_mul_15[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_15[0] <= 'd0;
    kernel_img_mul_15[1] <= 'd0;
    kernel_img_mul_15[2] <= 'd0;
    kernel_img_mul_15[3] <= 'd0;
    kernel_img_mul_15[4] <= 'd0;
    kernel_img_mul_15[5] <= 'd0;
    kernel_img_mul_15[6] <= 'd0;
    kernel_img_mul_15[7] <= 'd0;
    kernel_img_mul_15[8] <= 'd0;
    kernel_img_mul_15[9] <= 'd0;
    kernel_img_mul_15[10] <= 'd0;
    kernel_img_mul_15[11] <= 'd0;
    kernel_img_mul_15[12] <= 'd0;
    kernel_img_mul_15[13] <= 'd0;
    kernel_img_mul_15[14] <= 'd0;
    kernel_img_mul_15[15] <= 'd0;
    kernel_img_mul_15[16] <= 'd0;
    kernel_img_mul_15[17] <= 'd0;
    kernel_img_mul_15[18] <= 'd0;
    kernel_img_mul_15[19] <= 'd0;
    kernel_img_mul_15[20] <= 'd0;
    kernel_img_mul_15[21] <= 'd0;
    kernel_img_mul_15[22] <= 'd0;
    kernel_img_mul_15[23] <= 'd0;
    kernel_img_mul_15[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_15[0] <= { {8{1'b0}},layer0[15][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_15[1] <= { {8{1'b0}},layer0[15][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_15[2] <= { {8{1'b0}},layer0[15][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_15[3] <= { {8{1'b0}},layer0[15][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_15[4] <= { {8{1'b0}},layer0[15][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_15[5] <= { {8{1'b0}},layer1[15][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_15[6] <= { {8{1'b0}},layer1[15][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_15[7] <= { {8{1'b0}},layer1[15][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_15[8] <= { {8{1'b0}},layer1[15][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_15[9] <= { {8{1'b0}},layer1[15][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_15[10] <= { {8{1'b0}},layer2[15][7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_15[11] <= { {8{1'b0}},layer2[15][15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_15[12] <= { {8{1'b0}},layer2[15][23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_15[13] <= { {8{1'b0}},layer2[15][31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_15[14] <= { {8{1'b0}},layer2[15][39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_15[15] <= { {8{1'b0}},layer3[15][7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_15[16] <= { {8{1'b0}},layer3[15][15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_15[17] <= { {8{1'b0}},layer3[15][23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_15[18] <= { {8{1'b0}},layer3[15][31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_15[19] <= { {8{1'b0}},layer3[15][39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_15[20] <= { {8{1'b0}},layer4[15][7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_15[21] <= { {8{1'b0}},layer4[15][15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_15[22] <= { {8{1'b0}},layer4[15][23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_15[23] <= { {8{1'b0}},layer4[15][31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_15[24] <= { {8{1'b0}},layer4[15][39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_15;
reg  [15:0]  kernel_img_sum_2_15;
reg  [15:0]  kernel_img_sum_3_15;
reg  [15:0]  kernel_img_sum_4_15;
reg  [15:0]  kernel_img_sum_5_15;
reg  [15:0]  kernel_img_sum_6_15;
reg  [15:0]  kernel_img_sum_7_15;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_15 <= kernel_img_mul_15[0] + kernel_img_mul_15[1] + kernel_img_mul_15[2] + kernel_img_mul_15[3] + kernel_img_mul_15[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_15 <= kernel_img_mul_15[5] + kernel_img_mul_15[6] + kernel_img_mul_15[7] + kernel_img_mul_15[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_15 <= kernel_img_mul_15[9] + kernel_img_mul_15[10] + kernel_img_mul_15[11] + kernel_img_mul_15[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_15 <= kernel_img_mul_15[13] + kernel_img_mul_15[14] + kernel_img_mul_15[15] + kernel_img_mul_15[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_15 <= kernel_img_mul_15[17] + kernel_img_mul_15[18] + kernel_img_mul_15[19] + kernel_img_mul_15[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_15 <= kernel_img_mul_15[21] + kernel_img_mul_15[22] + kernel_img_mul_15[23] + kernel_img_mul_15[24];
  end
end
always@(*) begin
  kernel_img_sum_7_15 = kernel_img_sum_1_15 + kernel_img_sum_2_15 + kernel_img_sum_3_15 + kernel_img_sum_4_15 + kernel_img_sum_5_15 + kernel_img_sum_6_15;
end
always @(posedge clk) begin
  if(!rst_n) begin
    blur_out[7:0] <= 'd0;
    blur_out[15:8] <= 'd0;
    blur_out[23:16] <= 'd0;
    blur_out[31:24] <= 'd0;
    blur_out[39:32] <= 'd0;
    blur_out[47:40] <= 'd0;
    blur_out[55:48] <= 'd0;
    blur_out[63:56] <= 'd0;
    blur_out[71:64] <= 'd0;
    blur_out[79:72] <= 'd0;
    blur_out[87:80] <= 'd0;
    blur_out[95:88] <= 'd0;
    blur_out[103:96] <= 'd0;
    blur_out[111:104] <= 'd0;
    blur_out[119:112] <= 'd0;
    blur_out[127:120] <= 'd0;
  end
  else if(current_state==ST_UPDATE) begin
    blur_out[7:0] <= kernel_img_sum_7_0[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[15:8] <= kernel_img_sum_7_1[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[23:16] <= kernel_img_sum_7_2[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[31:24] <= kernel_img_sum_7_3[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[39:32] <= kernel_img_sum_7_4[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[47:40] <= kernel_img_sum_7_5[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[55:48] <= kernel_img_sum_7_6[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[63:56] <= kernel_img_sum_7_7[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[71:64] <= kernel_img_sum_7_8[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[79:72] <= kernel_img_sum_7_9[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[87:80] <= kernel_img_sum_7_10[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[95:88] <= kernel_img_sum_7_11[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[103:96] <= kernel_img_sum_7_12[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[111:104] <= kernel_img_sum_7_13[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[119:112] <= kernel_img_sum_7_14[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[127:120] <= kernel_img_sum_7_15[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
  end
end

/*
 *  FSM
 *
 */
always @(posedge clk) begin
  if (!rst_n) begin
    current_state <= ST_MUX;    
  end
  else begin
    current_state <= next_state;
  end
end
always @(*) begin
  case(current_state)
    ST_MUX: begin
      if(start)
        next_state = ST_MUL;
      else
        next_state = ST_MUX;
    end
    ST_MUL: begin
      if(current_state==ST_MUL)
        next_state = ST_ADD;
      else 
        next_state = ST_MUL;
    end
    ST_ADD: begin
      if(current_state==ST_ADD)
        next_state = ST_UPDATE;
      else 
        next_state = ST_ADD;
    end
    ST_UPDATE: begin
      if(current_state==ST_UPDATE)
        next_state = ST_MUL;
      else 
        next_state = ST_UPDATE;
    end
    default:
      next_state = ST_MUL;
  endcase
end

endmodule