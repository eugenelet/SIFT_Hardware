module detect_keypoint(
  layer_0_0, /*img*/
  layer_0_1,
  layer_0_2,
  layer_1_0, /*Blur 0*/
  layer_1_1,
  layer_1_2,
  layer_2_0, /*Blur 1*/
  layer_2_1,
  layer_2_2,
  layer_3_0, /*Blur 2*/
  layer_3_1,
  layer_3_2,
  current_col,
  is_keypoint
);

input       [5119:0]   layer_0_0,
                       layer_0_1,
                       layer_0_2,
                       layer_1_0,
                       layer_1_1,
                       layer_1_2,
                       layer_2_0,
                       layer_2_1,
                       layer_2_2,
                       layer_3_0,
                       layer_3_1,
                       layer_3_2;
input       [9:0]      current_col;
output                 is_keypoint;

reg signed [8:0]  top_0[0:2]; // wire
reg signed [8:0]  top_1[0:2]; // wire
reg signed [8:0]  top_2[0:2]; // wire
reg signed [8:0]  mid_0[0:2]; // wire
reg signed [8:0]  mid_1[0:2]; // wire
reg signed [8:0]  mid_2[0:2]; // wire
reg signed [8:0]  btm_0[0:2]; // wire
reg signed [8:0]  btm_1[0:2]; // wire
reg signed [8:0]  btm_2[0:2]; // wire

always@(*) begin
  case(current_col)
    'd8: begin
      top_0[0] = {1'b0,layer_1_0[63:56]} - {1'b0, layer_0_0[63:56]};
      top_0[1] = {1'b0,layer_1_0[71:64]} - {1'b0, layer_0_0[71:64]};
      top_0[2] = {1'b0,layer_1_0[79:72]} - {1'b0, layer_0_0[79:72]};
      top_1[0] = {1'b0,layer_1_1[63:56]} - {1'b0, layer_0_1[63:56]};
      top_1[1] = {1'b0,layer_1_1[71:64]} - {1'b0, layer_0_1[71:64]};
      top_1[2] = {1'b0,layer_1_1[79:72]} - {1'b0, layer_0_1[79:72]};
      top_2[0] = {1'b0,layer_1_2[63:56]} - {1'b0, layer_0_2[63:56]};
      top_2[1] = {1'b0,layer_1_2[71:64]} - {1'b0, layer_0_2[71:64]};
      top_2[2] = {1'b0,layer_1_2[79:72]} - {1'b0, layer_0_2[79:72]};
      mid_0[0] = {1'b0,layer_2_0[63:56]} - {1'b0, layer_1_0[63:56]};
      mid_0[1] = {1'b0,layer_2_0[71:64]} - {1'b0, layer_1_0[71:64]};
      mid_0[2] = {1'b0,layer_2_0[79:72]} - {1'b0, layer_1_0[79:72]};
      mid_1[0] = {1'b0,layer_2_1[63:56]} - {1'b0, layer_1_1[63:56]};
      mid_1[1] = {1'b0,layer_2_1[71:64]} - {1'b0, layer_1_1[71:64]};
      mid_1[2] = {1'b0,layer_2_1[79:72]} - {1'b0, layer_1_1[79:72]};
      mid_2[0] = {1'b0,layer_2_2[63:56]} - {1'b0, layer_1_2[63:56]};
      mid_2[1] = {1'b0,layer_2_2[71:64]} - {1'b0, layer_1_2[71:64]};
      mid_2[2] = {1'b0,layer_2_2[79:72]} - {1'b0, layer_1_2[79:72]};
      btm_0[0] = {1'b0,layer_3_0[63:56]} - {1'b0, layer_2_0[63:56]};
      btm_0[1] = {1'b0,layer_3_0[71:64]} - {1'b0, layer_2_0[71:64]};
      btm_0[2] = {1'b0,layer_3_0[79:72]} - {1'b0, layer_2_0[79:72]};
      btm_1[0] = {1'b0,layer_3_1[63:56]} - {1'b0, layer_2_1[63:56]};
      btm_1[1] = {1'b0,layer_3_1[71:64]} - {1'b0, layer_2_1[71:64]};
      btm_1[2] = {1'b0,layer_3_1[79:72]} - {1'b0, layer_2_1[79:72]};
      btm_2[0] = {1'b0,layer_3_2[63:56]} - {1'b0, layer_2_2[63:56]};
      btm_2[1] = {1'b0,layer_3_2[71:64]} - {1'b0, layer_2_2[71:64]};
      btm_2[2] = {1'b0,layer_3_2[79:72]} - {1'b0, layer_2_2[79:72]};
    end
    'd9: begin
      top_0[0] = {1'b0,layer_1_0[71:64]} - {1'b0, layer_0_0[71:64]};
      top_0[1] = {1'b0,layer_1_0[79:72]} - {1'b0, layer_0_0[79:72]};
      top_0[2] = {1'b0,layer_1_0[87:80]} - {1'b0, layer_0_0[87:80]};
      top_1[0] = {1'b0,layer_1_1[71:64]} - {1'b0, layer_0_1[71:64]};
      top_1[1] = {1'b0,layer_1_1[79:72]} - {1'b0, layer_0_1[79:72]};
      top_1[2] = {1'b0,layer_1_1[87:80]} - {1'b0, layer_0_1[87:80]};
      top_2[0] = {1'b0,layer_1_2[71:64]} - {1'b0, layer_0_2[71:64]};
      top_2[1] = {1'b0,layer_1_2[79:72]} - {1'b0, layer_0_2[79:72]};
      top_2[2] = {1'b0,layer_1_2[87:80]} - {1'b0, layer_0_2[87:80]};
      mid_0[0] = {1'b0,layer_2_0[71:64]} - {1'b0, layer_1_0[71:64]};
      mid_0[1] = {1'b0,layer_2_0[79:72]} - {1'b0, layer_1_0[79:72]};
      mid_0[2] = {1'b0,layer_2_0[87:80]} - {1'b0, layer_1_0[87:80]};
      mid_1[0] = {1'b0,layer_2_1[71:64]} - {1'b0, layer_1_1[71:64]};
      mid_1[1] = {1'b0,layer_2_1[79:72]} - {1'b0, layer_1_1[79:72]};
      mid_1[2] = {1'b0,layer_2_1[87:80]} - {1'b0, layer_1_1[87:80]};
      mid_2[0] = {1'b0,layer_2_2[71:64]} - {1'b0, layer_1_2[71:64]};
      mid_2[1] = {1'b0,layer_2_2[79:72]} - {1'b0, layer_1_2[79:72]};
      mid_2[2] = {1'b0,layer_2_2[87:80]} - {1'b0, layer_1_2[87:80]};
      btm_0[0] = {1'b0,layer_3_0[71:64]} - {1'b0, layer_2_0[71:64]};
      btm_0[1] = {1'b0,layer_3_0[79:72]} - {1'b0, layer_2_0[79:72]};
      btm_0[2] = {1'b0,layer_3_0[87:80]} - {1'b0, layer_2_0[87:80]};
      btm_1[0] = {1'b0,layer_3_1[71:64]} - {1'b0, layer_2_1[71:64]};
      btm_1[1] = {1'b0,layer_3_1[79:72]} - {1'b0, layer_2_1[79:72]};
      btm_1[2] = {1'b0,layer_3_1[87:80]} - {1'b0, layer_2_1[87:80]};
      btm_2[0] = {1'b0,layer_3_2[71:64]} - {1'b0, layer_2_2[71:64]};
      btm_2[1] = {1'b0,layer_3_2[79:72]} - {1'b0, layer_2_2[79:72]};
      btm_2[2] = {1'b0,layer_3_2[87:80]} - {1'b0, layer_2_2[87:80]};
    end
    'd10: begin
      top_0[0] = {1'b0,layer_1_0[79:72]} - {1'b0, layer_0_0[79:72]};
      top_0[1] = {1'b0,layer_1_0[87:80]} - {1'b0, layer_0_0[87:80]};
      top_0[2] = {1'b0,layer_1_0[95:88]} - {1'b0, layer_0_0[95:88]};
      top_1[0] = {1'b0,layer_1_1[79:72]} - {1'b0, layer_0_1[79:72]};
      top_1[1] = {1'b0,layer_1_1[87:80]} - {1'b0, layer_0_1[87:80]};
      top_1[2] = {1'b0,layer_1_1[95:88]} - {1'b0, layer_0_1[95:88]};
      top_2[0] = {1'b0,layer_1_2[79:72]} - {1'b0, layer_0_2[79:72]};
      top_2[1] = {1'b0,layer_1_2[87:80]} - {1'b0, layer_0_2[87:80]};
      top_2[2] = {1'b0,layer_1_2[95:88]} - {1'b0, layer_0_2[95:88]};
      mid_0[0] = {1'b0,layer_2_0[79:72]} - {1'b0, layer_1_0[79:72]};
      mid_0[1] = {1'b0,layer_2_0[87:80]} - {1'b0, layer_1_0[87:80]};
      mid_0[2] = {1'b0,layer_2_0[95:88]} - {1'b0, layer_1_0[95:88]};
      mid_1[0] = {1'b0,layer_2_1[79:72]} - {1'b0, layer_1_1[79:72]};
      mid_1[1] = {1'b0,layer_2_1[87:80]} - {1'b0, layer_1_1[87:80]};
      mid_1[2] = {1'b0,layer_2_1[95:88]} - {1'b0, layer_1_1[95:88]};
      mid_2[0] = {1'b0,layer_2_2[79:72]} - {1'b0, layer_1_2[79:72]};
      mid_2[1] = {1'b0,layer_2_2[87:80]} - {1'b0, layer_1_2[87:80]};
      mid_2[2] = {1'b0,layer_2_2[95:88]} - {1'b0, layer_1_2[95:88]};
      btm_0[0] = {1'b0,layer_3_0[79:72]} - {1'b0, layer_2_0[79:72]};
      btm_0[1] = {1'b0,layer_3_0[87:80]} - {1'b0, layer_2_0[87:80]};
      btm_0[2] = {1'b0,layer_3_0[95:88]} - {1'b0, layer_2_0[95:88]};
      btm_1[0] = {1'b0,layer_3_1[79:72]} - {1'b0, layer_2_1[79:72]};
      btm_1[1] = {1'b0,layer_3_1[87:80]} - {1'b0, layer_2_1[87:80]};
      btm_1[2] = {1'b0,layer_3_1[95:88]} - {1'b0, layer_2_1[95:88]};
      btm_2[0] = {1'b0,layer_3_2[79:72]} - {1'b0, layer_2_2[79:72]};
      btm_2[1] = {1'b0,layer_3_2[87:80]} - {1'b0, layer_2_2[87:80]};
      btm_2[2] = {1'b0,layer_3_2[95:88]} - {1'b0, layer_2_2[95:88]};
    end
    'd11: begin
      top_0[0] = {1'b0,layer_1_0[87:80]} - {1'b0, layer_0_0[87:80]};
      top_0[1] = {1'b0,layer_1_0[95:88]} - {1'b0, layer_0_0[95:88]};
      top_0[2] = {1'b0,layer_1_0[103:96]} - {1'b0, layer_0_0[103:96]};
      top_1[0] = {1'b0,layer_1_1[87:80]} - {1'b0, layer_0_1[87:80]};
      top_1[1] = {1'b0,layer_1_1[95:88]} - {1'b0, layer_0_1[95:88]};
      top_1[2] = {1'b0,layer_1_1[103:96]} - {1'b0, layer_0_1[103:96]};
      top_2[0] = {1'b0,layer_1_2[87:80]} - {1'b0, layer_0_2[87:80]};
      top_2[1] = {1'b0,layer_1_2[95:88]} - {1'b0, layer_0_2[95:88]};
      top_2[2] = {1'b0,layer_1_2[103:96]} - {1'b0, layer_0_2[103:96]};
      mid_0[0] = {1'b0,layer_2_0[87:80]} - {1'b0, layer_1_0[87:80]};
      mid_0[1] = {1'b0,layer_2_0[95:88]} - {1'b0, layer_1_0[95:88]};
      mid_0[2] = {1'b0,layer_2_0[103:96]} - {1'b0, layer_1_0[103:96]};
      mid_1[0] = {1'b0,layer_2_1[87:80]} - {1'b0, layer_1_1[87:80]};
      mid_1[1] = {1'b0,layer_2_1[95:88]} - {1'b0, layer_1_1[95:88]};
      mid_1[2] = {1'b0,layer_2_1[103:96]} - {1'b0, layer_1_1[103:96]};
      mid_2[0] = {1'b0,layer_2_2[87:80]} - {1'b0, layer_1_2[87:80]};
      mid_2[1] = {1'b0,layer_2_2[95:88]} - {1'b0, layer_1_2[95:88]};
      mid_2[2] = {1'b0,layer_2_2[103:96]} - {1'b0, layer_1_2[103:96]};
      btm_0[0] = {1'b0,layer_3_0[87:80]} - {1'b0, layer_2_0[87:80]};
      btm_0[1] = {1'b0,layer_3_0[95:88]} - {1'b0, layer_2_0[95:88]};
      btm_0[2] = {1'b0,layer_3_0[103:96]} - {1'b0, layer_2_0[103:96]};
      btm_1[0] = {1'b0,layer_3_1[87:80]} - {1'b0, layer_2_1[87:80]};
      btm_1[1] = {1'b0,layer_3_1[95:88]} - {1'b0, layer_2_1[95:88]};
      btm_1[2] = {1'b0,layer_3_1[103:96]} - {1'b0, layer_2_1[103:96]};
      btm_2[0] = {1'b0,layer_3_2[87:80]} - {1'b0, layer_2_2[87:80]};
      btm_2[1] = {1'b0,layer_3_2[95:88]} - {1'b0, layer_2_2[95:88]};
      btm_2[2] = {1'b0,layer_3_2[103:96]} - {1'b0, layer_2_2[103:96]};
    end
    'd12: begin
      top_0[0] = {1'b0,layer_1_0[95:88]} - {1'b0, layer_0_0[95:88]};
      top_0[1] = {1'b0,layer_1_0[103:96]} - {1'b0, layer_0_0[103:96]};
      top_0[2] = {1'b0,layer_1_0[111:104]} - {1'b0, layer_0_0[111:104]};
      top_1[0] = {1'b0,layer_1_1[95:88]} - {1'b0, layer_0_1[95:88]};
      top_1[1] = {1'b0,layer_1_1[103:96]} - {1'b0, layer_0_1[103:96]};
      top_1[2] = {1'b0,layer_1_1[111:104]} - {1'b0, layer_0_1[111:104]};
      top_2[0] = {1'b0,layer_1_2[95:88]} - {1'b0, layer_0_2[95:88]};
      top_2[1] = {1'b0,layer_1_2[103:96]} - {1'b0, layer_0_2[103:96]};
      top_2[2] = {1'b0,layer_1_2[111:104]} - {1'b0, layer_0_2[111:104]};
      mid_0[0] = {1'b0,layer_2_0[95:88]} - {1'b0, layer_1_0[95:88]};
      mid_0[1] = {1'b0,layer_2_0[103:96]} - {1'b0, layer_1_0[103:96]};
      mid_0[2] = {1'b0,layer_2_0[111:104]} - {1'b0, layer_1_0[111:104]};
      mid_1[0] = {1'b0,layer_2_1[95:88]} - {1'b0, layer_1_1[95:88]};
      mid_1[1] = {1'b0,layer_2_1[103:96]} - {1'b0, layer_1_1[103:96]};
      mid_1[2] = {1'b0,layer_2_1[111:104]} - {1'b0, layer_1_1[111:104]};
      mid_2[0] = {1'b0,layer_2_2[95:88]} - {1'b0, layer_1_2[95:88]};
      mid_2[1] = {1'b0,layer_2_2[103:96]} - {1'b0, layer_1_2[103:96]};
      mid_2[2] = {1'b0,layer_2_2[111:104]} - {1'b0, layer_1_2[111:104]};
      btm_0[0] = {1'b0,layer_3_0[95:88]} - {1'b0, layer_2_0[95:88]};
      btm_0[1] = {1'b0,layer_3_0[103:96]} - {1'b0, layer_2_0[103:96]};
      btm_0[2] = {1'b0,layer_3_0[111:104]} - {1'b0, layer_2_0[111:104]};
      btm_1[0] = {1'b0,layer_3_1[95:88]} - {1'b0, layer_2_1[95:88]};
      btm_1[1] = {1'b0,layer_3_1[103:96]} - {1'b0, layer_2_1[103:96]};
      btm_1[2] = {1'b0,layer_3_1[111:104]} - {1'b0, layer_2_1[111:104]};
      btm_2[0] = {1'b0,layer_3_2[95:88]} - {1'b0, layer_2_2[95:88]};
      btm_2[1] = {1'b0,layer_3_2[103:96]} - {1'b0, layer_2_2[103:96]};
      btm_2[2] = {1'b0,layer_3_2[111:104]} - {1'b0, layer_2_2[111:104]};
    end
    'd13: begin
      top_0[0] = {1'b0,layer_1_0[103:96]} - {1'b0, layer_0_0[103:96]};
      top_0[1] = {1'b0,layer_1_0[111:104]} - {1'b0, layer_0_0[111:104]};
      top_0[2] = {1'b0,layer_1_0[119:112]} - {1'b0, layer_0_0[119:112]};
      top_1[0] = {1'b0,layer_1_1[103:96]} - {1'b0, layer_0_1[103:96]};
      top_1[1] = {1'b0,layer_1_1[111:104]} - {1'b0, layer_0_1[111:104]};
      top_1[2] = {1'b0,layer_1_1[119:112]} - {1'b0, layer_0_1[119:112]};
      top_2[0] = {1'b0,layer_1_2[103:96]} - {1'b0, layer_0_2[103:96]};
      top_2[1] = {1'b0,layer_1_2[111:104]} - {1'b0, layer_0_2[111:104]};
      top_2[2] = {1'b0,layer_1_2[119:112]} - {1'b0, layer_0_2[119:112]};
      mid_0[0] = {1'b0,layer_2_0[103:96]} - {1'b0, layer_1_0[103:96]};
      mid_0[1] = {1'b0,layer_2_0[111:104]} - {1'b0, layer_1_0[111:104]};
      mid_0[2] = {1'b0,layer_2_0[119:112]} - {1'b0, layer_1_0[119:112]};
      mid_1[0] = {1'b0,layer_2_1[103:96]} - {1'b0, layer_1_1[103:96]};
      mid_1[1] = {1'b0,layer_2_1[111:104]} - {1'b0, layer_1_1[111:104]};
      mid_1[2] = {1'b0,layer_2_1[119:112]} - {1'b0, layer_1_1[119:112]};
      mid_2[0] = {1'b0,layer_2_2[103:96]} - {1'b0, layer_1_2[103:96]};
      mid_2[1] = {1'b0,layer_2_2[111:104]} - {1'b0, layer_1_2[111:104]};
      mid_2[2] = {1'b0,layer_2_2[119:112]} - {1'b0, layer_1_2[119:112]};
      btm_0[0] = {1'b0,layer_3_0[103:96]} - {1'b0, layer_2_0[103:96]};
      btm_0[1] = {1'b0,layer_3_0[111:104]} - {1'b0, layer_2_0[111:104]};
      btm_0[2] = {1'b0,layer_3_0[119:112]} - {1'b0, layer_2_0[119:112]};
      btm_1[0] = {1'b0,layer_3_1[103:96]} - {1'b0, layer_2_1[103:96]};
      btm_1[1] = {1'b0,layer_3_1[111:104]} - {1'b0, layer_2_1[111:104]};
      btm_1[2] = {1'b0,layer_3_1[119:112]} - {1'b0, layer_2_1[119:112]};
      btm_2[0] = {1'b0,layer_3_2[103:96]} - {1'b0, layer_2_2[103:96]};
      btm_2[1] = {1'b0,layer_3_2[111:104]} - {1'b0, layer_2_2[111:104]};
      btm_2[2] = {1'b0,layer_3_2[119:112]} - {1'b0, layer_2_2[119:112]};
    end
    'd14: begin
      top_0[0] = {1'b0,layer_1_0[111:104]} - {1'b0, layer_0_0[111:104]};
      top_0[1] = {1'b0,layer_1_0[119:112]} - {1'b0, layer_0_0[119:112]};
      top_0[2] = {1'b0,layer_1_0[127:120]} - {1'b0, layer_0_0[127:120]};
      top_1[0] = {1'b0,layer_1_1[111:104]} - {1'b0, layer_0_1[111:104]};
      top_1[1] = {1'b0,layer_1_1[119:112]} - {1'b0, layer_0_1[119:112]};
      top_1[2] = {1'b0,layer_1_1[127:120]} - {1'b0, layer_0_1[127:120]};
      top_2[0] = {1'b0,layer_1_2[111:104]} - {1'b0, layer_0_2[111:104]};
      top_2[1] = {1'b0,layer_1_2[119:112]} - {1'b0, layer_0_2[119:112]};
      top_2[2] = {1'b0,layer_1_2[127:120]} - {1'b0, layer_0_2[127:120]};
      mid_0[0] = {1'b0,layer_2_0[111:104]} - {1'b0, layer_1_0[111:104]};
      mid_0[1] = {1'b0,layer_2_0[119:112]} - {1'b0, layer_1_0[119:112]};
      mid_0[2] = {1'b0,layer_2_0[127:120]} - {1'b0, layer_1_0[127:120]};
      mid_1[0] = {1'b0,layer_2_1[111:104]} - {1'b0, layer_1_1[111:104]};
      mid_1[1] = {1'b0,layer_2_1[119:112]} - {1'b0, layer_1_1[119:112]};
      mid_1[2] = {1'b0,layer_2_1[127:120]} - {1'b0, layer_1_1[127:120]};
      mid_2[0] = {1'b0,layer_2_2[111:104]} - {1'b0, layer_1_2[111:104]};
      mid_2[1] = {1'b0,layer_2_2[119:112]} - {1'b0, layer_1_2[119:112]};
      mid_2[2] = {1'b0,layer_2_2[127:120]} - {1'b0, layer_1_2[127:120]};
      btm_0[0] = {1'b0,layer_3_0[111:104]} - {1'b0, layer_2_0[111:104]};
      btm_0[1] = {1'b0,layer_3_0[119:112]} - {1'b0, layer_2_0[119:112]};
      btm_0[2] = {1'b0,layer_3_0[127:120]} - {1'b0, layer_2_0[127:120]};
      btm_1[0] = {1'b0,layer_3_1[111:104]} - {1'b0, layer_2_1[111:104]};
      btm_1[1] = {1'b0,layer_3_1[119:112]} - {1'b0, layer_2_1[119:112]};
      btm_1[2] = {1'b0,layer_3_1[127:120]} - {1'b0, layer_2_1[127:120]};
      btm_2[0] = {1'b0,layer_3_2[111:104]} - {1'b0, layer_2_2[111:104]};
      btm_2[1] = {1'b0,layer_3_2[119:112]} - {1'b0, layer_2_2[119:112]};
      btm_2[2] = {1'b0,layer_3_2[127:120]} - {1'b0, layer_2_2[127:120]};
    end
    'd15: begin
      top_0[0] = {1'b0,layer_1_0[119:112]} - {1'b0, layer_0_0[119:112]};
      top_0[1] = {1'b0,layer_1_0[127:120]} - {1'b0, layer_0_0[127:120]};
      top_0[2] = {1'b0,layer_1_0[135:128]} - {1'b0, layer_0_0[135:128]};
      top_1[0] = {1'b0,layer_1_1[119:112]} - {1'b0, layer_0_1[119:112]};
      top_1[1] = {1'b0,layer_1_1[127:120]} - {1'b0, layer_0_1[127:120]};
      top_1[2] = {1'b0,layer_1_1[135:128]} - {1'b0, layer_0_1[135:128]};
      top_2[0] = {1'b0,layer_1_2[119:112]} - {1'b0, layer_0_2[119:112]};
      top_2[1] = {1'b0,layer_1_2[127:120]} - {1'b0, layer_0_2[127:120]};
      top_2[2] = {1'b0,layer_1_2[135:128]} - {1'b0, layer_0_2[135:128]};
      mid_0[0] = {1'b0,layer_2_0[119:112]} - {1'b0, layer_1_0[119:112]};
      mid_0[1] = {1'b0,layer_2_0[127:120]} - {1'b0, layer_1_0[127:120]};
      mid_0[2] = {1'b0,layer_2_0[135:128]} - {1'b0, layer_1_0[135:128]};
      mid_1[0] = {1'b0,layer_2_1[119:112]} - {1'b0, layer_1_1[119:112]};
      mid_1[1] = {1'b0,layer_2_1[127:120]} - {1'b0, layer_1_1[127:120]};
      mid_1[2] = {1'b0,layer_2_1[135:128]} - {1'b0, layer_1_1[135:128]};
      mid_2[0] = {1'b0,layer_2_2[119:112]} - {1'b0, layer_1_2[119:112]};
      mid_2[1] = {1'b0,layer_2_2[127:120]} - {1'b0, layer_1_2[127:120]};
      mid_2[2] = {1'b0,layer_2_2[135:128]} - {1'b0, layer_1_2[135:128]};
      btm_0[0] = {1'b0,layer_3_0[119:112]} - {1'b0, layer_2_0[119:112]};
      btm_0[1] = {1'b0,layer_3_0[127:120]} - {1'b0, layer_2_0[127:120]};
      btm_0[2] = {1'b0,layer_3_0[135:128]} - {1'b0, layer_2_0[135:128]};
      btm_1[0] = {1'b0,layer_3_1[119:112]} - {1'b0, layer_2_1[119:112]};
      btm_1[1] = {1'b0,layer_3_1[127:120]} - {1'b0, layer_2_1[127:120]};
      btm_1[2] = {1'b0,layer_3_1[135:128]} - {1'b0, layer_2_1[135:128]};
      btm_2[0] = {1'b0,layer_3_2[119:112]} - {1'b0, layer_2_2[119:112]};
      btm_2[1] = {1'b0,layer_3_2[127:120]} - {1'b0, layer_2_2[127:120]};
      btm_2[2] = {1'b0,layer_3_2[135:128]} - {1'b0, layer_2_2[135:128]};
    end
    'd16: begin
      top_0[0] = {1'b0,layer_1_0[127:120]} - {1'b0, layer_0_0[127:120]};
      top_0[1] = {1'b0,layer_1_0[135:128]} - {1'b0, layer_0_0[135:128]};
      top_0[2] = {1'b0,layer_1_0[143:136]} - {1'b0, layer_0_0[143:136]};
      top_1[0] = {1'b0,layer_1_1[127:120]} - {1'b0, layer_0_1[127:120]};
      top_1[1] = {1'b0,layer_1_1[135:128]} - {1'b0, layer_0_1[135:128]};
      top_1[2] = {1'b0,layer_1_1[143:136]} - {1'b0, layer_0_1[143:136]};
      top_2[0] = {1'b0,layer_1_2[127:120]} - {1'b0, layer_0_2[127:120]};
      top_2[1] = {1'b0,layer_1_2[135:128]} - {1'b0, layer_0_2[135:128]};
      top_2[2] = {1'b0,layer_1_2[143:136]} - {1'b0, layer_0_2[143:136]};
      mid_0[0] = {1'b0,layer_2_0[127:120]} - {1'b0, layer_1_0[127:120]};
      mid_0[1] = {1'b0,layer_2_0[135:128]} - {1'b0, layer_1_0[135:128]};
      mid_0[2] = {1'b0,layer_2_0[143:136]} - {1'b0, layer_1_0[143:136]};
      mid_1[0] = {1'b0,layer_2_1[127:120]} - {1'b0, layer_1_1[127:120]};
      mid_1[1] = {1'b0,layer_2_1[135:128]} - {1'b0, layer_1_1[135:128]};
      mid_1[2] = {1'b0,layer_2_1[143:136]} - {1'b0, layer_1_1[143:136]};
      mid_2[0] = {1'b0,layer_2_2[127:120]} - {1'b0, layer_1_2[127:120]};
      mid_2[1] = {1'b0,layer_2_2[135:128]} - {1'b0, layer_1_2[135:128]};
      mid_2[2] = {1'b0,layer_2_2[143:136]} - {1'b0, layer_1_2[143:136]};
      btm_0[0] = {1'b0,layer_3_0[127:120]} - {1'b0, layer_2_0[127:120]};
      btm_0[1] = {1'b0,layer_3_0[135:128]} - {1'b0, layer_2_0[135:128]};
      btm_0[2] = {1'b0,layer_3_0[143:136]} - {1'b0, layer_2_0[143:136]};
      btm_1[0] = {1'b0,layer_3_1[127:120]} - {1'b0, layer_2_1[127:120]};
      btm_1[1] = {1'b0,layer_3_1[135:128]} - {1'b0, layer_2_1[135:128]};
      btm_1[2] = {1'b0,layer_3_1[143:136]} - {1'b0, layer_2_1[143:136]};
      btm_2[0] = {1'b0,layer_3_2[127:120]} - {1'b0, layer_2_2[127:120]};
      btm_2[1] = {1'b0,layer_3_2[135:128]} - {1'b0, layer_2_2[135:128]};
      btm_2[2] = {1'b0,layer_3_2[143:136]} - {1'b0, layer_2_2[143:136]};
    end
    'd17: begin
      top_0[0] = {1'b0,layer_1_0[135:128]} - {1'b0, layer_0_0[135:128]};
      top_0[1] = {1'b0,layer_1_0[143:136]} - {1'b0, layer_0_0[143:136]};
      top_0[2] = {1'b0,layer_1_0[151:144]} - {1'b0, layer_0_0[151:144]};
      top_1[0] = {1'b0,layer_1_1[135:128]} - {1'b0, layer_0_1[135:128]};
      top_1[1] = {1'b0,layer_1_1[143:136]} - {1'b0, layer_0_1[143:136]};
      top_1[2] = {1'b0,layer_1_1[151:144]} - {1'b0, layer_0_1[151:144]};
      top_2[0] = {1'b0,layer_1_2[135:128]} - {1'b0, layer_0_2[135:128]};
      top_2[1] = {1'b0,layer_1_2[143:136]} - {1'b0, layer_0_2[143:136]};
      top_2[2] = {1'b0,layer_1_2[151:144]} - {1'b0, layer_0_2[151:144]};
      mid_0[0] = {1'b0,layer_2_0[135:128]} - {1'b0, layer_1_0[135:128]};
      mid_0[1] = {1'b0,layer_2_0[143:136]} - {1'b0, layer_1_0[143:136]};
      mid_0[2] = {1'b0,layer_2_0[151:144]} - {1'b0, layer_1_0[151:144]};
      mid_1[0] = {1'b0,layer_2_1[135:128]} - {1'b0, layer_1_1[135:128]};
      mid_1[1] = {1'b0,layer_2_1[143:136]} - {1'b0, layer_1_1[143:136]};
      mid_1[2] = {1'b0,layer_2_1[151:144]} - {1'b0, layer_1_1[151:144]};
      mid_2[0] = {1'b0,layer_2_2[135:128]} - {1'b0, layer_1_2[135:128]};
      mid_2[1] = {1'b0,layer_2_2[143:136]} - {1'b0, layer_1_2[143:136]};
      mid_2[2] = {1'b0,layer_2_2[151:144]} - {1'b0, layer_1_2[151:144]};
      btm_0[0] = {1'b0,layer_3_0[135:128]} - {1'b0, layer_2_0[135:128]};
      btm_0[1] = {1'b0,layer_3_0[143:136]} - {1'b0, layer_2_0[143:136]};
      btm_0[2] = {1'b0,layer_3_0[151:144]} - {1'b0, layer_2_0[151:144]};
      btm_1[0] = {1'b0,layer_3_1[135:128]} - {1'b0, layer_2_1[135:128]};
      btm_1[1] = {1'b0,layer_3_1[143:136]} - {1'b0, layer_2_1[143:136]};
      btm_1[2] = {1'b0,layer_3_1[151:144]} - {1'b0, layer_2_1[151:144]};
      btm_2[0] = {1'b0,layer_3_2[135:128]} - {1'b0, layer_2_2[135:128]};
      btm_2[1] = {1'b0,layer_3_2[143:136]} - {1'b0, layer_2_2[143:136]};
      btm_2[2] = {1'b0,layer_3_2[151:144]} - {1'b0, layer_2_2[151:144]};
    end
    'd18: begin
      top_0[0] = {1'b0,layer_1_0[143:136]} - {1'b0, layer_0_0[143:136]};
      top_0[1] = {1'b0,layer_1_0[151:144]} - {1'b0, layer_0_0[151:144]};
      top_0[2] = {1'b0,layer_1_0[159:152]} - {1'b0, layer_0_0[159:152]};
      top_1[0] = {1'b0,layer_1_1[143:136]} - {1'b0, layer_0_1[143:136]};
      top_1[1] = {1'b0,layer_1_1[151:144]} - {1'b0, layer_0_1[151:144]};
      top_1[2] = {1'b0,layer_1_1[159:152]} - {1'b0, layer_0_1[159:152]};
      top_2[0] = {1'b0,layer_1_2[143:136]} - {1'b0, layer_0_2[143:136]};
      top_2[1] = {1'b0,layer_1_2[151:144]} - {1'b0, layer_0_2[151:144]};
      top_2[2] = {1'b0,layer_1_2[159:152]} - {1'b0, layer_0_2[159:152]};
      mid_0[0] = {1'b0,layer_2_0[143:136]} - {1'b0, layer_1_0[143:136]};
      mid_0[1] = {1'b0,layer_2_0[151:144]} - {1'b0, layer_1_0[151:144]};
      mid_0[2] = {1'b0,layer_2_0[159:152]} - {1'b0, layer_1_0[159:152]};
      mid_1[0] = {1'b0,layer_2_1[143:136]} - {1'b0, layer_1_1[143:136]};
      mid_1[1] = {1'b0,layer_2_1[151:144]} - {1'b0, layer_1_1[151:144]};
      mid_1[2] = {1'b0,layer_2_1[159:152]} - {1'b0, layer_1_1[159:152]};
      mid_2[0] = {1'b0,layer_2_2[143:136]} - {1'b0, layer_1_2[143:136]};
      mid_2[1] = {1'b0,layer_2_2[151:144]} - {1'b0, layer_1_2[151:144]};
      mid_2[2] = {1'b0,layer_2_2[159:152]} - {1'b0, layer_1_2[159:152]};
      btm_0[0] = {1'b0,layer_3_0[143:136]} - {1'b0, layer_2_0[143:136]};
      btm_0[1] = {1'b0,layer_3_0[151:144]} - {1'b0, layer_2_0[151:144]};
      btm_0[2] = {1'b0,layer_3_0[159:152]} - {1'b0, layer_2_0[159:152]};
      btm_1[0] = {1'b0,layer_3_1[143:136]} - {1'b0, layer_2_1[143:136]};
      btm_1[1] = {1'b0,layer_3_1[151:144]} - {1'b0, layer_2_1[151:144]};
      btm_1[2] = {1'b0,layer_3_1[159:152]} - {1'b0, layer_2_1[159:152]};
      btm_2[0] = {1'b0,layer_3_2[143:136]} - {1'b0, layer_2_2[143:136]};
      btm_2[1] = {1'b0,layer_3_2[151:144]} - {1'b0, layer_2_2[151:144]};
      btm_2[2] = {1'b0,layer_3_2[159:152]} - {1'b0, layer_2_2[159:152]};
    end
    'd19: begin
      top_0[0] = {1'b0,layer_1_0[151:144]} - {1'b0, layer_0_0[151:144]};
      top_0[1] = {1'b0,layer_1_0[159:152]} - {1'b0, layer_0_0[159:152]};
      top_0[2] = {1'b0,layer_1_0[167:160]} - {1'b0, layer_0_0[167:160]};
      top_1[0] = {1'b0,layer_1_1[151:144]} - {1'b0, layer_0_1[151:144]};
      top_1[1] = {1'b0,layer_1_1[159:152]} - {1'b0, layer_0_1[159:152]};
      top_1[2] = {1'b0,layer_1_1[167:160]} - {1'b0, layer_0_1[167:160]};
      top_2[0] = {1'b0,layer_1_2[151:144]} - {1'b0, layer_0_2[151:144]};
      top_2[1] = {1'b0,layer_1_2[159:152]} - {1'b0, layer_0_2[159:152]};
      top_2[2] = {1'b0,layer_1_2[167:160]} - {1'b0, layer_0_2[167:160]};
      mid_0[0] = {1'b0,layer_2_0[151:144]} - {1'b0, layer_1_0[151:144]};
      mid_0[1] = {1'b0,layer_2_0[159:152]} - {1'b0, layer_1_0[159:152]};
      mid_0[2] = {1'b0,layer_2_0[167:160]} - {1'b0, layer_1_0[167:160]};
      mid_1[0] = {1'b0,layer_2_1[151:144]} - {1'b0, layer_1_1[151:144]};
      mid_1[1] = {1'b0,layer_2_1[159:152]} - {1'b0, layer_1_1[159:152]};
      mid_1[2] = {1'b0,layer_2_1[167:160]} - {1'b0, layer_1_1[167:160]};
      mid_2[0] = {1'b0,layer_2_2[151:144]} - {1'b0, layer_1_2[151:144]};
      mid_2[1] = {1'b0,layer_2_2[159:152]} - {1'b0, layer_1_2[159:152]};
      mid_2[2] = {1'b0,layer_2_2[167:160]} - {1'b0, layer_1_2[167:160]};
      btm_0[0] = {1'b0,layer_3_0[151:144]} - {1'b0, layer_2_0[151:144]};
      btm_0[1] = {1'b0,layer_3_0[159:152]} - {1'b0, layer_2_0[159:152]};
      btm_0[2] = {1'b0,layer_3_0[167:160]} - {1'b0, layer_2_0[167:160]};
      btm_1[0] = {1'b0,layer_3_1[151:144]} - {1'b0, layer_2_1[151:144]};
      btm_1[1] = {1'b0,layer_3_1[159:152]} - {1'b0, layer_2_1[159:152]};
      btm_1[2] = {1'b0,layer_3_1[167:160]} - {1'b0, layer_2_1[167:160]};
      btm_2[0] = {1'b0,layer_3_2[151:144]} - {1'b0, layer_2_2[151:144]};
      btm_2[1] = {1'b0,layer_3_2[159:152]} - {1'b0, layer_2_2[159:152]};
      btm_2[2] = {1'b0,layer_3_2[167:160]} - {1'b0, layer_2_2[167:160]};
    end
    'd20: begin
      top_0[0] = {1'b0,layer_1_0[159:152]} - {1'b0, layer_0_0[159:152]};
      top_0[1] = {1'b0,layer_1_0[167:160]} - {1'b0, layer_0_0[167:160]};
      top_0[2] = {1'b0,layer_1_0[175:168]} - {1'b0, layer_0_0[175:168]};
      top_1[0] = {1'b0,layer_1_1[159:152]} - {1'b0, layer_0_1[159:152]};
      top_1[1] = {1'b0,layer_1_1[167:160]} - {1'b0, layer_0_1[167:160]};
      top_1[2] = {1'b0,layer_1_1[175:168]} - {1'b0, layer_0_1[175:168]};
      top_2[0] = {1'b0,layer_1_2[159:152]} - {1'b0, layer_0_2[159:152]};
      top_2[1] = {1'b0,layer_1_2[167:160]} - {1'b0, layer_0_2[167:160]};
      top_2[2] = {1'b0,layer_1_2[175:168]} - {1'b0, layer_0_2[175:168]};
      mid_0[0] = {1'b0,layer_2_0[159:152]} - {1'b0, layer_1_0[159:152]};
      mid_0[1] = {1'b0,layer_2_0[167:160]} - {1'b0, layer_1_0[167:160]};
      mid_0[2] = {1'b0,layer_2_0[175:168]} - {1'b0, layer_1_0[175:168]};
      mid_1[0] = {1'b0,layer_2_1[159:152]} - {1'b0, layer_1_1[159:152]};
      mid_1[1] = {1'b0,layer_2_1[167:160]} - {1'b0, layer_1_1[167:160]};
      mid_1[2] = {1'b0,layer_2_1[175:168]} - {1'b0, layer_1_1[175:168]};
      mid_2[0] = {1'b0,layer_2_2[159:152]} - {1'b0, layer_1_2[159:152]};
      mid_2[1] = {1'b0,layer_2_2[167:160]} - {1'b0, layer_1_2[167:160]};
      mid_2[2] = {1'b0,layer_2_2[175:168]} - {1'b0, layer_1_2[175:168]};
      btm_0[0] = {1'b0,layer_3_0[159:152]} - {1'b0, layer_2_0[159:152]};
      btm_0[1] = {1'b0,layer_3_0[167:160]} - {1'b0, layer_2_0[167:160]};
      btm_0[2] = {1'b0,layer_3_0[175:168]} - {1'b0, layer_2_0[175:168]};
      btm_1[0] = {1'b0,layer_3_1[159:152]} - {1'b0, layer_2_1[159:152]};
      btm_1[1] = {1'b0,layer_3_1[167:160]} - {1'b0, layer_2_1[167:160]};
      btm_1[2] = {1'b0,layer_3_1[175:168]} - {1'b0, layer_2_1[175:168]};
      btm_2[0] = {1'b0,layer_3_2[159:152]} - {1'b0, layer_2_2[159:152]};
      btm_2[1] = {1'b0,layer_3_2[167:160]} - {1'b0, layer_2_2[167:160]};
      btm_2[2] = {1'b0,layer_3_2[175:168]} - {1'b0, layer_2_2[175:168]};
    end
    'd21: begin
      top_0[0] = {1'b0,layer_1_0[167:160]} - {1'b0, layer_0_0[167:160]};
      top_0[1] = {1'b0,layer_1_0[175:168]} - {1'b0, layer_0_0[175:168]};
      top_0[2] = {1'b0,layer_1_0[183:176]} - {1'b0, layer_0_0[183:176]};
      top_1[0] = {1'b0,layer_1_1[167:160]} - {1'b0, layer_0_1[167:160]};
      top_1[1] = {1'b0,layer_1_1[175:168]} - {1'b0, layer_0_1[175:168]};
      top_1[2] = {1'b0,layer_1_1[183:176]} - {1'b0, layer_0_1[183:176]};
      top_2[0] = {1'b0,layer_1_2[167:160]} - {1'b0, layer_0_2[167:160]};
      top_2[1] = {1'b0,layer_1_2[175:168]} - {1'b0, layer_0_2[175:168]};
      top_2[2] = {1'b0,layer_1_2[183:176]} - {1'b0, layer_0_2[183:176]};
      mid_0[0] = {1'b0,layer_2_0[167:160]} - {1'b0, layer_1_0[167:160]};
      mid_0[1] = {1'b0,layer_2_0[175:168]} - {1'b0, layer_1_0[175:168]};
      mid_0[2] = {1'b0,layer_2_0[183:176]} - {1'b0, layer_1_0[183:176]};
      mid_1[0] = {1'b0,layer_2_1[167:160]} - {1'b0, layer_1_1[167:160]};
      mid_1[1] = {1'b0,layer_2_1[175:168]} - {1'b0, layer_1_1[175:168]};
      mid_1[2] = {1'b0,layer_2_1[183:176]} - {1'b0, layer_1_1[183:176]};
      mid_2[0] = {1'b0,layer_2_2[167:160]} - {1'b0, layer_1_2[167:160]};
      mid_2[1] = {1'b0,layer_2_2[175:168]} - {1'b0, layer_1_2[175:168]};
      mid_2[2] = {1'b0,layer_2_2[183:176]} - {1'b0, layer_1_2[183:176]};
      btm_0[0] = {1'b0,layer_3_0[167:160]} - {1'b0, layer_2_0[167:160]};
      btm_0[1] = {1'b0,layer_3_0[175:168]} - {1'b0, layer_2_0[175:168]};
      btm_0[2] = {1'b0,layer_3_0[183:176]} - {1'b0, layer_2_0[183:176]};
      btm_1[0] = {1'b0,layer_3_1[167:160]} - {1'b0, layer_2_1[167:160]};
      btm_1[1] = {1'b0,layer_3_1[175:168]} - {1'b0, layer_2_1[175:168]};
      btm_1[2] = {1'b0,layer_3_1[183:176]} - {1'b0, layer_2_1[183:176]};
      btm_2[0] = {1'b0,layer_3_2[167:160]} - {1'b0, layer_2_2[167:160]};
      btm_2[1] = {1'b0,layer_3_2[175:168]} - {1'b0, layer_2_2[175:168]};
      btm_2[2] = {1'b0,layer_3_2[183:176]} - {1'b0, layer_2_2[183:176]};
    end
    'd22: begin
      top_0[0] = {1'b0,layer_1_0[175:168]} - {1'b0, layer_0_0[175:168]};
      top_0[1] = {1'b0,layer_1_0[183:176]} - {1'b0, layer_0_0[183:176]};
      top_0[2] = {1'b0,layer_1_0[191:184]} - {1'b0, layer_0_0[191:184]};
      top_1[0] = {1'b0,layer_1_1[175:168]} - {1'b0, layer_0_1[175:168]};
      top_1[1] = {1'b0,layer_1_1[183:176]} - {1'b0, layer_0_1[183:176]};
      top_1[2] = {1'b0,layer_1_1[191:184]} - {1'b0, layer_0_1[191:184]};
      top_2[0] = {1'b0,layer_1_2[175:168]} - {1'b0, layer_0_2[175:168]};
      top_2[1] = {1'b0,layer_1_2[183:176]} - {1'b0, layer_0_2[183:176]};
      top_2[2] = {1'b0,layer_1_2[191:184]} - {1'b0, layer_0_2[191:184]};
      mid_0[0] = {1'b0,layer_2_0[175:168]} - {1'b0, layer_1_0[175:168]};
      mid_0[1] = {1'b0,layer_2_0[183:176]} - {1'b0, layer_1_0[183:176]};
      mid_0[2] = {1'b0,layer_2_0[191:184]} - {1'b0, layer_1_0[191:184]};
      mid_1[0] = {1'b0,layer_2_1[175:168]} - {1'b0, layer_1_1[175:168]};
      mid_1[1] = {1'b0,layer_2_1[183:176]} - {1'b0, layer_1_1[183:176]};
      mid_1[2] = {1'b0,layer_2_1[191:184]} - {1'b0, layer_1_1[191:184]};
      mid_2[0] = {1'b0,layer_2_2[175:168]} - {1'b0, layer_1_2[175:168]};
      mid_2[1] = {1'b0,layer_2_2[183:176]} - {1'b0, layer_1_2[183:176]};
      mid_2[2] = {1'b0,layer_2_2[191:184]} - {1'b0, layer_1_2[191:184]};
      btm_0[0] = {1'b0,layer_3_0[175:168]} - {1'b0, layer_2_0[175:168]};
      btm_0[1] = {1'b0,layer_3_0[183:176]} - {1'b0, layer_2_0[183:176]};
      btm_0[2] = {1'b0,layer_3_0[191:184]} - {1'b0, layer_2_0[191:184]};
      btm_1[0] = {1'b0,layer_3_1[175:168]} - {1'b0, layer_2_1[175:168]};
      btm_1[1] = {1'b0,layer_3_1[183:176]} - {1'b0, layer_2_1[183:176]};
      btm_1[2] = {1'b0,layer_3_1[191:184]} - {1'b0, layer_2_1[191:184]};
      btm_2[0] = {1'b0,layer_3_2[175:168]} - {1'b0, layer_2_2[175:168]};
      btm_2[1] = {1'b0,layer_3_2[183:176]} - {1'b0, layer_2_2[183:176]};
      btm_2[2] = {1'b0,layer_3_2[191:184]} - {1'b0, layer_2_2[191:184]};
    end
    'd23: begin
      top_0[0] = {1'b0,layer_1_0[183:176]} - {1'b0, layer_0_0[183:176]};
      top_0[1] = {1'b0,layer_1_0[191:184]} - {1'b0, layer_0_0[191:184]};
      top_0[2] = {1'b0,layer_1_0[199:192]} - {1'b0, layer_0_0[199:192]};
      top_1[0] = {1'b0,layer_1_1[183:176]} - {1'b0, layer_0_1[183:176]};
      top_1[1] = {1'b0,layer_1_1[191:184]} - {1'b0, layer_0_1[191:184]};
      top_1[2] = {1'b0,layer_1_1[199:192]} - {1'b0, layer_0_1[199:192]};
      top_2[0] = {1'b0,layer_1_2[183:176]} - {1'b0, layer_0_2[183:176]};
      top_2[1] = {1'b0,layer_1_2[191:184]} - {1'b0, layer_0_2[191:184]};
      top_2[2] = {1'b0,layer_1_2[199:192]} - {1'b0, layer_0_2[199:192]};
      mid_0[0] = {1'b0,layer_2_0[183:176]} - {1'b0, layer_1_0[183:176]};
      mid_0[1] = {1'b0,layer_2_0[191:184]} - {1'b0, layer_1_0[191:184]};
      mid_0[2] = {1'b0,layer_2_0[199:192]} - {1'b0, layer_1_0[199:192]};
      mid_1[0] = {1'b0,layer_2_1[183:176]} - {1'b0, layer_1_1[183:176]};
      mid_1[1] = {1'b0,layer_2_1[191:184]} - {1'b0, layer_1_1[191:184]};
      mid_1[2] = {1'b0,layer_2_1[199:192]} - {1'b0, layer_1_1[199:192]};
      mid_2[0] = {1'b0,layer_2_2[183:176]} - {1'b0, layer_1_2[183:176]};
      mid_2[1] = {1'b0,layer_2_2[191:184]} - {1'b0, layer_1_2[191:184]};
      mid_2[2] = {1'b0,layer_2_2[199:192]} - {1'b0, layer_1_2[199:192]};
      btm_0[0] = {1'b0,layer_3_0[183:176]} - {1'b0, layer_2_0[183:176]};
      btm_0[1] = {1'b0,layer_3_0[191:184]} - {1'b0, layer_2_0[191:184]};
      btm_0[2] = {1'b0,layer_3_0[199:192]} - {1'b0, layer_2_0[199:192]};
      btm_1[0] = {1'b0,layer_3_1[183:176]} - {1'b0, layer_2_1[183:176]};
      btm_1[1] = {1'b0,layer_3_1[191:184]} - {1'b0, layer_2_1[191:184]};
      btm_1[2] = {1'b0,layer_3_1[199:192]} - {1'b0, layer_2_1[199:192]};
      btm_2[0] = {1'b0,layer_3_2[183:176]} - {1'b0, layer_2_2[183:176]};
      btm_2[1] = {1'b0,layer_3_2[191:184]} - {1'b0, layer_2_2[191:184]};
      btm_2[2] = {1'b0,layer_3_2[199:192]} - {1'b0, layer_2_2[199:192]};
    end
    'd24: begin
      top_0[0] = {1'b0,layer_1_0[191:184]} - {1'b0, layer_0_0[191:184]};
      top_0[1] = {1'b0,layer_1_0[199:192]} - {1'b0, layer_0_0[199:192]};
      top_0[2] = {1'b0,layer_1_0[207:200]} - {1'b0, layer_0_0[207:200]};
      top_1[0] = {1'b0,layer_1_1[191:184]} - {1'b0, layer_0_1[191:184]};
      top_1[1] = {1'b0,layer_1_1[199:192]} - {1'b0, layer_0_1[199:192]};
      top_1[2] = {1'b0,layer_1_1[207:200]} - {1'b0, layer_0_1[207:200]};
      top_2[0] = {1'b0,layer_1_2[191:184]} - {1'b0, layer_0_2[191:184]};
      top_2[1] = {1'b0,layer_1_2[199:192]} - {1'b0, layer_0_2[199:192]};
      top_2[2] = {1'b0,layer_1_2[207:200]} - {1'b0, layer_0_2[207:200]};
      mid_0[0] = {1'b0,layer_2_0[191:184]} - {1'b0, layer_1_0[191:184]};
      mid_0[1] = {1'b0,layer_2_0[199:192]} - {1'b0, layer_1_0[199:192]};
      mid_0[2] = {1'b0,layer_2_0[207:200]} - {1'b0, layer_1_0[207:200]};
      mid_1[0] = {1'b0,layer_2_1[191:184]} - {1'b0, layer_1_1[191:184]};
      mid_1[1] = {1'b0,layer_2_1[199:192]} - {1'b0, layer_1_1[199:192]};
      mid_1[2] = {1'b0,layer_2_1[207:200]} - {1'b0, layer_1_1[207:200]};
      mid_2[0] = {1'b0,layer_2_2[191:184]} - {1'b0, layer_1_2[191:184]};
      mid_2[1] = {1'b0,layer_2_2[199:192]} - {1'b0, layer_1_2[199:192]};
      mid_2[2] = {1'b0,layer_2_2[207:200]} - {1'b0, layer_1_2[207:200]};
      btm_0[0] = {1'b0,layer_3_0[191:184]} - {1'b0, layer_2_0[191:184]};
      btm_0[1] = {1'b0,layer_3_0[199:192]} - {1'b0, layer_2_0[199:192]};
      btm_0[2] = {1'b0,layer_3_0[207:200]} - {1'b0, layer_2_0[207:200]};
      btm_1[0] = {1'b0,layer_3_1[191:184]} - {1'b0, layer_2_1[191:184]};
      btm_1[1] = {1'b0,layer_3_1[199:192]} - {1'b0, layer_2_1[199:192]};
      btm_1[2] = {1'b0,layer_3_1[207:200]} - {1'b0, layer_2_1[207:200]};
      btm_2[0] = {1'b0,layer_3_2[191:184]} - {1'b0, layer_2_2[191:184]};
      btm_2[1] = {1'b0,layer_3_2[199:192]} - {1'b0, layer_2_2[199:192]};
      btm_2[2] = {1'b0,layer_3_2[207:200]} - {1'b0, layer_2_2[207:200]};
    end
    'd25: begin
      top_0[0] = {1'b0,layer_1_0[199:192]} - {1'b0, layer_0_0[199:192]};
      top_0[1] = {1'b0,layer_1_0[207:200]} - {1'b0, layer_0_0[207:200]};
      top_0[2] = {1'b0,layer_1_0[215:208]} - {1'b0, layer_0_0[215:208]};
      top_1[0] = {1'b0,layer_1_1[199:192]} - {1'b0, layer_0_1[199:192]};
      top_1[1] = {1'b0,layer_1_1[207:200]} - {1'b0, layer_0_1[207:200]};
      top_1[2] = {1'b0,layer_1_1[215:208]} - {1'b0, layer_0_1[215:208]};
      top_2[0] = {1'b0,layer_1_2[199:192]} - {1'b0, layer_0_2[199:192]};
      top_2[1] = {1'b0,layer_1_2[207:200]} - {1'b0, layer_0_2[207:200]};
      top_2[2] = {1'b0,layer_1_2[215:208]} - {1'b0, layer_0_2[215:208]};
      mid_0[0] = {1'b0,layer_2_0[199:192]} - {1'b0, layer_1_0[199:192]};
      mid_0[1] = {1'b0,layer_2_0[207:200]} - {1'b0, layer_1_0[207:200]};
      mid_0[2] = {1'b0,layer_2_0[215:208]} - {1'b0, layer_1_0[215:208]};
      mid_1[0] = {1'b0,layer_2_1[199:192]} - {1'b0, layer_1_1[199:192]};
      mid_1[1] = {1'b0,layer_2_1[207:200]} - {1'b0, layer_1_1[207:200]};
      mid_1[2] = {1'b0,layer_2_1[215:208]} - {1'b0, layer_1_1[215:208]};
      mid_2[0] = {1'b0,layer_2_2[199:192]} - {1'b0, layer_1_2[199:192]};
      mid_2[1] = {1'b0,layer_2_2[207:200]} - {1'b0, layer_1_2[207:200]};
      mid_2[2] = {1'b0,layer_2_2[215:208]} - {1'b0, layer_1_2[215:208]};
      btm_0[0] = {1'b0,layer_3_0[199:192]} - {1'b0, layer_2_0[199:192]};
      btm_0[1] = {1'b0,layer_3_0[207:200]} - {1'b0, layer_2_0[207:200]};
      btm_0[2] = {1'b0,layer_3_0[215:208]} - {1'b0, layer_2_0[215:208]};
      btm_1[0] = {1'b0,layer_3_1[199:192]} - {1'b0, layer_2_1[199:192]};
      btm_1[1] = {1'b0,layer_3_1[207:200]} - {1'b0, layer_2_1[207:200]};
      btm_1[2] = {1'b0,layer_3_1[215:208]} - {1'b0, layer_2_1[215:208]};
      btm_2[0] = {1'b0,layer_3_2[199:192]} - {1'b0, layer_2_2[199:192]};
      btm_2[1] = {1'b0,layer_3_2[207:200]} - {1'b0, layer_2_2[207:200]};
      btm_2[2] = {1'b0,layer_3_2[215:208]} - {1'b0, layer_2_2[215:208]};
    end
    'd26: begin
      top_0[0] = {1'b0,layer_1_0[207:200]} - {1'b0, layer_0_0[207:200]};
      top_0[1] = {1'b0,layer_1_0[215:208]} - {1'b0, layer_0_0[215:208]};
      top_0[2] = {1'b0,layer_1_0[223:216]} - {1'b0, layer_0_0[223:216]};
      top_1[0] = {1'b0,layer_1_1[207:200]} - {1'b0, layer_0_1[207:200]};
      top_1[1] = {1'b0,layer_1_1[215:208]} - {1'b0, layer_0_1[215:208]};
      top_1[2] = {1'b0,layer_1_1[223:216]} - {1'b0, layer_0_1[223:216]};
      top_2[0] = {1'b0,layer_1_2[207:200]} - {1'b0, layer_0_2[207:200]};
      top_2[1] = {1'b0,layer_1_2[215:208]} - {1'b0, layer_0_2[215:208]};
      top_2[2] = {1'b0,layer_1_2[223:216]} - {1'b0, layer_0_2[223:216]};
      mid_0[0] = {1'b0,layer_2_0[207:200]} - {1'b0, layer_1_0[207:200]};
      mid_0[1] = {1'b0,layer_2_0[215:208]} - {1'b0, layer_1_0[215:208]};
      mid_0[2] = {1'b0,layer_2_0[223:216]} - {1'b0, layer_1_0[223:216]};
      mid_1[0] = {1'b0,layer_2_1[207:200]} - {1'b0, layer_1_1[207:200]};
      mid_1[1] = {1'b0,layer_2_1[215:208]} - {1'b0, layer_1_1[215:208]};
      mid_1[2] = {1'b0,layer_2_1[223:216]} - {1'b0, layer_1_1[223:216]};
      mid_2[0] = {1'b0,layer_2_2[207:200]} - {1'b0, layer_1_2[207:200]};
      mid_2[1] = {1'b0,layer_2_2[215:208]} - {1'b0, layer_1_2[215:208]};
      mid_2[2] = {1'b0,layer_2_2[223:216]} - {1'b0, layer_1_2[223:216]};
      btm_0[0] = {1'b0,layer_3_0[207:200]} - {1'b0, layer_2_0[207:200]};
      btm_0[1] = {1'b0,layer_3_0[215:208]} - {1'b0, layer_2_0[215:208]};
      btm_0[2] = {1'b0,layer_3_0[223:216]} - {1'b0, layer_2_0[223:216]};
      btm_1[0] = {1'b0,layer_3_1[207:200]} - {1'b0, layer_2_1[207:200]};
      btm_1[1] = {1'b0,layer_3_1[215:208]} - {1'b0, layer_2_1[215:208]};
      btm_1[2] = {1'b0,layer_3_1[223:216]} - {1'b0, layer_2_1[223:216]};
      btm_2[0] = {1'b0,layer_3_2[207:200]} - {1'b0, layer_2_2[207:200]};
      btm_2[1] = {1'b0,layer_3_2[215:208]} - {1'b0, layer_2_2[215:208]};
      btm_2[2] = {1'b0,layer_3_2[223:216]} - {1'b0, layer_2_2[223:216]};
    end
    'd27: begin
      top_0[0] = {1'b0,layer_1_0[215:208]} - {1'b0, layer_0_0[215:208]};
      top_0[1] = {1'b0,layer_1_0[223:216]} - {1'b0, layer_0_0[223:216]};
      top_0[2] = {1'b0,layer_1_0[231:224]} - {1'b0, layer_0_0[231:224]};
      top_1[0] = {1'b0,layer_1_1[215:208]} - {1'b0, layer_0_1[215:208]};
      top_1[1] = {1'b0,layer_1_1[223:216]} - {1'b0, layer_0_1[223:216]};
      top_1[2] = {1'b0,layer_1_1[231:224]} - {1'b0, layer_0_1[231:224]};
      top_2[0] = {1'b0,layer_1_2[215:208]} - {1'b0, layer_0_2[215:208]};
      top_2[1] = {1'b0,layer_1_2[223:216]} - {1'b0, layer_0_2[223:216]};
      top_2[2] = {1'b0,layer_1_2[231:224]} - {1'b0, layer_0_2[231:224]};
      mid_0[0] = {1'b0,layer_2_0[215:208]} - {1'b0, layer_1_0[215:208]};
      mid_0[1] = {1'b0,layer_2_0[223:216]} - {1'b0, layer_1_0[223:216]};
      mid_0[2] = {1'b0,layer_2_0[231:224]} - {1'b0, layer_1_0[231:224]};
      mid_1[0] = {1'b0,layer_2_1[215:208]} - {1'b0, layer_1_1[215:208]};
      mid_1[1] = {1'b0,layer_2_1[223:216]} - {1'b0, layer_1_1[223:216]};
      mid_1[2] = {1'b0,layer_2_1[231:224]} - {1'b0, layer_1_1[231:224]};
      mid_2[0] = {1'b0,layer_2_2[215:208]} - {1'b0, layer_1_2[215:208]};
      mid_2[1] = {1'b0,layer_2_2[223:216]} - {1'b0, layer_1_2[223:216]};
      mid_2[2] = {1'b0,layer_2_2[231:224]} - {1'b0, layer_1_2[231:224]};
      btm_0[0] = {1'b0,layer_3_0[215:208]} - {1'b0, layer_2_0[215:208]};
      btm_0[1] = {1'b0,layer_3_0[223:216]} - {1'b0, layer_2_0[223:216]};
      btm_0[2] = {1'b0,layer_3_0[231:224]} - {1'b0, layer_2_0[231:224]};
      btm_1[0] = {1'b0,layer_3_1[215:208]} - {1'b0, layer_2_1[215:208]};
      btm_1[1] = {1'b0,layer_3_1[223:216]} - {1'b0, layer_2_1[223:216]};
      btm_1[2] = {1'b0,layer_3_1[231:224]} - {1'b0, layer_2_1[231:224]};
      btm_2[0] = {1'b0,layer_3_2[215:208]} - {1'b0, layer_2_2[215:208]};
      btm_2[1] = {1'b0,layer_3_2[223:216]} - {1'b0, layer_2_2[223:216]};
      btm_2[2] = {1'b0,layer_3_2[231:224]} - {1'b0, layer_2_2[231:224]};
    end
    'd28: begin
      top_0[0] = {1'b0,layer_1_0[223:216]} - {1'b0, layer_0_0[223:216]};
      top_0[1] = {1'b0,layer_1_0[231:224]} - {1'b0, layer_0_0[231:224]};
      top_0[2] = {1'b0,layer_1_0[239:232]} - {1'b0, layer_0_0[239:232]};
      top_1[0] = {1'b0,layer_1_1[223:216]} - {1'b0, layer_0_1[223:216]};
      top_1[1] = {1'b0,layer_1_1[231:224]} - {1'b0, layer_0_1[231:224]};
      top_1[2] = {1'b0,layer_1_1[239:232]} - {1'b0, layer_0_1[239:232]};
      top_2[0] = {1'b0,layer_1_2[223:216]} - {1'b0, layer_0_2[223:216]};
      top_2[1] = {1'b0,layer_1_2[231:224]} - {1'b0, layer_0_2[231:224]};
      top_2[2] = {1'b0,layer_1_2[239:232]} - {1'b0, layer_0_2[239:232]};
      mid_0[0] = {1'b0,layer_2_0[223:216]} - {1'b0, layer_1_0[223:216]};
      mid_0[1] = {1'b0,layer_2_0[231:224]} - {1'b0, layer_1_0[231:224]};
      mid_0[2] = {1'b0,layer_2_0[239:232]} - {1'b0, layer_1_0[239:232]};
      mid_1[0] = {1'b0,layer_2_1[223:216]} - {1'b0, layer_1_1[223:216]};
      mid_1[1] = {1'b0,layer_2_1[231:224]} - {1'b0, layer_1_1[231:224]};
      mid_1[2] = {1'b0,layer_2_1[239:232]} - {1'b0, layer_1_1[239:232]};
      mid_2[0] = {1'b0,layer_2_2[223:216]} - {1'b0, layer_1_2[223:216]};
      mid_2[1] = {1'b0,layer_2_2[231:224]} - {1'b0, layer_1_2[231:224]};
      mid_2[2] = {1'b0,layer_2_2[239:232]} - {1'b0, layer_1_2[239:232]};
      btm_0[0] = {1'b0,layer_3_0[223:216]} - {1'b0, layer_2_0[223:216]};
      btm_0[1] = {1'b0,layer_3_0[231:224]} - {1'b0, layer_2_0[231:224]};
      btm_0[2] = {1'b0,layer_3_0[239:232]} - {1'b0, layer_2_0[239:232]};
      btm_1[0] = {1'b0,layer_3_1[223:216]} - {1'b0, layer_2_1[223:216]};
      btm_1[1] = {1'b0,layer_3_1[231:224]} - {1'b0, layer_2_1[231:224]};
      btm_1[2] = {1'b0,layer_3_1[239:232]} - {1'b0, layer_2_1[239:232]};
      btm_2[0] = {1'b0,layer_3_2[223:216]} - {1'b0, layer_2_2[223:216]};
      btm_2[1] = {1'b0,layer_3_2[231:224]} - {1'b0, layer_2_2[231:224]};
      btm_2[2] = {1'b0,layer_3_2[239:232]} - {1'b0, layer_2_2[239:232]};
    end
    'd29: begin
      top_0[0] = {1'b0,layer_1_0[231:224]} - {1'b0, layer_0_0[231:224]};
      top_0[1] = {1'b0,layer_1_0[239:232]} - {1'b0, layer_0_0[239:232]};
      top_0[2] = {1'b0,layer_1_0[247:240]} - {1'b0, layer_0_0[247:240]};
      top_1[0] = {1'b0,layer_1_1[231:224]} - {1'b0, layer_0_1[231:224]};
      top_1[1] = {1'b0,layer_1_1[239:232]} - {1'b0, layer_0_1[239:232]};
      top_1[2] = {1'b0,layer_1_1[247:240]} - {1'b0, layer_0_1[247:240]};
      top_2[0] = {1'b0,layer_1_2[231:224]} - {1'b0, layer_0_2[231:224]};
      top_2[1] = {1'b0,layer_1_2[239:232]} - {1'b0, layer_0_2[239:232]};
      top_2[2] = {1'b0,layer_1_2[247:240]} - {1'b0, layer_0_2[247:240]};
      mid_0[0] = {1'b0,layer_2_0[231:224]} - {1'b0, layer_1_0[231:224]};
      mid_0[1] = {1'b0,layer_2_0[239:232]} - {1'b0, layer_1_0[239:232]};
      mid_0[2] = {1'b0,layer_2_0[247:240]} - {1'b0, layer_1_0[247:240]};
      mid_1[0] = {1'b0,layer_2_1[231:224]} - {1'b0, layer_1_1[231:224]};
      mid_1[1] = {1'b0,layer_2_1[239:232]} - {1'b0, layer_1_1[239:232]};
      mid_1[2] = {1'b0,layer_2_1[247:240]} - {1'b0, layer_1_1[247:240]};
      mid_2[0] = {1'b0,layer_2_2[231:224]} - {1'b0, layer_1_2[231:224]};
      mid_2[1] = {1'b0,layer_2_2[239:232]} - {1'b0, layer_1_2[239:232]};
      mid_2[2] = {1'b0,layer_2_2[247:240]} - {1'b0, layer_1_2[247:240]};
      btm_0[0] = {1'b0,layer_3_0[231:224]} - {1'b0, layer_2_0[231:224]};
      btm_0[1] = {1'b0,layer_3_0[239:232]} - {1'b0, layer_2_0[239:232]};
      btm_0[2] = {1'b0,layer_3_0[247:240]} - {1'b0, layer_2_0[247:240]};
      btm_1[0] = {1'b0,layer_3_1[231:224]} - {1'b0, layer_2_1[231:224]};
      btm_1[1] = {1'b0,layer_3_1[239:232]} - {1'b0, layer_2_1[239:232]};
      btm_1[2] = {1'b0,layer_3_1[247:240]} - {1'b0, layer_2_1[247:240]};
      btm_2[0] = {1'b0,layer_3_2[231:224]} - {1'b0, layer_2_2[231:224]};
      btm_2[1] = {1'b0,layer_3_2[239:232]} - {1'b0, layer_2_2[239:232]};
      btm_2[2] = {1'b0,layer_3_2[247:240]} - {1'b0, layer_2_2[247:240]};
    end
    'd30: begin
      top_0[0] = {1'b0,layer_1_0[239:232]} - {1'b0, layer_0_0[239:232]};
      top_0[1] = {1'b0,layer_1_0[247:240]} - {1'b0, layer_0_0[247:240]};
      top_0[2] = {1'b0,layer_1_0[255:248]} - {1'b0, layer_0_0[255:248]};
      top_1[0] = {1'b0,layer_1_1[239:232]} - {1'b0, layer_0_1[239:232]};
      top_1[1] = {1'b0,layer_1_1[247:240]} - {1'b0, layer_0_1[247:240]};
      top_1[2] = {1'b0,layer_1_1[255:248]} - {1'b0, layer_0_1[255:248]};
      top_2[0] = {1'b0,layer_1_2[239:232]} - {1'b0, layer_0_2[239:232]};
      top_2[1] = {1'b0,layer_1_2[247:240]} - {1'b0, layer_0_2[247:240]};
      top_2[2] = {1'b0,layer_1_2[255:248]} - {1'b0, layer_0_2[255:248]};
      mid_0[0] = {1'b0,layer_2_0[239:232]} - {1'b0, layer_1_0[239:232]};
      mid_0[1] = {1'b0,layer_2_0[247:240]} - {1'b0, layer_1_0[247:240]};
      mid_0[2] = {1'b0,layer_2_0[255:248]} - {1'b0, layer_1_0[255:248]};
      mid_1[0] = {1'b0,layer_2_1[239:232]} - {1'b0, layer_1_1[239:232]};
      mid_1[1] = {1'b0,layer_2_1[247:240]} - {1'b0, layer_1_1[247:240]};
      mid_1[2] = {1'b0,layer_2_1[255:248]} - {1'b0, layer_1_1[255:248]};
      mid_2[0] = {1'b0,layer_2_2[239:232]} - {1'b0, layer_1_2[239:232]};
      mid_2[1] = {1'b0,layer_2_2[247:240]} - {1'b0, layer_1_2[247:240]};
      mid_2[2] = {1'b0,layer_2_2[255:248]} - {1'b0, layer_1_2[255:248]};
      btm_0[0] = {1'b0,layer_3_0[239:232]} - {1'b0, layer_2_0[239:232]};
      btm_0[1] = {1'b0,layer_3_0[247:240]} - {1'b0, layer_2_0[247:240]};
      btm_0[2] = {1'b0,layer_3_0[255:248]} - {1'b0, layer_2_0[255:248]};
      btm_1[0] = {1'b0,layer_3_1[239:232]} - {1'b0, layer_2_1[239:232]};
      btm_1[1] = {1'b0,layer_3_1[247:240]} - {1'b0, layer_2_1[247:240]};
      btm_1[2] = {1'b0,layer_3_1[255:248]} - {1'b0, layer_2_1[255:248]};
      btm_2[0] = {1'b0,layer_3_2[239:232]} - {1'b0, layer_2_2[239:232]};
      btm_2[1] = {1'b0,layer_3_2[247:240]} - {1'b0, layer_2_2[247:240]};
      btm_2[2] = {1'b0,layer_3_2[255:248]} - {1'b0, layer_2_2[255:248]};
    end
    'd31: begin
      top_0[0] = {1'b0,layer_1_0[247:240]} - {1'b0, layer_0_0[247:240]};
      top_0[1] = {1'b0,layer_1_0[255:248]} - {1'b0, layer_0_0[255:248]};
      top_0[2] = {1'b0,layer_1_0[263:256]} - {1'b0, layer_0_0[263:256]};
      top_1[0] = {1'b0,layer_1_1[247:240]} - {1'b0, layer_0_1[247:240]};
      top_1[1] = {1'b0,layer_1_1[255:248]} - {1'b0, layer_0_1[255:248]};
      top_1[2] = {1'b0,layer_1_1[263:256]} - {1'b0, layer_0_1[263:256]};
      top_2[0] = {1'b0,layer_1_2[247:240]} - {1'b0, layer_0_2[247:240]};
      top_2[1] = {1'b0,layer_1_2[255:248]} - {1'b0, layer_0_2[255:248]};
      top_2[2] = {1'b0,layer_1_2[263:256]} - {1'b0, layer_0_2[263:256]};
      mid_0[0] = {1'b0,layer_2_0[247:240]} - {1'b0, layer_1_0[247:240]};
      mid_0[1] = {1'b0,layer_2_0[255:248]} - {1'b0, layer_1_0[255:248]};
      mid_0[2] = {1'b0,layer_2_0[263:256]} - {1'b0, layer_1_0[263:256]};
      mid_1[0] = {1'b0,layer_2_1[247:240]} - {1'b0, layer_1_1[247:240]};
      mid_1[1] = {1'b0,layer_2_1[255:248]} - {1'b0, layer_1_1[255:248]};
      mid_1[2] = {1'b0,layer_2_1[263:256]} - {1'b0, layer_1_1[263:256]};
      mid_2[0] = {1'b0,layer_2_2[247:240]} - {1'b0, layer_1_2[247:240]};
      mid_2[1] = {1'b0,layer_2_2[255:248]} - {1'b0, layer_1_2[255:248]};
      mid_2[2] = {1'b0,layer_2_2[263:256]} - {1'b0, layer_1_2[263:256]};
      btm_0[0] = {1'b0,layer_3_0[247:240]} - {1'b0, layer_2_0[247:240]};
      btm_0[1] = {1'b0,layer_3_0[255:248]} - {1'b0, layer_2_0[255:248]};
      btm_0[2] = {1'b0,layer_3_0[263:256]} - {1'b0, layer_2_0[263:256]};
      btm_1[0] = {1'b0,layer_3_1[247:240]} - {1'b0, layer_2_1[247:240]};
      btm_1[1] = {1'b0,layer_3_1[255:248]} - {1'b0, layer_2_1[255:248]};
      btm_1[2] = {1'b0,layer_3_1[263:256]} - {1'b0, layer_2_1[263:256]};
      btm_2[0] = {1'b0,layer_3_2[247:240]} - {1'b0, layer_2_2[247:240]};
      btm_2[1] = {1'b0,layer_3_2[255:248]} - {1'b0, layer_2_2[255:248]};
      btm_2[2] = {1'b0,layer_3_2[263:256]} - {1'b0, layer_2_2[263:256]};
    end
    'd32: begin
      top_0[0] = {1'b0,layer_1_0[255:248]} - {1'b0, layer_0_0[255:248]};
      top_0[1] = {1'b0,layer_1_0[263:256]} - {1'b0, layer_0_0[263:256]};
      top_0[2] = {1'b0,layer_1_0[271:264]} - {1'b0, layer_0_0[271:264]};
      top_1[0] = {1'b0,layer_1_1[255:248]} - {1'b0, layer_0_1[255:248]};
      top_1[1] = {1'b0,layer_1_1[263:256]} - {1'b0, layer_0_1[263:256]};
      top_1[2] = {1'b0,layer_1_1[271:264]} - {1'b0, layer_0_1[271:264]};
      top_2[0] = {1'b0,layer_1_2[255:248]} - {1'b0, layer_0_2[255:248]};
      top_2[1] = {1'b0,layer_1_2[263:256]} - {1'b0, layer_0_2[263:256]};
      top_2[2] = {1'b0,layer_1_2[271:264]} - {1'b0, layer_0_2[271:264]};
      mid_0[0] = {1'b0,layer_2_0[255:248]} - {1'b0, layer_1_0[255:248]};
      mid_0[1] = {1'b0,layer_2_0[263:256]} - {1'b0, layer_1_0[263:256]};
      mid_0[2] = {1'b0,layer_2_0[271:264]} - {1'b0, layer_1_0[271:264]};
      mid_1[0] = {1'b0,layer_2_1[255:248]} - {1'b0, layer_1_1[255:248]};
      mid_1[1] = {1'b0,layer_2_1[263:256]} - {1'b0, layer_1_1[263:256]};
      mid_1[2] = {1'b0,layer_2_1[271:264]} - {1'b0, layer_1_1[271:264]};
      mid_2[0] = {1'b0,layer_2_2[255:248]} - {1'b0, layer_1_2[255:248]};
      mid_2[1] = {1'b0,layer_2_2[263:256]} - {1'b0, layer_1_2[263:256]};
      mid_2[2] = {1'b0,layer_2_2[271:264]} - {1'b0, layer_1_2[271:264]};
      btm_0[0] = {1'b0,layer_3_0[255:248]} - {1'b0, layer_2_0[255:248]};
      btm_0[1] = {1'b0,layer_3_0[263:256]} - {1'b0, layer_2_0[263:256]};
      btm_0[2] = {1'b0,layer_3_0[271:264]} - {1'b0, layer_2_0[271:264]};
      btm_1[0] = {1'b0,layer_3_1[255:248]} - {1'b0, layer_2_1[255:248]};
      btm_1[1] = {1'b0,layer_3_1[263:256]} - {1'b0, layer_2_1[263:256]};
      btm_1[2] = {1'b0,layer_3_1[271:264]} - {1'b0, layer_2_1[271:264]};
      btm_2[0] = {1'b0,layer_3_2[255:248]} - {1'b0, layer_2_2[255:248]};
      btm_2[1] = {1'b0,layer_3_2[263:256]} - {1'b0, layer_2_2[263:256]};
      btm_2[2] = {1'b0,layer_3_2[271:264]} - {1'b0, layer_2_2[271:264]};
    end
    'd33: begin
      top_0[0] = {1'b0,layer_1_0[263:256]} - {1'b0, layer_0_0[263:256]};
      top_0[1] = {1'b0,layer_1_0[271:264]} - {1'b0, layer_0_0[271:264]};
      top_0[2] = {1'b0,layer_1_0[279:272]} - {1'b0, layer_0_0[279:272]};
      top_1[0] = {1'b0,layer_1_1[263:256]} - {1'b0, layer_0_1[263:256]};
      top_1[1] = {1'b0,layer_1_1[271:264]} - {1'b0, layer_0_1[271:264]};
      top_1[2] = {1'b0,layer_1_1[279:272]} - {1'b0, layer_0_1[279:272]};
      top_2[0] = {1'b0,layer_1_2[263:256]} - {1'b0, layer_0_2[263:256]};
      top_2[1] = {1'b0,layer_1_2[271:264]} - {1'b0, layer_0_2[271:264]};
      top_2[2] = {1'b0,layer_1_2[279:272]} - {1'b0, layer_0_2[279:272]};
      mid_0[0] = {1'b0,layer_2_0[263:256]} - {1'b0, layer_1_0[263:256]};
      mid_0[1] = {1'b0,layer_2_0[271:264]} - {1'b0, layer_1_0[271:264]};
      mid_0[2] = {1'b0,layer_2_0[279:272]} - {1'b0, layer_1_0[279:272]};
      mid_1[0] = {1'b0,layer_2_1[263:256]} - {1'b0, layer_1_1[263:256]};
      mid_1[1] = {1'b0,layer_2_1[271:264]} - {1'b0, layer_1_1[271:264]};
      mid_1[2] = {1'b0,layer_2_1[279:272]} - {1'b0, layer_1_1[279:272]};
      mid_2[0] = {1'b0,layer_2_2[263:256]} - {1'b0, layer_1_2[263:256]};
      mid_2[1] = {1'b0,layer_2_2[271:264]} - {1'b0, layer_1_2[271:264]};
      mid_2[2] = {1'b0,layer_2_2[279:272]} - {1'b0, layer_1_2[279:272]};
      btm_0[0] = {1'b0,layer_3_0[263:256]} - {1'b0, layer_2_0[263:256]};
      btm_0[1] = {1'b0,layer_3_0[271:264]} - {1'b0, layer_2_0[271:264]};
      btm_0[2] = {1'b0,layer_3_0[279:272]} - {1'b0, layer_2_0[279:272]};
      btm_1[0] = {1'b0,layer_3_1[263:256]} - {1'b0, layer_2_1[263:256]};
      btm_1[1] = {1'b0,layer_3_1[271:264]} - {1'b0, layer_2_1[271:264]};
      btm_1[2] = {1'b0,layer_3_1[279:272]} - {1'b0, layer_2_1[279:272]};
      btm_2[0] = {1'b0,layer_3_2[263:256]} - {1'b0, layer_2_2[263:256]};
      btm_2[1] = {1'b0,layer_3_2[271:264]} - {1'b0, layer_2_2[271:264]};
      btm_2[2] = {1'b0,layer_3_2[279:272]} - {1'b0, layer_2_2[279:272]};
    end
    'd34: begin
      top_0[0] = {1'b0,layer_1_0[271:264]} - {1'b0, layer_0_0[271:264]};
      top_0[1] = {1'b0,layer_1_0[279:272]} - {1'b0, layer_0_0[279:272]};
      top_0[2] = {1'b0,layer_1_0[287:280]} - {1'b0, layer_0_0[287:280]};
      top_1[0] = {1'b0,layer_1_1[271:264]} - {1'b0, layer_0_1[271:264]};
      top_1[1] = {1'b0,layer_1_1[279:272]} - {1'b0, layer_0_1[279:272]};
      top_1[2] = {1'b0,layer_1_1[287:280]} - {1'b0, layer_0_1[287:280]};
      top_2[0] = {1'b0,layer_1_2[271:264]} - {1'b0, layer_0_2[271:264]};
      top_2[1] = {1'b0,layer_1_2[279:272]} - {1'b0, layer_0_2[279:272]};
      top_2[2] = {1'b0,layer_1_2[287:280]} - {1'b0, layer_0_2[287:280]};
      mid_0[0] = {1'b0,layer_2_0[271:264]} - {1'b0, layer_1_0[271:264]};
      mid_0[1] = {1'b0,layer_2_0[279:272]} - {1'b0, layer_1_0[279:272]};
      mid_0[2] = {1'b0,layer_2_0[287:280]} - {1'b0, layer_1_0[287:280]};
      mid_1[0] = {1'b0,layer_2_1[271:264]} - {1'b0, layer_1_1[271:264]};
      mid_1[1] = {1'b0,layer_2_1[279:272]} - {1'b0, layer_1_1[279:272]};
      mid_1[2] = {1'b0,layer_2_1[287:280]} - {1'b0, layer_1_1[287:280]};
      mid_2[0] = {1'b0,layer_2_2[271:264]} - {1'b0, layer_1_2[271:264]};
      mid_2[1] = {1'b0,layer_2_2[279:272]} - {1'b0, layer_1_2[279:272]};
      mid_2[2] = {1'b0,layer_2_2[287:280]} - {1'b0, layer_1_2[287:280]};
      btm_0[0] = {1'b0,layer_3_0[271:264]} - {1'b0, layer_2_0[271:264]};
      btm_0[1] = {1'b0,layer_3_0[279:272]} - {1'b0, layer_2_0[279:272]};
      btm_0[2] = {1'b0,layer_3_0[287:280]} - {1'b0, layer_2_0[287:280]};
      btm_1[0] = {1'b0,layer_3_1[271:264]} - {1'b0, layer_2_1[271:264]};
      btm_1[1] = {1'b0,layer_3_1[279:272]} - {1'b0, layer_2_1[279:272]};
      btm_1[2] = {1'b0,layer_3_1[287:280]} - {1'b0, layer_2_1[287:280]};
      btm_2[0] = {1'b0,layer_3_2[271:264]} - {1'b0, layer_2_2[271:264]};
      btm_2[1] = {1'b0,layer_3_2[279:272]} - {1'b0, layer_2_2[279:272]};
      btm_2[2] = {1'b0,layer_3_2[287:280]} - {1'b0, layer_2_2[287:280]};
    end
    'd35: begin
      top_0[0] = {1'b0,layer_1_0[279:272]} - {1'b0, layer_0_0[279:272]};
      top_0[1] = {1'b0,layer_1_0[287:280]} - {1'b0, layer_0_0[287:280]};
      top_0[2] = {1'b0,layer_1_0[295:288]} - {1'b0, layer_0_0[295:288]};
      top_1[0] = {1'b0,layer_1_1[279:272]} - {1'b0, layer_0_1[279:272]};
      top_1[1] = {1'b0,layer_1_1[287:280]} - {1'b0, layer_0_1[287:280]};
      top_1[2] = {1'b0,layer_1_1[295:288]} - {1'b0, layer_0_1[295:288]};
      top_2[0] = {1'b0,layer_1_2[279:272]} - {1'b0, layer_0_2[279:272]};
      top_2[1] = {1'b0,layer_1_2[287:280]} - {1'b0, layer_0_2[287:280]};
      top_2[2] = {1'b0,layer_1_2[295:288]} - {1'b0, layer_0_2[295:288]};
      mid_0[0] = {1'b0,layer_2_0[279:272]} - {1'b0, layer_1_0[279:272]};
      mid_0[1] = {1'b0,layer_2_0[287:280]} - {1'b0, layer_1_0[287:280]};
      mid_0[2] = {1'b0,layer_2_0[295:288]} - {1'b0, layer_1_0[295:288]};
      mid_1[0] = {1'b0,layer_2_1[279:272]} - {1'b0, layer_1_1[279:272]};
      mid_1[1] = {1'b0,layer_2_1[287:280]} - {1'b0, layer_1_1[287:280]};
      mid_1[2] = {1'b0,layer_2_1[295:288]} - {1'b0, layer_1_1[295:288]};
      mid_2[0] = {1'b0,layer_2_2[279:272]} - {1'b0, layer_1_2[279:272]};
      mid_2[1] = {1'b0,layer_2_2[287:280]} - {1'b0, layer_1_2[287:280]};
      mid_2[2] = {1'b0,layer_2_2[295:288]} - {1'b0, layer_1_2[295:288]};
      btm_0[0] = {1'b0,layer_3_0[279:272]} - {1'b0, layer_2_0[279:272]};
      btm_0[1] = {1'b0,layer_3_0[287:280]} - {1'b0, layer_2_0[287:280]};
      btm_0[2] = {1'b0,layer_3_0[295:288]} - {1'b0, layer_2_0[295:288]};
      btm_1[0] = {1'b0,layer_3_1[279:272]} - {1'b0, layer_2_1[279:272]};
      btm_1[1] = {1'b0,layer_3_1[287:280]} - {1'b0, layer_2_1[287:280]};
      btm_1[2] = {1'b0,layer_3_1[295:288]} - {1'b0, layer_2_1[295:288]};
      btm_2[0] = {1'b0,layer_3_2[279:272]} - {1'b0, layer_2_2[279:272]};
      btm_2[1] = {1'b0,layer_3_2[287:280]} - {1'b0, layer_2_2[287:280]};
      btm_2[2] = {1'b0,layer_3_2[295:288]} - {1'b0, layer_2_2[295:288]};
    end
    'd36: begin
      top_0[0] = {1'b0,layer_1_0[287:280]} - {1'b0, layer_0_0[287:280]};
      top_0[1] = {1'b0,layer_1_0[295:288]} - {1'b0, layer_0_0[295:288]};
      top_0[2] = {1'b0,layer_1_0[303:296]} - {1'b0, layer_0_0[303:296]};
      top_1[0] = {1'b0,layer_1_1[287:280]} - {1'b0, layer_0_1[287:280]};
      top_1[1] = {1'b0,layer_1_1[295:288]} - {1'b0, layer_0_1[295:288]};
      top_1[2] = {1'b0,layer_1_1[303:296]} - {1'b0, layer_0_1[303:296]};
      top_2[0] = {1'b0,layer_1_2[287:280]} - {1'b0, layer_0_2[287:280]};
      top_2[1] = {1'b0,layer_1_2[295:288]} - {1'b0, layer_0_2[295:288]};
      top_2[2] = {1'b0,layer_1_2[303:296]} - {1'b0, layer_0_2[303:296]};
      mid_0[0] = {1'b0,layer_2_0[287:280]} - {1'b0, layer_1_0[287:280]};
      mid_0[1] = {1'b0,layer_2_0[295:288]} - {1'b0, layer_1_0[295:288]};
      mid_0[2] = {1'b0,layer_2_0[303:296]} - {1'b0, layer_1_0[303:296]};
      mid_1[0] = {1'b0,layer_2_1[287:280]} - {1'b0, layer_1_1[287:280]};
      mid_1[1] = {1'b0,layer_2_1[295:288]} - {1'b0, layer_1_1[295:288]};
      mid_1[2] = {1'b0,layer_2_1[303:296]} - {1'b0, layer_1_1[303:296]};
      mid_2[0] = {1'b0,layer_2_2[287:280]} - {1'b0, layer_1_2[287:280]};
      mid_2[1] = {1'b0,layer_2_2[295:288]} - {1'b0, layer_1_2[295:288]};
      mid_2[2] = {1'b0,layer_2_2[303:296]} - {1'b0, layer_1_2[303:296]};
      btm_0[0] = {1'b0,layer_3_0[287:280]} - {1'b0, layer_2_0[287:280]};
      btm_0[1] = {1'b0,layer_3_0[295:288]} - {1'b0, layer_2_0[295:288]};
      btm_0[2] = {1'b0,layer_3_0[303:296]} - {1'b0, layer_2_0[303:296]};
      btm_1[0] = {1'b0,layer_3_1[287:280]} - {1'b0, layer_2_1[287:280]};
      btm_1[1] = {1'b0,layer_3_1[295:288]} - {1'b0, layer_2_1[295:288]};
      btm_1[2] = {1'b0,layer_3_1[303:296]} - {1'b0, layer_2_1[303:296]};
      btm_2[0] = {1'b0,layer_3_2[287:280]} - {1'b0, layer_2_2[287:280]};
      btm_2[1] = {1'b0,layer_3_2[295:288]} - {1'b0, layer_2_2[295:288]};
      btm_2[2] = {1'b0,layer_3_2[303:296]} - {1'b0, layer_2_2[303:296]};
    end
    'd37: begin
      top_0[0] = {1'b0,layer_1_0[295:288]} - {1'b0, layer_0_0[295:288]};
      top_0[1] = {1'b0,layer_1_0[303:296]} - {1'b0, layer_0_0[303:296]};
      top_0[2] = {1'b0,layer_1_0[311:304]} - {1'b0, layer_0_0[311:304]};
      top_1[0] = {1'b0,layer_1_1[295:288]} - {1'b0, layer_0_1[295:288]};
      top_1[1] = {1'b0,layer_1_1[303:296]} - {1'b0, layer_0_1[303:296]};
      top_1[2] = {1'b0,layer_1_1[311:304]} - {1'b0, layer_0_1[311:304]};
      top_2[0] = {1'b0,layer_1_2[295:288]} - {1'b0, layer_0_2[295:288]};
      top_2[1] = {1'b0,layer_1_2[303:296]} - {1'b0, layer_0_2[303:296]};
      top_2[2] = {1'b0,layer_1_2[311:304]} - {1'b0, layer_0_2[311:304]};
      mid_0[0] = {1'b0,layer_2_0[295:288]} - {1'b0, layer_1_0[295:288]};
      mid_0[1] = {1'b0,layer_2_0[303:296]} - {1'b0, layer_1_0[303:296]};
      mid_0[2] = {1'b0,layer_2_0[311:304]} - {1'b0, layer_1_0[311:304]};
      mid_1[0] = {1'b0,layer_2_1[295:288]} - {1'b0, layer_1_1[295:288]};
      mid_1[1] = {1'b0,layer_2_1[303:296]} - {1'b0, layer_1_1[303:296]};
      mid_1[2] = {1'b0,layer_2_1[311:304]} - {1'b0, layer_1_1[311:304]};
      mid_2[0] = {1'b0,layer_2_2[295:288]} - {1'b0, layer_1_2[295:288]};
      mid_2[1] = {1'b0,layer_2_2[303:296]} - {1'b0, layer_1_2[303:296]};
      mid_2[2] = {1'b0,layer_2_2[311:304]} - {1'b0, layer_1_2[311:304]};
      btm_0[0] = {1'b0,layer_3_0[295:288]} - {1'b0, layer_2_0[295:288]};
      btm_0[1] = {1'b0,layer_3_0[303:296]} - {1'b0, layer_2_0[303:296]};
      btm_0[2] = {1'b0,layer_3_0[311:304]} - {1'b0, layer_2_0[311:304]};
      btm_1[0] = {1'b0,layer_3_1[295:288]} - {1'b0, layer_2_1[295:288]};
      btm_1[1] = {1'b0,layer_3_1[303:296]} - {1'b0, layer_2_1[303:296]};
      btm_1[2] = {1'b0,layer_3_1[311:304]} - {1'b0, layer_2_1[311:304]};
      btm_2[0] = {1'b0,layer_3_2[295:288]} - {1'b0, layer_2_2[295:288]};
      btm_2[1] = {1'b0,layer_3_2[303:296]} - {1'b0, layer_2_2[303:296]};
      btm_2[2] = {1'b0,layer_3_2[311:304]} - {1'b0, layer_2_2[311:304]};
    end
    'd38: begin
      top_0[0] = {1'b0,layer_1_0[303:296]} - {1'b0, layer_0_0[303:296]};
      top_0[1] = {1'b0,layer_1_0[311:304]} - {1'b0, layer_0_0[311:304]};
      top_0[2] = {1'b0,layer_1_0[319:312]} - {1'b0, layer_0_0[319:312]};
      top_1[0] = {1'b0,layer_1_1[303:296]} - {1'b0, layer_0_1[303:296]};
      top_1[1] = {1'b0,layer_1_1[311:304]} - {1'b0, layer_0_1[311:304]};
      top_1[2] = {1'b0,layer_1_1[319:312]} - {1'b0, layer_0_1[319:312]};
      top_2[0] = {1'b0,layer_1_2[303:296]} - {1'b0, layer_0_2[303:296]};
      top_2[1] = {1'b0,layer_1_2[311:304]} - {1'b0, layer_0_2[311:304]};
      top_2[2] = {1'b0,layer_1_2[319:312]} - {1'b0, layer_0_2[319:312]};
      mid_0[0] = {1'b0,layer_2_0[303:296]} - {1'b0, layer_1_0[303:296]};
      mid_0[1] = {1'b0,layer_2_0[311:304]} - {1'b0, layer_1_0[311:304]};
      mid_0[2] = {1'b0,layer_2_0[319:312]} - {1'b0, layer_1_0[319:312]};
      mid_1[0] = {1'b0,layer_2_1[303:296]} - {1'b0, layer_1_1[303:296]};
      mid_1[1] = {1'b0,layer_2_1[311:304]} - {1'b0, layer_1_1[311:304]};
      mid_1[2] = {1'b0,layer_2_1[319:312]} - {1'b0, layer_1_1[319:312]};
      mid_2[0] = {1'b0,layer_2_2[303:296]} - {1'b0, layer_1_2[303:296]};
      mid_2[1] = {1'b0,layer_2_2[311:304]} - {1'b0, layer_1_2[311:304]};
      mid_2[2] = {1'b0,layer_2_2[319:312]} - {1'b0, layer_1_2[319:312]};
      btm_0[0] = {1'b0,layer_3_0[303:296]} - {1'b0, layer_2_0[303:296]};
      btm_0[1] = {1'b0,layer_3_0[311:304]} - {1'b0, layer_2_0[311:304]};
      btm_0[2] = {1'b0,layer_3_0[319:312]} - {1'b0, layer_2_0[319:312]};
      btm_1[0] = {1'b0,layer_3_1[303:296]} - {1'b0, layer_2_1[303:296]};
      btm_1[1] = {1'b0,layer_3_1[311:304]} - {1'b0, layer_2_1[311:304]};
      btm_1[2] = {1'b0,layer_3_1[319:312]} - {1'b0, layer_2_1[319:312]};
      btm_2[0] = {1'b0,layer_3_2[303:296]} - {1'b0, layer_2_2[303:296]};
      btm_2[1] = {1'b0,layer_3_2[311:304]} - {1'b0, layer_2_2[311:304]};
      btm_2[2] = {1'b0,layer_3_2[319:312]} - {1'b0, layer_2_2[319:312]};
    end
    'd39: begin
      top_0[0] = {1'b0,layer_1_0[311:304]} - {1'b0, layer_0_0[311:304]};
      top_0[1] = {1'b0,layer_1_0[319:312]} - {1'b0, layer_0_0[319:312]};
      top_0[2] = {1'b0,layer_1_0[327:320]} - {1'b0, layer_0_0[327:320]};
      top_1[0] = {1'b0,layer_1_1[311:304]} - {1'b0, layer_0_1[311:304]};
      top_1[1] = {1'b0,layer_1_1[319:312]} - {1'b0, layer_0_1[319:312]};
      top_1[2] = {1'b0,layer_1_1[327:320]} - {1'b0, layer_0_1[327:320]};
      top_2[0] = {1'b0,layer_1_2[311:304]} - {1'b0, layer_0_2[311:304]};
      top_2[1] = {1'b0,layer_1_2[319:312]} - {1'b0, layer_0_2[319:312]};
      top_2[2] = {1'b0,layer_1_2[327:320]} - {1'b0, layer_0_2[327:320]};
      mid_0[0] = {1'b0,layer_2_0[311:304]} - {1'b0, layer_1_0[311:304]};
      mid_0[1] = {1'b0,layer_2_0[319:312]} - {1'b0, layer_1_0[319:312]};
      mid_0[2] = {1'b0,layer_2_0[327:320]} - {1'b0, layer_1_0[327:320]};
      mid_1[0] = {1'b0,layer_2_1[311:304]} - {1'b0, layer_1_1[311:304]};
      mid_1[1] = {1'b0,layer_2_1[319:312]} - {1'b0, layer_1_1[319:312]};
      mid_1[2] = {1'b0,layer_2_1[327:320]} - {1'b0, layer_1_1[327:320]};
      mid_2[0] = {1'b0,layer_2_2[311:304]} - {1'b0, layer_1_2[311:304]};
      mid_2[1] = {1'b0,layer_2_2[319:312]} - {1'b0, layer_1_2[319:312]};
      mid_2[2] = {1'b0,layer_2_2[327:320]} - {1'b0, layer_1_2[327:320]};
      btm_0[0] = {1'b0,layer_3_0[311:304]} - {1'b0, layer_2_0[311:304]};
      btm_0[1] = {1'b0,layer_3_0[319:312]} - {1'b0, layer_2_0[319:312]};
      btm_0[2] = {1'b0,layer_3_0[327:320]} - {1'b0, layer_2_0[327:320]};
      btm_1[0] = {1'b0,layer_3_1[311:304]} - {1'b0, layer_2_1[311:304]};
      btm_1[1] = {1'b0,layer_3_1[319:312]} - {1'b0, layer_2_1[319:312]};
      btm_1[2] = {1'b0,layer_3_1[327:320]} - {1'b0, layer_2_1[327:320]};
      btm_2[0] = {1'b0,layer_3_2[311:304]} - {1'b0, layer_2_2[311:304]};
      btm_2[1] = {1'b0,layer_3_2[319:312]} - {1'b0, layer_2_2[319:312]};
      btm_2[2] = {1'b0,layer_3_2[327:320]} - {1'b0, layer_2_2[327:320]};
    end
    'd40: begin
      top_0[0] = {1'b0,layer_1_0[319:312]} - {1'b0, layer_0_0[319:312]};
      top_0[1] = {1'b0,layer_1_0[327:320]} - {1'b0, layer_0_0[327:320]};
      top_0[2] = {1'b0,layer_1_0[335:328]} - {1'b0, layer_0_0[335:328]};
      top_1[0] = {1'b0,layer_1_1[319:312]} - {1'b0, layer_0_1[319:312]};
      top_1[1] = {1'b0,layer_1_1[327:320]} - {1'b0, layer_0_1[327:320]};
      top_1[2] = {1'b0,layer_1_1[335:328]} - {1'b0, layer_0_1[335:328]};
      top_2[0] = {1'b0,layer_1_2[319:312]} - {1'b0, layer_0_2[319:312]};
      top_2[1] = {1'b0,layer_1_2[327:320]} - {1'b0, layer_0_2[327:320]};
      top_2[2] = {1'b0,layer_1_2[335:328]} - {1'b0, layer_0_2[335:328]};
      mid_0[0] = {1'b0,layer_2_0[319:312]} - {1'b0, layer_1_0[319:312]};
      mid_0[1] = {1'b0,layer_2_0[327:320]} - {1'b0, layer_1_0[327:320]};
      mid_0[2] = {1'b0,layer_2_0[335:328]} - {1'b0, layer_1_0[335:328]};
      mid_1[0] = {1'b0,layer_2_1[319:312]} - {1'b0, layer_1_1[319:312]};
      mid_1[1] = {1'b0,layer_2_1[327:320]} - {1'b0, layer_1_1[327:320]};
      mid_1[2] = {1'b0,layer_2_1[335:328]} - {1'b0, layer_1_1[335:328]};
      mid_2[0] = {1'b0,layer_2_2[319:312]} - {1'b0, layer_1_2[319:312]};
      mid_2[1] = {1'b0,layer_2_2[327:320]} - {1'b0, layer_1_2[327:320]};
      mid_2[2] = {1'b0,layer_2_2[335:328]} - {1'b0, layer_1_2[335:328]};
      btm_0[0] = {1'b0,layer_3_0[319:312]} - {1'b0, layer_2_0[319:312]};
      btm_0[1] = {1'b0,layer_3_0[327:320]} - {1'b0, layer_2_0[327:320]};
      btm_0[2] = {1'b0,layer_3_0[335:328]} - {1'b0, layer_2_0[335:328]};
      btm_1[0] = {1'b0,layer_3_1[319:312]} - {1'b0, layer_2_1[319:312]};
      btm_1[1] = {1'b0,layer_3_1[327:320]} - {1'b0, layer_2_1[327:320]};
      btm_1[2] = {1'b0,layer_3_1[335:328]} - {1'b0, layer_2_1[335:328]};
      btm_2[0] = {1'b0,layer_3_2[319:312]} - {1'b0, layer_2_2[319:312]};
      btm_2[1] = {1'b0,layer_3_2[327:320]} - {1'b0, layer_2_2[327:320]};
      btm_2[2] = {1'b0,layer_3_2[335:328]} - {1'b0, layer_2_2[335:328]};
    end
    'd41: begin
      top_0[0] = {1'b0,layer_1_0[327:320]} - {1'b0, layer_0_0[327:320]};
      top_0[1] = {1'b0,layer_1_0[335:328]} - {1'b0, layer_0_0[335:328]};
      top_0[2] = {1'b0,layer_1_0[343:336]} - {1'b0, layer_0_0[343:336]};
      top_1[0] = {1'b0,layer_1_1[327:320]} - {1'b0, layer_0_1[327:320]};
      top_1[1] = {1'b0,layer_1_1[335:328]} - {1'b0, layer_0_1[335:328]};
      top_1[2] = {1'b0,layer_1_1[343:336]} - {1'b0, layer_0_1[343:336]};
      top_2[0] = {1'b0,layer_1_2[327:320]} - {1'b0, layer_0_2[327:320]};
      top_2[1] = {1'b0,layer_1_2[335:328]} - {1'b0, layer_0_2[335:328]};
      top_2[2] = {1'b0,layer_1_2[343:336]} - {1'b0, layer_0_2[343:336]};
      mid_0[0] = {1'b0,layer_2_0[327:320]} - {1'b0, layer_1_0[327:320]};
      mid_0[1] = {1'b0,layer_2_0[335:328]} - {1'b0, layer_1_0[335:328]};
      mid_0[2] = {1'b0,layer_2_0[343:336]} - {1'b0, layer_1_0[343:336]};
      mid_1[0] = {1'b0,layer_2_1[327:320]} - {1'b0, layer_1_1[327:320]};
      mid_1[1] = {1'b0,layer_2_1[335:328]} - {1'b0, layer_1_1[335:328]};
      mid_1[2] = {1'b0,layer_2_1[343:336]} - {1'b0, layer_1_1[343:336]};
      mid_2[0] = {1'b0,layer_2_2[327:320]} - {1'b0, layer_1_2[327:320]};
      mid_2[1] = {1'b0,layer_2_2[335:328]} - {1'b0, layer_1_2[335:328]};
      mid_2[2] = {1'b0,layer_2_2[343:336]} - {1'b0, layer_1_2[343:336]};
      btm_0[0] = {1'b0,layer_3_0[327:320]} - {1'b0, layer_2_0[327:320]};
      btm_0[1] = {1'b0,layer_3_0[335:328]} - {1'b0, layer_2_0[335:328]};
      btm_0[2] = {1'b0,layer_3_0[343:336]} - {1'b0, layer_2_0[343:336]};
      btm_1[0] = {1'b0,layer_3_1[327:320]} - {1'b0, layer_2_1[327:320]};
      btm_1[1] = {1'b0,layer_3_1[335:328]} - {1'b0, layer_2_1[335:328]};
      btm_1[2] = {1'b0,layer_3_1[343:336]} - {1'b0, layer_2_1[343:336]};
      btm_2[0] = {1'b0,layer_3_2[327:320]} - {1'b0, layer_2_2[327:320]};
      btm_2[1] = {1'b0,layer_3_2[335:328]} - {1'b0, layer_2_2[335:328]};
      btm_2[2] = {1'b0,layer_3_2[343:336]} - {1'b0, layer_2_2[343:336]};
    end
    'd42: begin
      top_0[0] = {1'b0,layer_1_0[335:328]} - {1'b0, layer_0_0[335:328]};
      top_0[1] = {1'b0,layer_1_0[343:336]} - {1'b0, layer_0_0[343:336]};
      top_0[2] = {1'b0,layer_1_0[351:344]} - {1'b0, layer_0_0[351:344]};
      top_1[0] = {1'b0,layer_1_1[335:328]} - {1'b0, layer_0_1[335:328]};
      top_1[1] = {1'b0,layer_1_1[343:336]} - {1'b0, layer_0_1[343:336]};
      top_1[2] = {1'b0,layer_1_1[351:344]} - {1'b0, layer_0_1[351:344]};
      top_2[0] = {1'b0,layer_1_2[335:328]} - {1'b0, layer_0_2[335:328]};
      top_2[1] = {1'b0,layer_1_2[343:336]} - {1'b0, layer_0_2[343:336]};
      top_2[2] = {1'b0,layer_1_2[351:344]} - {1'b0, layer_0_2[351:344]};
      mid_0[0] = {1'b0,layer_2_0[335:328]} - {1'b0, layer_1_0[335:328]};
      mid_0[1] = {1'b0,layer_2_0[343:336]} - {1'b0, layer_1_0[343:336]};
      mid_0[2] = {1'b0,layer_2_0[351:344]} - {1'b0, layer_1_0[351:344]};
      mid_1[0] = {1'b0,layer_2_1[335:328]} - {1'b0, layer_1_1[335:328]};
      mid_1[1] = {1'b0,layer_2_1[343:336]} - {1'b0, layer_1_1[343:336]};
      mid_1[2] = {1'b0,layer_2_1[351:344]} - {1'b0, layer_1_1[351:344]};
      mid_2[0] = {1'b0,layer_2_2[335:328]} - {1'b0, layer_1_2[335:328]};
      mid_2[1] = {1'b0,layer_2_2[343:336]} - {1'b0, layer_1_2[343:336]};
      mid_2[2] = {1'b0,layer_2_2[351:344]} - {1'b0, layer_1_2[351:344]};
      btm_0[0] = {1'b0,layer_3_0[335:328]} - {1'b0, layer_2_0[335:328]};
      btm_0[1] = {1'b0,layer_3_0[343:336]} - {1'b0, layer_2_0[343:336]};
      btm_0[2] = {1'b0,layer_3_0[351:344]} - {1'b0, layer_2_0[351:344]};
      btm_1[0] = {1'b0,layer_3_1[335:328]} - {1'b0, layer_2_1[335:328]};
      btm_1[1] = {1'b0,layer_3_1[343:336]} - {1'b0, layer_2_1[343:336]};
      btm_1[2] = {1'b0,layer_3_1[351:344]} - {1'b0, layer_2_1[351:344]};
      btm_2[0] = {1'b0,layer_3_2[335:328]} - {1'b0, layer_2_2[335:328]};
      btm_2[1] = {1'b0,layer_3_2[343:336]} - {1'b0, layer_2_2[343:336]};
      btm_2[2] = {1'b0,layer_3_2[351:344]} - {1'b0, layer_2_2[351:344]};
    end
    'd43: begin
      top_0[0] = {1'b0,layer_1_0[343:336]} - {1'b0, layer_0_0[343:336]};
      top_0[1] = {1'b0,layer_1_0[351:344]} - {1'b0, layer_0_0[351:344]};
      top_0[2] = {1'b0,layer_1_0[359:352]} - {1'b0, layer_0_0[359:352]};
      top_1[0] = {1'b0,layer_1_1[343:336]} - {1'b0, layer_0_1[343:336]};
      top_1[1] = {1'b0,layer_1_1[351:344]} - {1'b0, layer_0_1[351:344]};
      top_1[2] = {1'b0,layer_1_1[359:352]} - {1'b0, layer_0_1[359:352]};
      top_2[0] = {1'b0,layer_1_2[343:336]} - {1'b0, layer_0_2[343:336]};
      top_2[1] = {1'b0,layer_1_2[351:344]} - {1'b0, layer_0_2[351:344]};
      top_2[2] = {1'b0,layer_1_2[359:352]} - {1'b0, layer_0_2[359:352]};
      mid_0[0] = {1'b0,layer_2_0[343:336]} - {1'b0, layer_1_0[343:336]};
      mid_0[1] = {1'b0,layer_2_0[351:344]} - {1'b0, layer_1_0[351:344]};
      mid_0[2] = {1'b0,layer_2_0[359:352]} - {1'b0, layer_1_0[359:352]};
      mid_1[0] = {1'b0,layer_2_1[343:336]} - {1'b0, layer_1_1[343:336]};
      mid_1[1] = {1'b0,layer_2_1[351:344]} - {1'b0, layer_1_1[351:344]};
      mid_1[2] = {1'b0,layer_2_1[359:352]} - {1'b0, layer_1_1[359:352]};
      mid_2[0] = {1'b0,layer_2_2[343:336]} - {1'b0, layer_1_2[343:336]};
      mid_2[1] = {1'b0,layer_2_2[351:344]} - {1'b0, layer_1_2[351:344]};
      mid_2[2] = {1'b0,layer_2_2[359:352]} - {1'b0, layer_1_2[359:352]};
      btm_0[0] = {1'b0,layer_3_0[343:336]} - {1'b0, layer_2_0[343:336]};
      btm_0[1] = {1'b0,layer_3_0[351:344]} - {1'b0, layer_2_0[351:344]};
      btm_0[2] = {1'b0,layer_3_0[359:352]} - {1'b0, layer_2_0[359:352]};
      btm_1[0] = {1'b0,layer_3_1[343:336]} - {1'b0, layer_2_1[343:336]};
      btm_1[1] = {1'b0,layer_3_1[351:344]} - {1'b0, layer_2_1[351:344]};
      btm_1[2] = {1'b0,layer_3_1[359:352]} - {1'b0, layer_2_1[359:352]};
      btm_2[0] = {1'b0,layer_3_2[343:336]} - {1'b0, layer_2_2[343:336]};
      btm_2[1] = {1'b0,layer_3_2[351:344]} - {1'b0, layer_2_2[351:344]};
      btm_2[2] = {1'b0,layer_3_2[359:352]} - {1'b0, layer_2_2[359:352]};
    end
    'd44: begin
      top_0[0] = {1'b0,layer_1_0[351:344]} - {1'b0, layer_0_0[351:344]};
      top_0[1] = {1'b0,layer_1_0[359:352]} - {1'b0, layer_0_0[359:352]};
      top_0[2] = {1'b0,layer_1_0[367:360]} - {1'b0, layer_0_0[367:360]};
      top_1[0] = {1'b0,layer_1_1[351:344]} - {1'b0, layer_0_1[351:344]};
      top_1[1] = {1'b0,layer_1_1[359:352]} - {1'b0, layer_0_1[359:352]};
      top_1[2] = {1'b0,layer_1_1[367:360]} - {1'b0, layer_0_1[367:360]};
      top_2[0] = {1'b0,layer_1_2[351:344]} - {1'b0, layer_0_2[351:344]};
      top_2[1] = {1'b0,layer_1_2[359:352]} - {1'b0, layer_0_2[359:352]};
      top_2[2] = {1'b0,layer_1_2[367:360]} - {1'b0, layer_0_2[367:360]};
      mid_0[0] = {1'b0,layer_2_0[351:344]} - {1'b0, layer_1_0[351:344]};
      mid_0[1] = {1'b0,layer_2_0[359:352]} - {1'b0, layer_1_0[359:352]};
      mid_0[2] = {1'b0,layer_2_0[367:360]} - {1'b0, layer_1_0[367:360]};
      mid_1[0] = {1'b0,layer_2_1[351:344]} - {1'b0, layer_1_1[351:344]};
      mid_1[1] = {1'b0,layer_2_1[359:352]} - {1'b0, layer_1_1[359:352]};
      mid_1[2] = {1'b0,layer_2_1[367:360]} - {1'b0, layer_1_1[367:360]};
      mid_2[0] = {1'b0,layer_2_2[351:344]} - {1'b0, layer_1_2[351:344]};
      mid_2[1] = {1'b0,layer_2_2[359:352]} - {1'b0, layer_1_2[359:352]};
      mid_2[2] = {1'b0,layer_2_2[367:360]} - {1'b0, layer_1_2[367:360]};
      btm_0[0] = {1'b0,layer_3_0[351:344]} - {1'b0, layer_2_0[351:344]};
      btm_0[1] = {1'b0,layer_3_0[359:352]} - {1'b0, layer_2_0[359:352]};
      btm_0[2] = {1'b0,layer_3_0[367:360]} - {1'b0, layer_2_0[367:360]};
      btm_1[0] = {1'b0,layer_3_1[351:344]} - {1'b0, layer_2_1[351:344]};
      btm_1[1] = {1'b0,layer_3_1[359:352]} - {1'b0, layer_2_1[359:352]};
      btm_1[2] = {1'b0,layer_3_1[367:360]} - {1'b0, layer_2_1[367:360]};
      btm_2[0] = {1'b0,layer_3_2[351:344]} - {1'b0, layer_2_2[351:344]};
      btm_2[1] = {1'b0,layer_3_2[359:352]} - {1'b0, layer_2_2[359:352]};
      btm_2[2] = {1'b0,layer_3_2[367:360]} - {1'b0, layer_2_2[367:360]};
    end
    'd45: begin
      top_0[0] = {1'b0,layer_1_0[359:352]} - {1'b0, layer_0_0[359:352]};
      top_0[1] = {1'b0,layer_1_0[367:360]} - {1'b0, layer_0_0[367:360]};
      top_0[2] = {1'b0,layer_1_0[375:368]} - {1'b0, layer_0_0[375:368]};
      top_1[0] = {1'b0,layer_1_1[359:352]} - {1'b0, layer_0_1[359:352]};
      top_1[1] = {1'b0,layer_1_1[367:360]} - {1'b0, layer_0_1[367:360]};
      top_1[2] = {1'b0,layer_1_1[375:368]} - {1'b0, layer_0_1[375:368]};
      top_2[0] = {1'b0,layer_1_2[359:352]} - {1'b0, layer_0_2[359:352]};
      top_2[1] = {1'b0,layer_1_2[367:360]} - {1'b0, layer_0_2[367:360]};
      top_2[2] = {1'b0,layer_1_2[375:368]} - {1'b0, layer_0_2[375:368]};
      mid_0[0] = {1'b0,layer_2_0[359:352]} - {1'b0, layer_1_0[359:352]};
      mid_0[1] = {1'b0,layer_2_0[367:360]} - {1'b0, layer_1_0[367:360]};
      mid_0[2] = {1'b0,layer_2_0[375:368]} - {1'b0, layer_1_0[375:368]};
      mid_1[0] = {1'b0,layer_2_1[359:352]} - {1'b0, layer_1_1[359:352]};
      mid_1[1] = {1'b0,layer_2_1[367:360]} - {1'b0, layer_1_1[367:360]};
      mid_1[2] = {1'b0,layer_2_1[375:368]} - {1'b0, layer_1_1[375:368]};
      mid_2[0] = {1'b0,layer_2_2[359:352]} - {1'b0, layer_1_2[359:352]};
      mid_2[1] = {1'b0,layer_2_2[367:360]} - {1'b0, layer_1_2[367:360]};
      mid_2[2] = {1'b0,layer_2_2[375:368]} - {1'b0, layer_1_2[375:368]};
      btm_0[0] = {1'b0,layer_3_0[359:352]} - {1'b0, layer_2_0[359:352]};
      btm_0[1] = {1'b0,layer_3_0[367:360]} - {1'b0, layer_2_0[367:360]};
      btm_0[2] = {1'b0,layer_3_0[375:368]} - {1'b0, layer_2_0[375:368]};
      btm_1[0] = {1'b0,layer_3_1[359:352]} - {1'b0, layer_2_1[359:352]};
      btm_1[1] = {1'b0,layer_3_1[367:360]} - {1'b0, layer_2_1[367:360]};
      btm_1[2] = {1'b0,layer_3_1[375:368]} - {1'b0, layer_2_1[375:368]};
      btm_2[0] = {1'b0,layer_3_2[359:352]} - {1'b0, layer_2_2[359:352]};
      btm_2[1] = {1'b0,layer_3_2[367:360]} - {1'b0, layer_2_2[367:360]};
      btm_2[2] = {1'b0,layer_3_2[375:368]} - {1'b0, layer_2_2[375:368]};
    end
    'd46: begin
      top_0[0] = {1'b0,layer_1_0[367:360]} - {1'b0, layer_0_0[367:360]};
      top_0[1] = {1'b0,layer_1_0[375:368]} - {1'b0, layer_0_0[375:368]};
      top_0[2] = {1'b0,layer_1_0[383:376]} - {1'b0, layer_0_0[383:376]};
      top_1[0] = {1'b0,layer_1_1[367:360]} - {1'b0, layer_0_1[367:360]};
      top_1[1] = {1'b0,layer_1_1[375:368]} - {1'b0, layer_0_1[375:368]};
      top_1[2] = {1'b0,layer_1_1[383:376]} - {1'b0, layer_0_1[383:376]};
      top_2[0] = {1'b0,layer_1_2[367:360]} - {1'b0, layer_0_2[367:360]};
      top_2[1] = {1'b0,layer_1_2[375:368]} - {1'b0, layer_0_2[375:368]};
      top_2[2] = {1'b0,layer_1_2[383:376]} - {1'b0, layer_0_2[383:376]};
      mid_0[0] = {1'b0,layer_2_0[367:360]} - {1'b0, layer_1_0[367:360]};
      mid_0[1] = {1'b0,layer_2_0[375:368]} - {1'b0, layer_1_0[375:368]};
      mid_0[2] = {1'b0,layer_2_0[383:376]} - {1'b0, layer_1_0[383:376]};
      mid_1[0] = {1'b0,layer_2_1[367:360]} - {1'b0, layer_1_1[367:360]};
      mid_1[1] = {1'b0,layer_2_1[375:368]} - {1'b0, layer_1_1[375:368]};
      mid_1[2] = {1'b0,layer_2_1[383:376]} - {1'b0, layer_1_1[383:376]};
      mid_2[0] = {1'b0,layer_2_2[367:360]} - {1'b0, layer_1_2[367:360]};
      mid_2[1] = {1'b0,layer_2_2[375:368]} - {1'b0, layer_1_2[375:368]};
      mid_2[2] = {1'b0,layer_2_2[383:376]} - {1'b0, layer_1_2[383:376]};
      btm_0[0] = {1'b0,layer_3_0[367:360]} - {1'b0, layer_2_0[367:360]};
      btm_0[1] = {1'b0,layer_3_0[375:368]} - {1'b0, layer_2_0[375:368]};
      btm_0[2] = {1'b0,layer_3_0[383:376]} - {1'b0, layer_2_0[383:376]};
      btm_1[0] = {1'b0,layer_3_1[367:360]} - {1'b0, layer_2_1[367:360]};
      btm_1[1] = {1'b0,layer_3_1[375:368]} - {1'b0, layer_2_1[375:368]};
      btm_1[2] = {1'b0,layer_3_1[383:376]} - {1'b0, layer_2_1[383:376]};
      btm_2[0] = {1'b0,layer_3_2[367:360]} - {1'b0, layer_2_2[367:360]};
      btm_2[1] = {1'b0,layer_3_2[375:368]} - {1'b0, layer_2_2[375:368]};
      btm_2[2] = {1'b0,layer_3_2[383:376]} - {1'b0, layer_2_2[383:376]};
    end
    'd47: begin
      top_0[0] = {1'b0,layer_1_0[375:368]} - {1'b0, layer_0_0[375:368]};
      top_0[1] = {1'b0,layer_1_0[383:376]} - {1'b0, layer_0_0[383:376]};
      top_0[2] = {1'b0,layer_1_0[391:384]} - {1'b0, layer_0_0[391:384]};
      top_1[0] = {1'b0,layer_1_1[375:368]} - {1'b0, layer_0_1[375:368]};
      top_1[1] = {1'b0,layer_1_1[383:376]} - {1'b0, layer_0_1[383:376]};
      top_1[2] = {1'b0,layer_1_1[391:384]} - {1'b0, layer_0_1[391:384]};
      top_2[0] = {1'b0,layer_1_2[375:368]} - {1'b0, layer_0_2[375:368]};
      top_2[1] = {1'b0,layer_1_2[383:376]} - {1'b0, layer_0_2[383:376]};
      top_2[2] = {1'b0,layer_1_2[391:384]} - {1'b0, layer_0_2[391:384]};
      mid_0[0] = {1'b0,layer_2_0[375:368]} - {1'b0, layer_1_0[375:368]};
      mid_0[1] = {1'b0,layer_2_0[383:376]} - {1'b0, layer_1_0[383:376]};
      mid_0[2] = {1'b0,layer_2_0[391:384]} - {1'b0, layer_1_0[391:384]};
      mid_1[0] = {1'b0,layer_2_1[375:368]} - {1'b0, layer_1_1[375:368]};
      mid_1[1] = {1'b0,layer_2_1[383:376]} - {1'b0, layer_1_1[383:376]};
      mid_1[2] = {1'b0,layer_2_1[391:384]} - {1'b0, layer_1_1[391:384]};
      mid_2[0] = {1'b0,layer_2_2[375:368]} - {1'b0, layer_1_2[375:368]};
      mid_2[1] = {1'b0,layer_2_2[383:376]} - {1'b0, layer_1_2[383:376]};
      mid_2[2] = {1'b0,layer_2_2[391:384]} - {1'b0, layer_1_2[391:384]};
      btm_0[0] = {1'b0,layer_3_0[375:368]} - {1'b0, layer_2_0[375:368]};
      btm_0[1] = {1'b0,layer_3_0[383:376]} - {1'b0, layer_2_0[383:376]};
      btm_0[2] = {1'b0,layer_3_0[391:384]} - {1'b0, layer_2_0[391:384]};
      btm_1[0] = {1'b0,layer_3_1[375:368]} - {1'b0, layer_2_1[375:368]};
      btm_1[1] = {1'b0,layer_3_1[383:376]} - {1'b0, layer_2_1[383:376]};
      btm_1[2] = {1'b0,layer_3_1[391:384]} - {1'b0, layer_2_1[391:384]};
      btm_2[0] = {1'b0,layer_3_2[375:368]} - {1'b0, layer_2_2[375:368]};
      btm_2[1] = {1'b0,layer_3_2[383:376]} - {1'b0, layer_2_2[383:376]};
      btm_2[2] = {1'b0,layer_3_2[391:384]} - {1'b0, layer_2_2[391:384]};
    end
    'd48: begin
      top_0[0] = {1'b0,layer_1_0[383:376]} - {1'b0, layer_0_0[383:376]};
      top_0[1] = {1'b0,layer_1_0[391:384]} - {1'b0, layer_0_0[391:384]};
      top_0[2] = {1'b0,layer_1_0[399:392]} - {1'b0, layer_0_0[399:392]};
      top_1[0] = {1'b0,layer_1_1[383:376]} - {1'b0, layer_0_1[383:376]};
      top_1[1] = {1'b0,layer_1_1[391:384]} - {1'b0, layer_0_1[391:384]};
      top_1[2] = {1'b0,layer_1_1[399:392]} - {1'b0, layer_0_1[399:392]};
      top_2[0] = {1'b0,layer_1_2[383:376]} - {1'b0, layer_0_2[383:376]};
      top_2[1] = {1'b0,layer_1_2[391:384]} - {1'b0, layer_0_2[391:384]};
      top_2[2] = {1'b0,layer_1_2[399:392]} - {1'b0, layer_0_2[399:392]};
      mid_0[0] = {1'b0,layer_2_0[383:376]} - {1'b0, layer_1_0[383:376]};
      mid_0[1] = {1'b0,layer_2_0[391:384]} - {1'b0, layer_1_0[391:384]};
      mid_0[2] = {1'b0,layer_2_0[399:392]} - {1'b0, layer_1_0[399:392]};
      mid_1[0] = {1'b0,layer_2_1[383:376]} - {1'b0, layer_1_1[383:376]};
      mid_1[1] = {1'b0,layer_2_1[391:384]} - {1'b0, layer_1_1[391:384]};
      mid_1[2] = {1'b0,layer_2_1[399:392]} - {1'b0, layer_1_1[399:392]};
      mid_2[0] = {1'b0,layer_2_2[383:376]} - {1'b0, layer_1_2[383:376]};
      mid_2[1] = {1'b0,layer_2_2[391:384]} - {1'b0, layer_1_2[391:384]};
      mid_2[2] = {1'b0,layer_2_2[399:392]} - {1'b0, layer_1_2[399:392]};
      btm_0[0] = {1'b0,layer_3_0[383:376]} - {1'b0, layer_2_0[383:376]};
      btm_0[1] = {1'b0,layer_3_0[391:384]} - {1'b0, layer_2_0[391:384]};
      btm_0[2] = {1'b0,layer_3_0[399:392]} - {1'b0, layer_2_0[399:392]};
      btm_1[0] = {1'b0,layer_3_1[383:376]} - {1'b0, layer_2_1[383:376]};
      btm_1[1] = {1'b0,layer_3_1[391:384]} - {1'b0, layer_2_1[391:384]};
      btm_1[2] = {1'b0,layer_3_1[399:392]} - {1'b0, layer_2_1[399:392]};
      btm_2[0] = {1'b0,layer_3_2[383:376]} - {1'b0, layer_2_2[383:376]};
      btm_2[1] = {1'b0,layer_3_2[391:384]} - {1'b0, layer_2_2[391:384]};
      btm_2[2] = {1'b0,layer_3_2[399:392]} - {1'b0, layer_2_2[399:392]};
    end
    'd49: begin
      top_0[0] = {1'b0,layer_1_0[391:384]} - {1'b0, layer_0_0[391:384]};
      top_0[1] = {1'b0,layer_1_0[399:392]} - {1'b0, layer_0_0[399:392]};
      top_0[2] = {1'b0,layer_1_0[407:400]} - {1'b0, layer_0_0[407:400]};
      top_1[0] = {1'b0,layer_1_1[391:384]} - {1'b0, layer_0_1[391:384]};
      top_1[1] = {1'b0,layer_1_1[399:392]} - {1'b0, layer_0_1[399:392]};
      top_1[2] = {1'b0,layer_1_1[407:400]} - {1'b0, layer_0_1[407:400]};
      top_2[0] = {1'b0,layer_1_2[391:384]} - {1'b0, layer_0_2[391:384]};
      top_2[1] = {1'b0,layer_1_2[399:392]} - {1'b0, layer_0_2[399:392]};
      top_2[2] = {1'b0,layer_1_2[407:400]} - {1'b0, layer_0_2[407:400]};
      mid_0[0] = {1'b0,layer_2_0[391:384]} - {1'b0, layer_1_0[391:384]};
      mid_0[1] = {1'b0,layer_2_0[399:392]} - {1'b0, layer_1_0[399:392]};
      mid_0[2] = {1'b0,layer_2_0[407:400]} - {1'b0, layer_1_0[407:400]};
      mid_1[0] = {1'b0,layer_2_1[391:384]} - {1'b0, layer_1_1[391:384]};
      mid_1[1] = {1'b0,layer_2_1[399:392]} - {1'b0, layer_1_1[399:392]};
      mid_1[2] = {1'b0,layer_2_1[407:400]} - {1'b0, layer_1_1[407:400]};
      mid_2[0] = {1'b0,layer_2_2[391:384]} - {1'b0, layer_1_2[391:384]};
      mid_2[1] = {1'b0,layer_2_2[399:392]} - {1'b0, layer_1_2[399:392]};
      mid_2[2] = {1'b0,layer_2_2[407:400]} - {1'b0, layer_1_2[407:400]};
      btm_0[0] = {1'b0,layer_3_0[391:384]} - {1'b0, layer_2_0[391:384]};
      btm_0[1] = {1'b0,layer_3_0[399:392]} - {1'b0, layer_2_0[399:392]};
      btm_0[2] = {1'b0,layer_3_0[407:400]} - {1'b0, layer_2_0[407:400]};
      btm_1[0] = {1'b0,layer_3_1[391:384]} - {1'b0, layer_2_1[391:384]};
      btm_1[1] = {1'b0,layer_3_1[399:392]} - {1'b0, layer_2_1[399:392]};
      btm_1[2] = {1'b0,layer_3_1[407:400]} - {1'b0, layer_2_1[407:400]};
      btm_2[0] = {1'b0,layer_3_2[391:384]} - {1'b0, layer_2_2[391:384]};
      btm_2[1] = {1'b0,layer_3_2[399:392]} - {1'b0, layer_2_2[399:392]};
      btm_2[2] = {1'b0,layer_3_2[407:400]} - {1'b0, layer_2_2[407:400]};
    end
    'd50: begin
      top_0[0] = {1'b0,layer_1_0[399:392]} - {1'b0, layer_0_0[399:392]};
      top_0[1] = {1'b0,layer_1_0[407:400]} - {1'b0, layer_0_0[407:400]};
      top_0[2] = {1'b0,layer_1_0[415:408]} - {1'b0, layer_0_0[415:408]};
      top_1[0] = {1'b0,layer_1_1[399:392]} - {1'b0, layer_0_1[399:392]};
      top_1[1] = {1'b0,layer_1_1[407:400]} - {1'b0, layer_0_1[407:400]};
      top_1[2] = {1'b0,layer_1_1[415:408]} - {1'b0, layer_0_1[415:408]};
      top_2[0] = {1'b0,layer_1_2[399:392]} - {1'b0, layer_0_2[399:392]};
      top_2[1] = {1'b0,layer_1_2[407:400]} - {1'b0, layer_0_2[407:400]};
      top_2[2] = {1'b0,layer_1_2[415:408]} - {1'b0, layer_0_2[415:408]};
      mid_0[0] = {1'b0,layer_2_0[399:392]} - {1'b0, layer_1_0[399:392]};
      mid_0[1] = {1'b0,layer_2_0[407:400]} - {1'b0, layer_1_0[407:400]};
      mid_0[2] = {1'b0,layer_2_0[415:408]} - {1'b0, layer_1_0[415:408]};
      mid_1[0] = {1'b0,layer_2_1[399:392]} - {1'b0, layer_1_1[399:392]};
      mid_1[1] = {1'b0,layer_2_1[407:400]} - {1'b0, layer_1_1[407:400]};
      mid_1[2] = {1'b0,layer_2_1[415:408]} - {1'b0, layer_1_1[415:408]};
      mid_2[0] = {1'b0,layer_2_2[399:392]} - {1'b0, layer_1_2[399:392]};
      mid_2[1] = {1'b0,layer_2_2[407:400]} - {1'b0, layer_1_2[407:400]};
      mid_2[2] = {1'b0,layer_2_2[415:408]} - {1'b0, layer_1_2[415:408]};
      btm_0[0] = {1'b0,layer_3_0[399:392]} - {1'b0, layer_2_0[399:392]};
      btm_0[1] = {1'b0,layer_3_0[407:400]} - {1'b0, layer_2_0[407:400]};
      btm_0[2] = {1'b0,layer_3_0[415:408]} - {1'b0, layer_2_0[415:408]};
      btm_1[0] = {1'b0,layer_3_1[399:392]} - {1'b0, layer_2_1[399:392]};
      btm_1[1] = {1'b0,layer_3_1[407:400]} - {1'b0, layer_2_1[407:400]};
      btm_1[2] = {1'b0,layer_3_1[415:408]} - {1'b0, layer_2_1[415:408]};
      btm_2[0] = {1'b0,layer_3_2[399:392]} - {1'b0, layer_2_2[399:392]};
      btm_2[1] = {1'b0,layer_3_2[407:400]} - {1'b0, layer_2_2[407:400]};
      btm_2[2] = {1'b0,layer_3_2[415:408]} - {1'b0, layer_2_2[415:408]};
    end
    'd51: begin
      top_0[0] = {1'b0,layer_1_0[407:400]} - {1'b0, layer_0_0[407:400]};
      top_0[1] = {1'b0,layer_1_0[415:408]} - {1'b0, layer_0_0[415:408]};
      top_0[2] = {1'b0,layer_1_0[423:416]} - {1'b0, layer_0_0[423:416]};
      top_1[0] = {1'b0,layer_1_1[407:400]} - {1'b0, layer_0_1[407:400]};
      top_1[1] = {1'b0,layer_1_1[415:408]} - {1'b0, layer_0_1[415:408]};
      top_1[2] = {1'b0,layer_1_1[423:416]} - {1'b0, layer_0_1[423:416]};
      top_2[0] = {1'b0,layer_1_2[407:400]} - {1'b0, layer_0_2[407:400]};
      top_2[1] = {1'b0,layer_1_2[415:408]} - {1'b0, layer_0_2[415:408]};
      top_2[2] = {1'b0,layer_1_2[423:416]} - {1'b0, layer_0_2[423:416]};
      mid_0[0] = {1'b0,layer_2_0[407:400]} - {1'b0, layer_1_0[407:400]};
      mid_0[1] = {1'b0,layer_2_0[415:408]} - {1'b0, layer_1_0[415:408]};
      mid_0[2] = {1'b0,layer_2_0[423:416]} - {1'b0, layer_1_0[423:416]};
      mid_1[0] = {1'b0,layer_2_1[407:400]} - {1'b0, layer_1_1[407:400]};
      mid_1[1] = {1'b0,layer_2_1[415:408]} - {1'b0, layer_1_1[415:408]};
      mid_1[2] = {1'b0,layer_2_1[423:416]} - {1'b0, layer_1_1[423:416]};
      mid_2[0] = {1'b0,layer_2_2[407:400]} - {1'b0, layer_1_2[407:400]};
      mid_2[1] = {1'b0,layer_2_2[415:408]} - {1'b0, layer_1_2[415:408]};
      mid_2[2] = {1'b0,layer_2_2[423:416]} - {1'b0, layer_1_2[423:416]};
      btm_0[0] = {1'b0,layer_3_0[407:400]} - {1'b0, layer_2_0[407:400]};
      btm_0[1] = {1'b0,layer_3_0[415:408]} - {1'b0, layer_2_0[415:408]};
      btm_0[2] = {1'b0,layer_3_0[423:416]} - {1'b0, layer_2_0[423:416]};
      btm_1[0] = {1'b0,layer_3_1[407:400]} - {1'b0, layer_2_1[407:400]};
      btm_1[1] = {1'b0,layer_3_1[415:408]} - {1'b0, layer_2_1[415:408]};
      btm_1[2] = {1'b0,layer_3_1[423:416]} - {1'b0, layer_2_1[423:416]};
      btm_2[0] = {1'b0,layer_3_2[407:400]} - {1'b0, layer_2_2[407:400]};
      btm_2[1] = {1'b0,layer_3_2[415:408]} - {1'b0, layer_2_2[415:408]};
      btm_2[2] = {1'b0,layer_3_2[423:416]} - {1'b0, layer_2_2[423:416]};
    end
    'd52: begin
      top_0[0] = {1'b0,layer_1_0[415:408]} - {1'b0, layer_0_0[415:408]};
      top_0[1] = {1'b0,layer_1_0[423:416]} - {1'b0, layer_0_0[423:416]};
      top_0[2] = {1'b0,layer_1_0[431:424]} - {1'b0, layer_0_0[431:424]};
      top_1[0] = {1'b0,layer_1_1[415:408]} - {1'b0, layer_0_1[415:408]};
      top_1[1] = {1'b0,layer_1_1[423:416]} - {1'b0, layer_0_1[423:416]};
      top_1[2] = {1'b0,layer_1_1[431:424]} - {1'b0, layer_0_1[431:424]};
      top_2[0] = {1'b0,layer_1_2[415:408]} - {1'b0, layer_0_2[415:408]};
      top_2[1] = {1'b0,layer_1_2[423:416]} - {1'b0, layer_0_2[423:416]};
      top_2[2] = {1'b0,layer_1_2[431:424]} - {1'b0, layer_0_2[431:424]};
      mid_0[0] = {1'b0,layer_2_0[415:408]} - {1'b0, layer_1_0[415:408]};
      mid_0[1] = {1'b0,layer_2_0[423:416]} - {1'b0, layer_1_0[423:416]};
      mid_0[2] = {1'b0,layer_2_0[431:424]} - {1'b0, layer_1_0[431:424]};
      mid_1[0] = {1'b0,layer_2_1[415:408]} - {1'b0, layer_1_1[415:408]};
      mid_1[1] = {1'b0,layer_2_1[423:416]} - {1'b0, layer_1_1[423:416]};
      mid_1[2] = {1'b0,layer_2_1[431:424]} - {1'b0, layer_1_1[431:424]};
      mid_2[0] = {1'b0,layer_2_2[415:408]} - {1'b0, layer_1_2[415:408]};
      mid_2[1] = {1'b0,layer_2_2[423:416]} - {1'b0, layer_1_2[423:416]};
      mid_2[2] = {1'b0,layer_2_2[431:424]} - {1'b0, layer_1_2[431:424]};
      btm_0[0] = {1'b0,layer_3_0[415:408]} - {1'b0, layer_2_0[415:408]};
      btm_0[1] = {1'b0,layer_3_0[423:416]} - {1'b0, layer_2_0[423:416]};
      btm_0[2] = {1'b0,layer_3_0[431:424]} - {1'b0, layer_2_0[431:424]};
      btm_1[0] = {1'b0,layer_3_1[415:408]} - {1'b0, layer_2_1[415:408]};
      btm_1[1] = {1'b0,layer_3_1[423:416]} - {1'b0, layer_2_1[423:416]};
      btm_1[2] = {1'b0,layer_3_1[431:424]} - {1'b0, layer_2_1[431:424]};
      btm_2[0] = {1'b0,layer_3_2[415:408]} - {1'b0, layer_2_2[415:408]};
      btm_2[1] = {1'b0,layer_3_2[423:416]} - {1'b0, layer_2_2[423:416]};
      btm_2[2] = {1'b0,layer_3_2[431:424]} - {1'b0, layer_2_2[431:424]};
    end
    'd53: begin
      top_0[0] = {1'b0,layer_1_0[423:416]} - {1'b0, layer_0_0[423:416]};
      top_0[1] = {1'b0,layer_1_0[431:424]} - {1'b0, layer_0_0[431:424]};
      top_0[2] = {1'b0,layer_1_0[439:432]} - {1'b0, layer_0_0[439:432]};
      top_1[0] = {1'b0,layer_1_1[423:416]} - {1'b0, layer_0_1[423:416]};
      top_1[1] = {1'b0,layer_1_1[431:424]} - {1'b0, layer_0_1[431:424]};
      top_1[2] = {1'b0,layer_1_1[439:432]} - {1'b0, layer_0_1[439:432]};
      top_2[0] = {1'b0,layer_1_2[423:416]} - {1'b0, layer_0_2[423:416]};
      top_2[1] = {1'b0,layer_1_2[431:424]} - {1'b0, layer_0_2[431:424]};
      top_2[2] = {1'b0,layer_1_2[439:432]} - {1'b0, layer_0_2[439:432]};
      mid_0[0] = {1'b0,layer_2_0[423:416]} - {1'b0, layer_1_0[423:416]};
      mid_0[1] = {1'b0,layer_2_0[431:424]} - {1'b0, layer_1_0[431:424]};
      mid_0[2] = {1'b0,layer_2_0[439:432]} - {1'b0, layer_1_0[439:432]};
      mid_1[0] = {1'b0,layer_2_1[423:416]} - {1'b0, layer_1_1[423:416]};
      mid_1[1] = {1'b0,layer_2_1[431:424]} - {1'b0, layer_1_1[431:424]};
      mid_1[2] = {1'b0,layer_2_1[439:432]} - {1'b0, layer_1_1[439:432]};
      mid_2[0] = {1'b0,layer_2_2[423:416]} - {1'b0, layer_1_2[423:416]};
      mid_2[1] = {1'b0,layer_2_2[431:424]} - {1'b0, layer_1_2[431:424]};
      mid_2[2] = {1'b0,layer_2_2[439:432]} - {1'b0, layer_1_2[439:432]};
      btm_0[0] = {1'b0,layer_3_0[423:416]} - {1'b0, layer_2_0[423:416]};
      btm_0[1] = {1'b0,layer_3_0[431:424]} - {1'b0, layer_2_0[431:424]};
      btm_0[2] = {1'b0,layer_3_0[439:432]} - {1'b0, layer_2_0[439:432]};
      btm_1[0] = {1'b0,layer_3_1[423:416]} - {1'b0, layer_2_1[423:416]};
      btm_1[1] = {1'b0,layer_3_1[431:424]} - {1'b0, layer_2_1[431:424]};
      btm_1[2] = {1'b0,layer_3_1[439:432]} - {1'b0, layer_2_1[439:432]};
      btm_2[0] = {1'b0,layer_3_2[423:416]} - {1'b0, layer_2_2[423:416]};
      btm_2[1] = {1'b0,layer_3_2[431:424]} - {1'b0, layer_2_2[431:424]};
      btm_2[2] = {1'b0,layer_3_2[439:432]} - {1'b0, layer_2_2[439:432]};
    end
    'd54: begin
      top_0[0] = {1'b0,layer_1_0[431:424]} - {1'b0, layer_0_0[431:424]};
      top_0[1] = {1'b0,layer_1_0[439:432]} - {1'b0, layer_0_0[439:432]};
      top_0[2] = {1'b0,layer_1_0[447:440]} - {1'b0, layer_0_0[447:440]};
      top_1[0] = {1'b0,layer_1_1[431:424]} - {1'b0, layer_0_1[431:424]};
      top_1[1] = {1'b0,layer_1_1[439:432]} - {1'b0, layer_0_1[439:432]};
      top_1[2] = {1'b0,layer_1_1[447:440]} - {1'b0, layer_0_1[447:440]};
      top_2[0] = {1'b0,layer_1_2[431:424]} - {1'b0, layer_0_2[431:424]};
      top_2[1] = {1'b0,layer_1_2[439:432]} - {1'b0, layer_0_2[439:432]};
      top_2[2] = {1'b0,layer_1_2[447:440]} - {1'b0, layer_0_2[447:440]};
      mid_0[0] = {1'b0,layer_2_0[431:424]} - {1'b0, layer_1_0[431:424]};
      mid_0[1] = {1'b0,layer_2_0[439:432]} - {1'b0, layer_1_0[439:432]};
      mid_0[2] = {1'b0,layer_2_0[447:440]} - {1'b0, layer_1_0[447:440]};
      mid_1[0] = {1'b0,layer_2_1[431:424]} - {1'b0, layer_1_1[431:424]};
      mid_1[1] = {1'b0,layer_2_1[439:432]} - {1'b0, layer_1_1[439:432]};
      mid_1[2] = {1'b0,layer_2_1[447:440]} - {1'b0, layer_1_1[447:440]};
      mid_2[0] = {1'b0,layer_2_2[431:424]} - {1'b0, layer_1_2[431:424]};
      mid_2[1] = {1'b0,layer_2_2[439:432]} - {1'b0, layer_1_2[439:432]};
      mid_2[2] = {1'b0,layer_2_2[447:440]} - {1'b0, layer_1_2[447:440]};
      btm_0[0] = {1'b0,layer_3_0[431:424]} - {1'b0, layer_2_0[431:424]};
      btm_0[1] = {1'b0,layer_3_0[439:432]} - {1'b0, layer_2_0[439:432]};
      btm_0[2] = {1'b0,layer_3_0[447:440]} - {1'b0, layer_2_0[447:440]};
      btm_1[0] = {1'b0,layer_3_1[431:424]} - {1'b0, layer_2_1[431:424]};
      btm_1[1] = {1'b0,layer_3_1[439:432]} - {1'b0, layer_2_1[439:432]};
      btm_1[2] = {1'b0,layer_3_1[447:440]} - {1'b0, layer_2_1[447:440]};
      btm_2[0] = {1'b0,layer_3_2[431:424]} - {1'b0, layer_2_2[431:424]};
      btm_2[1] = {1'b0,layer_3_2[439:432]} - {1'b0, layer_2_2[439:432]};
      btm_2[2] = {1'b0,layer_3_2[447:440]} - {1'b0, layer_2_2[447:440]};
    end
    'd55: begin
      top_0[0] = {1'b0,layer_1_0[439:432]} - {1'b0, layer_0_0[439:432]};
      top_0[1] = {1'b0,layer_1_0[447:440]} - {1'b0, layer_0_0[447:440]};
      top_0[2] = {1'b0,layer_1_0[455:448]} - {1'b0, layer_0_0[455:448]};
      top_1[0] = {1'b0,layer_1_1[439:432]} - {1'b0, layer_0_1[439:432]};
      top_1[1] = {1'b0,layer_1_1[447:440]} - {1'b0, layer_0_1[447:440]};
      top_1[2] = {1'b0,layer_1_1[455:448]} - {1'b0, layer_0_1[455:448]};
      top_2[0] = {1'b0,layer_1_2[439:432]} - {1'b0, layer_0_2[439:432]};
      top_2[1] = {1'b0,layer_1_2[447:440]} - {1'b0, layer_0_2[447:440]};
      top_2[2] = {1'b0,layer_1_2[455:448]} - {1'b0, layer_0_2[455:448]};
      mid_0[0] = {1'b0,layer_2_0[439:432]} - {1'b0, layer_1_0[439:432]};
      mid_0[1] = {1'b0,layer_2_0[447:440]} - {1'b0, layer_1_0[447:440]};
      mid_0[2] = {1'b0,layer_2_0[455:448]} - {1'b0, layer_1_0[455:448]};
      mid_1[0] = {1'b0,layer_2_1[439:432]} - {1'b0, layer_1_1[439:432]};
      mid_1[1] = {1'b0,layer_2_1[447:440]} - {1'b0, layer_1_1[447:440]};
      mid_1[2] = {1'b0,layer_2_1[455:448]} - {1'b0, layer_1_1[455:448]};
      mid_2[0] = {1'b0,layer_2_2[439:432]} - {1'b0, layer_1_2[439:432]};
      mid_2[1] = {1'b0,layer_2_2[447:440]} - {1'b0, layer_1_2[447:440]};
      mid_2[2] = {1'b0,layer_2_2[455:448]} - {1'b0, layer_1_2[455:448]};
      btm_0[0] = {1'b0,layer_3_0[439:432]} - {1'b0, layer_2_0[439:432]};
      btm_0[1] = {1'b0,layer_3_0[447:440]} - {1'b0, layer_2_0[447:440]};
      btm_0[2] = {1'b0,layer_3_0[455:448]} - {1'b0, layer_2_0[455:448]};
      btm_1[0] = {1'b0,layer_3_1[439:432]} - {1'b0, layer_2_1[439:432]};
      btm_1[1] = {1'b0,layer_3_1[447:440]} - {1'b0, layer_2_1[447:440]};
      btm_1[2] = {1'b0,layer_3_1[455:448]} - {1'b0, layer_2_1[455:448]};
      btm_2[0] = {1'b0,layer_3_2[439:432]} - {1'b0, layer_2_2[439:432]};
      btm_2[1] = {1'b0,layer_3_2[447:440]} - {1'b0, layer_2_2[447:440]};
      btm_2[2] = {1'b0,layer_3_2[455:448]} - {1'b0, layer_2_2[455:448]};
    end
    'd56: begin
      top_0[0] = {1'b0,layer_1_0[447:440]} - {1'b0, layer_0_0[447:440]};
      top_0[1] = {1'b0,layer_1_0[455:448]} - {1'b0, layer_0_0[455:448]};
      top_0[2] = {1'b0,layer_1_0[463:456]} - {1'b0, layer_0_0[463:456]};
      top_1[0] = {1'b0,layer_1_1[447:440]} - {1'b0, layer_0_1[447:440]};
      top_1[1] = {1'b0,layer_1_1[455:448]} - {1'b0, layer_0_1[455:448]};
      top_1[2] = {1'b0,layer_1_1[463:456]} - {1'b0, layer_0_1[463:456]};
      top_2[0] = {1'b0,layer_1_2[447:440]} - {1'b0, layer_0_2[447:440]};
      top_2[1] = {1'b0,layer_1_2[455:448]} - {1'b0, layer_0_2[455:448]};
      top_2[2] = {1'b0,layer_1_2[463:456]} - {1'b0, layer_0_2[463:456]};
      mid_0[0] = {1'b0,layer_2_0[447:440]} - {1'b0, layer_1_0[447:440]};
      mid_0[1] = {1'b0,layer_2_0[455:448]} - {1'b0, layer_1_0[455:448]};
      mid_0[2] = {1'b0,layer_2_0[463:456]} - {1'b0, layer_1_0[463:456]};
      mid_1[0] = {1'b0,layer_2_1[447:440]} - {1'b0, layer_1_1[447:440]};
      mid_1[1] = {1'b0,layer_2_1[455:448]} - {1'b0, layer_1_1[455:448]};
      mid_1[2] = {1'b0,layer_2_1[463:456]} - {1'b0, layer_1_1[463:456]};
      mid_2[0] = {1'b0,layer_2_2[447:440]} - {1'b0, layer_1_2[447:440]};
      mid_2[1] = {1'b0,layer_2_2[455:448]} - {1'b0, layer_1_2[455:448]};
      mid_2[2] = {1'b0,layer_2_2[463:456]} - {1'b0, layer_1_2[463:456]};
      btm_0[0] = {1'b0,layer_3_0[447:440]} - {1'b0, layer_2_0[447:440]};
      btm_0[1] = {1'b0,layer_3_0[455:448]} - {1'b0, layer_2_0[455:448]};
      btm_0[2] = {1'b0,layer_3_0[463:456]} - {1'b0, layer_2_0[463:456]};
      btm_1[0] = {1'b0,layer_3_1[447:440]} - {1'b0, layer_2_1[447:440]};
      btm_1[1] = {1'b0,layer_3_1[455:448]} - {1'b0, layer_2_1[455:448]};
      btm_1[2] = {1'b0,layer_3_1[463:456]} - {1'b0, layer_2_1[463:456]};
      btm_2[0] = {1'b0,layer_3_2[447:440]} - {1'b0, layer_2_2[447:440]};
      btm_2[1] = {1'b0,layer_3_2[455:448]} - {1'b0, layer_2_2[455:448]};
      btm_2[2] = {1'b0,layer_3_2[463:456]} - {1'b0, layer_2_2[463:456]};
    end
    'd57: begin
      top_0[0] = {1'b0,layer_1_0[455:448]} - {1'b0, layer_0_0[455:448]};
      top_0[1] = {1'b0,layer_1_0[463:456]} - {1'b0, layer_0_0[463:456]};
      top_0[2] = {1'b0,layer_1_0[471:464]} - {1'b0, layer_0_0[471:464]};
      top_1[0] = {1'b0,layer_1_1[455:448]} - {1'b0, layer_0_1[455:448]};
      top_1[1] = {1'b0,layer_1_1[463:456]} - {1'b0, layer_0_1[463:456]};
      top_1[2] = {1'b0,layer_1_1[471:464]} - {1'b0, layer_0_1[471:464]};
      top_2[0] = {1'b0,layer_1_2[455:448]} - {1'b0, layer_0_2[455:448]};
      top_2[1] = {1'b0,layer_1_2[463:456]} - {1'b0, layer_0_2[463:456]};
      top_2[2] = {1'b0,layer_1_2[471:464]} - {1'b0, layer_0_2[471:464]};
      mid_0[0] = {1'b0,layer_2_0[455:448]} - {1'b0, layer_1_0[455:448]};
      mid_0[1] = {1'b0,layer_2_0[463:456]} - {1'b0, layer_1_0[463:456]};
      mid_0[2] = {1'b0,layer_2_0[471:464]} - {1'b0, layer_1_0[471:464]};
      mid_1[0] = {1'b0,layer_2_1[455:448]} - {1'b0, layer_1_1[455:448]};
      mid_1[1] = {1'b0,layer_2_1[463:456]} - {1'b0, layer_1_1[463:456]};
      mid_1[2] = {1'b0,layer_2_1[471:464]} - {1'b0, layer_1_1[471:464]};
      mid_2[0] = {1'b0,layer_2_2[455:448]} - {1'b0, layer_1_2[455:448]};
      mid_2[1] = {1'b0,layer_2_2[463:456]} - {1'b0, layer_1_2[463:456]};
      mid_2[2] = {1'b0,layer_2_2[471:464]} - {1'b0, layer_1_2[471:464]};
      btm_0[0] = {1'b0,layer_3_0[455:448]} - {1'b0, layer_2_0[455:448]};
      btm_0[1] = {1'b0,layer_3_0[463:456]} - {1'b0, layer_2_0[463:456]};
      btm_0[2] = {1'b0,layer_3_0[471:464]} - {1'b0, layer_2_0[471:464]};
      btm_1[0] = {1'b0,layer_3_1[455:448]} - {1'b0, layer_2_1[455:448]};
      btm_1[1] = {1'b0,layer_3_1[463:456]} - {1'b0, layer_2_1[463:456]};
      btm_1[2] = {1'b0,layer_3_1[471:464]} - {1'b0, layer_2_1[471:464]};
      btm_2[0] = {1'b0,layer_3_2[455:448]} - {1'b0, layer_2_2[455:448]};
      btm_2[1] = {1'b0,layer_3_2[463:456]} - {1'b0, layer_2_2[463:456]};
      btm_2[2] = {1'b0,layer_3_2[471:464]} - {1'b0, layer_2_2[471:464]};
    end
    'd58: begin
      top_0[0] = {1'b0,layer_1_0[463:456]} - {1'b0, layer_0_0[463:456]};
      top_0[1] = {1'b0,layer_1_0[471:464]} - {1'b0, layer_0_0[471:464]};
      top_0[2] = {1'b0,layer_1_0[479:472]} - {1'b0, layer_0_0[479:472]};
      top_1[0] = {1'b0,layer_1_1[463:456]} - {1'b0, layer_0_1[463:456]};
      top_1[1] = {1'b0,layer_1_1[471:464]} - {1'b0, layer_0_1[471:464]};
      top_1[2] = {1'b0,layer_1_1[479:472]} - {1'b0, layer_0_1[479:472]};
      top_2[0] = {1'b0,layer_1_2[463:456]} - {1'b0, layer_0_2[463:456]};
      top_2[1] = {1'b0,layer_1_2[471:464]} - {1'b0, layer_0_2[471:464]};
      top_2[2] = {1'b0,layer_1_2[479:472]} - {1'b0, layer_0_2[479:472]};
      mid_0[0] = {1'b0,layer_2_0[463:456]} - {1'b0, layer_1_0[463:456]};
      mid_0[1] = {1'b0,layer_2_0[471:464]} - {1'b0, layer_1_0[471:464]};
      mid_0[2] = {1'b0,layer_2_0[479:472]} - {1'b0, layer_1_0[479:472]};
      mid_1[0] = {1'b0,layer_2_1[463:456]} - {1'b0, layer_1_1[463:456]};
      mid_1[1] = {1'b0,layer_2_1[471:464]} - {1'b0, layer_1_1[471:464]};
      mid_1[2] = {1'b0,layer_2_1[479:472]} - {1'b0, layer_1_1[479:472]};
      mid_2[0] = {1'b0,layer_2_2[463:456]} - {1'b0, layer_1_2[463:456]};
      mid_2[1] = {1'b0,layer_2_2[471:464]} - {1'b0, layer_1_2[471:464]};
      mid_2[2] = {1'b0,layer_2_2[479:472]} - {1'b0, layer_1_2[479:472]};
      btm_0[0] = {1'b0,layer_3_0[463:456]} - {1'b0, layer_2_0[463:456]};
      btm_0[1] = {1'b0,layer_3_0[471:464]} - {1'b0, layer_2_0[471:464]};
      btm_0[2] = {1'b0,layer_3_0[479:472]} - {1'b0, layer_2_0[479:472]};
      btm_1[0] = {1'b0,layer_3_1[463:456]} - {1'b0, layer_2_1[463:456]};
      btm_1[1] = {1'b0,layer_3_1[471:464]} - {1'b0, layer_2_1[471:464]};
      btm_1[2] = {1'b0,layer_3_1[479:472]} - {1'b0, layer_2_1[479:472]};
      btm_2[0] = {1'b0,layer_3_2[463:456]} - {1'b0, layer_2_2[463:456]};
      btm_2[1] = {1'b0,layer_3_2[471:464]} - {1'b0, layer_2_2[471:464]};
      btm_2[2] = {1'b0,layer_3_2[479:472]} - {1'b0, layer_2_2[479:472]};
    end
    'd59: begin
      top_0[0] = {1'b0,layer_1_0[471:464]} - {1'b0, layer_0_0[471:464]};
      top_0[1] = {1'b0,layer_1_0[479:472]} - {1'b0, layer_0_0[479:472]};
      top_0[2] = {1'b0,layer_1_0[487:480]} - {1'b0, layer_0_0[487:480]};
      top_1[0] = {1'b0,layer_1_1[471:464]} - {1'b0, layer_0_1[471:464]};
      top_1[1] = {1'b0,layer_1_1[479:472]} - {1'b0, layer_0_1[479:472]};
      top_1[2] = {1'b0,layer_1_1[487:480]} - {1'b0, layer_0_1[487:480]};
      top_2[0] = {1'b0,layer_1_2[471:464]} - {1'b0, layer_0_2[471:464]};
      top_2[1] = {1'b0,layer_1_2[479:472]} - {1'b0, layer_0_2[479:472]};
      top_2[2] = {1'b0,layer_1_2[487:480]} - {1'b0, layer_0_2[487:480]};
      mid_0[0] = {1'b0,layer_2_0[471:464]} - {1'b0, layer_1_0[471:464]};
      mid_0[1] = {1'b0,layer_2_0[479:472]} - {1'b0, layer_1_0[479:472]};
      mid_0[2] = {1'b0,layer_2_0[487:480]} - {1'b0, layer_1_0[487:480]};
      mid_1[0] = {1'b0,layer_2_1[471:464]} - {1'b0, layer_1_1[471:464]};
      mid_1[1] = {1'b0,layer_2_1[479:472]} - {1'b0, layer_1_1[479:472]};
      mid_1[2] = {1'b0,layer_2_1[487:480]} - {1'b0, layer_1_1[487:480]};
      mid_2[0] = {1'b0,layer_2_2[471:464]} - {1'b0, layer_1_2[471:464]};
      mid_2[1] = {1'b0,layer_2_2[479:472]} - {1'b0, layer_1_2[479:472]};
      mid_2[2] = {1'b0,layer_2_2[487:480]} - {1'b0, layer_1_2[487:480]};
      btm_0[0] = {1'b0,layer_3_0[471:464]} - {1'b0, layer_2_0[471:464]};
      btm_0[1] = {1'b0,layer_3_0[479:472]} - {1'b0, layer_2_0[479:472]};
      btm_0[2] = {1'b0,layer_3_0[487:480]} - {1'b0, layer_2_0[487:480]};
      btm_1[0] = {1'b0,layer_3_1[471:464]} - {1'b0, layer_2_1[471:464]};
      btm_1[1] = {1'b0,layer_3_1[479:472]} - {1'b0, layer_2_1[479:472]};
      btm_1[2] = {1'b0,layer_3_1[487:480]} - {1'b0, layer_2_1[487:480]};
      btm_2[0] = {1'b0,layer_3_2[471:464]} - {1'b0, layer_2_2[471:464]};
      btm_2[1] = {1'b0,layer_3_2[479:472]} - {1'b0, layer_2_2[479:472]};
      btm_2[2] = {1'b0,layer_3_2[487:480]} - {1'b0, layer_2_2[487:480]};
    end
    'd60: begin
      top_0[0] = {1'b0,layer_1_0[479:472]} - {1'b0, layer_0_0[479:472]};
      top_0[1] = {1'b0,layer_1_0[487:480]} - {1'b0, layer_0_0[487:480]};
      top_0[2] = {1'b0,layer_1_0[495:488]} - {1'b0, layer_0_0[495:488]};
      top_1[0] = {1'b0,layer_1_1[479:472]} - {1'b0, layer_0_1[479:472]};
      top_1[1] = {1'b0,layer_1_1[487:480]} - {1'b0, layer_0_1[487:480]};
      top_1[2] = {1'b0,layer_1_1[495:488]} - {1'b0, layer_0_1[495:488]};
      top_2[0] = {1'b0,layer_1_2[479:472]} - {1'b0, layer_0_2[479:472]};
      top_2[1] = {1'b0,layer_1_2[487:480]} - {1'b0, layer_0_2[487:480]};
      top_2[2] = {1'b0,layer_1_2[495:488]} - {1'b0, layer_0_2[495:488]};
      mid_0[0] = {1'b0,layer_2_0[479:472]} - {1'b0, layer_1_0[479:472]};
      mid_0[1] = {1'b0,layer_2_0[487:480]} - {1'b0, layer_1_0[487:480]};
      mid_0[2] = {1'b0,layer_2_0[495:488]} - {1'b0, layer_1_0[495:488]};
      mid_1[0] = {1'b0,layer_2_1[479:472]} - {1'b0, layer_1_1[479:472]};
      mid_1[1] = {1'b0,layer_2_1[487:480]} - {1'b0, layer_1_1[487:480]};
      mid_1[2] = {1'b0,layer_2_1[495:488]} - {1'b0, layer_1_1[495:488]};
      mid_2[0] = {1'b0,layer_2_2[479:472]} - {1'b0, layer_1_2[479:472]};
      mid_2[1] = {1'b0,layer_2_2[487:480]} - {1'b0, layer_1_2[487:480]};
      mid_2[2] = {1'b0,layer_2_2[495:488]} - {1'b0, layer_1_2[495:488]};
      btm_0[0] = {1'b0,layer_3_0[479:472]} - {1'b0, layer_2_0[479:472]};
      btm_0[1] = {1'b0,layer_3_0[487:480]} - {1'b0, layer_2_0[487:480]};
      btm_0[2] = {1'b0,layer_3_0[495:488]} - {1'b0, layer_2_0[495:488]};
      btm_1[0] = {1'b0,layer_3_1[479:472]} - {1'b0, layer_2_1[479:472]};
      btm_1[1] = {1'b0,layer_3_1[487:480]} - {1'b0, layer_2_1[487:480]};
      btm_1[2] = {1'b0,layer_3_1[495:488]} - {1'b0, layer_2_1[495:488]};
      btm_2[0] = {1'b0,layer_3_2[479:472]} - {1'b0, layer_2_2[479:472]};
      btm_2[1] = {1'b0,layer_3_2[487:480]} - {1'b0, layer_2_2[487:480]};
      btm_2[2] = {1'b0,layer_3_2[495:488]} - {1'b0, layer_2_2[495:488]};
    end
    'd61: begin
      top_0[0] = {1'b0,layer_1_0[487:480]} - {1'b0, layer_0_0[487:480]};
      top_0[1] = {1'b0,layer_1_0[495:488]} - {1'b0, layer_0_0[495:488]};
      top_0[2] = {1'b0,layer_1_0[503:496]} - {1'b0, layer_0_0[503:496]};
      top_1[0] = {1'b0,layer_1_1[487:480]} - {1'b0, layer_0_1[487:480]};
      top_1[1] = {1'b0,layer_1_1[495:488]} - {1'b0, layer_0_1[495:488]};
      top_1[2] = {1'b0,layer_1_1[503:496]} - {1'b0, layer_0_1[503:496]};
      top_2[0] = {1'b0,layer_1_2[487:480]} - {1'b0, layer_0_2[487:480]};
      top_2[1] = {1'b0,layer_1_2[495:488]} - {1'b0, layer_0_2[495:488]};
      top_2[2] = {1'b0,layer_1_2[503:496]} - {1'b0, layer_0_2[503:496]};
      mid_0[0] = {1'b0,layer_2_0[487:480]} - {1'b0, layer_1_0[487:480]};
      mid_0[1] = {1'b0,layer_2_0[495:488]} - {1'b0, layer_1_0[495:488]};
      mid_0[2] = {1'b0,layer_2_0[503:496]} - {1'b0, layer_1_0[503:496]};
      mid_1[0] = {1'b0,layer_2_1[487:480]} - {1'b0, layer_1_1[487:480]};
      mid_1[1] = {1'b0,layer_2_1[495:488]} - {1'b0, layer_1_1[495:488]};
      mid_1[2] = {1'b0,layer_2_1[503:496]} - {1'b0, layer_1_1[503:496]};
      mid_2[0] = {1'b0,layer_2_2[487:480]} - {1'b0, layer_1_2[487:480]};
      mid_2[1] = {1'b0,layer_2_2[495:488]} - {1'b0, layer_1_2[495:488]};
      mid_2[2] = {1'b0,layer_2_2[503:496]} - {1'b0, layer_1_2[503:496]};
      btm_0[0] = {1'b0,layer_3_0[487:480]} - {1'b0, layer_2_0[487:480]};
      btm_0[1] = {1'b0,layer_3_0[495:488]} - {1'b0, layer_2_0[495:488]};
      btm_0[2] = {1'b0,layer_3_0[503:496]} - {1'b0, layer_2_0[503:496]};
      btm_1[0] = {1'b0,layer_3_1[487:480]} - {1'b0, layer_2_1[487:480]};
      btm_1[1] = {1'b0,layer_3_1[495:488]} - {1'b0, layer_2_1[495:488]};
      btm_1[2] = {1'b0,layer_3_1[503:496]} - {1'b0, layer_2_1[503:496]};
      btm_2[0] = {1'b0,layer_3_2[487:480]} - {1'b0, layer_2_2[487:480]};
      btm_2[1] = {1'b0,layer_3_2[495:488]} - {1'b0, layer_2_2[495:488]};
      btm_2[2] = {1'b0,layer_3_2[503:496]} - {1'b0, layer_2_2[503:496]};
    end
    'd62: begin
      top_0[0] = {1'b0,layer_1_0[495:488]} - {1'b0, layer_0_0[495:488]};
      top_0[1] = {1'b0,layer_1_0[503:496]} - {1'b0, layer_0_0[503:496]};
      top_0[2] = {1'b0,layer_1_0[511:504]} - {1'b0, layer_0_0[511:504]};
      top_1[0] = {1'b0,layer_1_1[495:488]} - {1'b0, layer_0_1[495:488]};
      top_1[1] = {1'b0,layer_1_1[503:496]} - {1'b0, layer_0_1[503:496]};
      top_1[2] = {1'b0,layer_1_1[511:504]} - {1'b0, layer_0_1[511:504]};
      top_2[0] = {1'b0,layer_1_2[495:488]} - {1'b0, layer_0_2[495:488]};
      top_2[1] = {1'b0,layer_1_2[503:496]} - {1'b0, layer_0_2[503:496]};
      top_2[2] = {1'b0,layer_1_2[511:504]} - {1'b0, layer_0_2[511:504]};
      mid_0[0] = {1'b0,layer_2_0[495:488]} - {1'b0, layer_1_0[495:488]};
      mid_0[1] = {1'b0,layer_2_0[503:496]} - {1'b0, layer_1_0[503:496]};
      mid_0[2] = {1'b0,layer_2_0[511:504]} - {1'b0, layer_1_0[511:504]};
      mid_1[0] = {1'b0,layer_2_1[495:488]} - {1'b0, layer_1_1[495:488]};
      mid_1[1] = {1'b0,layer_2_1[503:496]} - {1'b0, layer_1_1[503:496]};
      mid_1[2] = {1'b0,layer_2_1[511:504]} - {1'b0, layer_1_1[511:504]};
      mid_2[0] = {1'b0,layer_2_2[495:488]} - {1'b0, layer_1_2[495:488]};
      mid_2[1] = {1'b0,layer_2_2[503:496]} - {1'b0, layer_1_2[503:496]};
      mid_2[2] = {1'b0,layer_2_2[511:504]} - {1'b0, layer_1_2[511:504]};
      btm_0[0] = {1'b0,layer_3_0[495:488]} - {1'b0, layer_2_0[495:488]};
      btm_0[1] = {1'b0,layer_3_0[503:496]} - {1'b0, layer_2_0[503:496]};
      btm_0[2] = {1'b0,layer_3_0[511:504]} - {1'b0, layer_2_0[511:504]};
      btm_1[0] = {1'b0,layer_3_1[495:488]} - {1'b0, layer_2_1[495:488]};
      btm_1[1] = {1'b0,layer_3_1[503:496]} - {1'b0, layer_2_1[503:496]};
      btm_1[2] = {1'b0,layer_3_1[511:504]} - {1'b0, layer_2_1[511:504]};
      btm_2[0] = {1'b0,layer_3_2[495:488]} - {1'b0, layer_2_2[495:488]};
      btm_2[1] = {1'b0,layer_3_2[503:496]} - {1'b0, layer_2_2[503:496]};
      btm_2[2] = {1'b0,layer_3_2[511:504]} - {1'b0, layer_2_2[511:504]};
    end
    'd63: begin
      top_0[0] = {1'b0,layer_1_0[503:496]} - {1'b0, layer_0_0[503:496]};
      top_0[1] = {1'b0,layer_1_0[511:504]} - {1'b0, layer_0_0[511:504]};
      top_0[2] = {1'b0,layer_1_0[519:512]} - {1'b0, layer_0_0[519:512]};
      top_1[0] = {1'b0,layer_1_1[503:496]} - {1'b0, layer_0_1[503:496]};
      top_1[1] = {1'b0,layer_1_1[511:504]} - {1'b0, layer_0_1[511:504]};
      top_1[2] = {1'b0,layer_1_1[519:512]} - {1'b0, layer_0_1[519:512]};
      top_2[0] = {1'b0,layer_1_2[503:496]} - {1'b0, layer_0_2[503:496]};
      top_2[1] = {1'b0,layer_1_2[511:504]} - {1'b0, layer_0_2[511:504]};
      top_2[2] = {1'b0,layer_1_2[519:512]} - {1'b0, layer_0_2[519:512]};
      mid_0[0] = {1'b0,layer_2_0[503:496]} - {1'b0, layer_1_0[503:496]};
      mid_0[1] = {1'b0,layer_2_0[511:504]} - {1'b0, layer_1_0[511:504]};
      mid_0[2] = {1'b0,layer_2_0[519:512]} - {1'b0, layer_1_0[519:512]};
      mid_1[0] = {1'b0,layer_2_1[503:496]} - {1'b0, layer_1_1[503:496]};
      mid_1[1] = {1'b0,layer_2_1[511:504]} - {1'b0, layer_1_1[511:504]};
      mid_1[2] = {1'b0,layer_2_1[519:512]} - {1'b0, layer_1_1[519:512]};
      mid_2[0] = {1'b0,layer_2_2[503:496]} - {1'b0, layer_1_2[503:496]};
      mid_2[1] = {1'b0,layer_2_2[511:504]} - {1'b0, layer_1_2[511:504]};
      mid_2[2] = {1'b0,layer_2_2[519:512]} - {1'b0, layer_1_2[519:512]};
      btm_0[0] = {1'b0,layer_3_0[503:496]} - {1'b0, layer_2_0[503:496]};
      btm_0[1] = {1'b0,layer_3_0[511:504]} - {1'b0, layer_2_0[511:504]};
      btm_0[2] = {1'b0,layer_3_0[519:512]} - {1'b0, layer_2_0[519:512]};
      btm_1[0] = {1'b0,layer_3_1[503:496]} - {1'b0, layer_2_1[503:496]};
      btm_1[1] = {1'b0,layer_3_1[511:504]} - {1'b0, layer_2_1[511:504]};
      btm_1[2] = {1'b0,layer_3_1[519:512]} - {1'b0, layer_2_1[519:512]};
      btm_2[0] = {1'b0,layer_3_2[503:496]} - {1'b0, layer_2_2[503:496]};
      btm_2[1] = {1'b0,layer_3_2[511:504]} - {1'b0, layer_2_2[511:504]};
      btm_2[2] = {1'b0,layer_3_2[519:512]} - {1'b0, layer_2_2[519:512]};
    end
    'd64: begin
      top_0[0] = {1'b0,layer_1_0[511:504]} - {1'b0, layer_0_0[511:504]};
      top_0[1] = {1'b0,layer_1_0[519:512]} - {1'b0, layer_0_0[519:512]};
      top_0[2] = {1'b0,layer_1_0[527:520]} - {1'b0, layer_0_0[527:520]};
      top_1[0] = {1'b0,layer_1_1[511:504]} - {1'b0, layer_0_1[511:504]};
      top_1[1] = {1'b0,layer_1_1[519:512]} - {1'b0, layer_0_1[519:512]};
      top_1[2] = {1'b0,layer_1_1[527:520]} - {1'b0, layer_0_1[527:520]};
      top_2[0] = {1'b0,layer_1_2[511:504]} - {1'b0, layer_0_2[511:504]};
      top_2[1] = {1'b0,layer_1_2[519:512]} - {1'b0, layer_0_2[519:512]};
      top_2[2] = {1'b0,layer_1_2[527:520]} - {1'b0, layer_0_2[527:520]};
      mid_0[0] = {1'b0,layer_2_0[511:504]} - {1'b0, layer_1_0[511:504]};
      mid_0[1] = {1'b0,layer_2_0[519:512]} - {1'b0, layer_1_0[519:512]};
      mid_0[2] = {1'b0,layer_2_0[527:520]} - {1'b0, layer_1_0[527:520]};
      mid_1[0] = {1'b0,layer_2_1[511:504]} - {1'b0, layer_1_1[511:504]};
      mid_1[1] = {1'b0,layer_2_1[519:512]} - {1'b0, layer_1_1[519:512]};
      mid_1[2] = {1'b0,layer_2_1[527:520]} - {1'b0, layer_1_1[527:520]};
      mid_2[0] = {1'b0,layer_2_2[511:504]} - {1'b0, layer_1_2[511:504]};
      mid_2[1] = {1'b0,layer_2_2[519:512]} - {1'b0, layer_1_2[519:512]};
      mid_2[2] = {1'b0,layer_2_2[527:520]} - {1'b0, layer_1_2[527:520]};
      btm_0[0] = {1'b0,layer_3_0[511:504]} - {1'b0, layer_2_0[511:504]};
      btm_0[1] = {1'b0,layer_3_0[519:512]} - {1'b0, layer_2_0[519:512]};
      btm_0[2] = {1'b0,layer_3_0[527:520]} - {1'b0, layer_2_0[527:520]};
      btm_1[0] = {1'b0,layer_3_1[511:504]} - {1'b0, layer_2_1[511:504]};
      btm_1[1] = {1'b0,layer_3_1[519:512]} - {1'b0, layer_2_1[519:512]};
      btm_1[2] = {1'b0,layer_3_1[527:520]} - {1'b0, layer_2_1[527:520]};
      btm_2[0] = {1'b0,layer_3_2[511:504]} - {1'b0, layer_2_2[511:504]};
      btm_2[1] = {1'b0,layer_3_2[519:512]} - {1'b0, layer_2_2[519:512]};
      btm_2[2] = {1'b0,layer_3_2[527:520]} - {1'b0, layer_2_2[527:520]};
    end
    'd65: begin
      top_0[0] = {1'b0,layer_1_0[519:512]} - {1'b0, layer_0_0[519:512]};
      top_0[1] = {1'b0,layer_1_0[527:520]} - {1'b0, layer_0_0[527:520]};
      top_0[2] = {1'b0,layer_1_0[535:528]} - {1'b0, layer_0_0[535:528]};
      top_1[0] = {1'b0,layer_1_1[519:512]} - {1'b0, layer_0_1[519:512]};
      top_1[1] = {1'b0,layer_1_1[527:520]} - {1'b0, layer_0_1[527:520]};
      top_1[2] = {1'b0,layer_1_1[535:528]} - {1'b0, layer_0_1[535:528]};
      top_2[0] = {1'b0,layer_1_2[519:512]} - {1'b0, layer_0_2[519:512]};
      top_2[1] = {1'b0,layer_1_2[527:520]} - {1'b0, layer_0_2[527:520]};
      top_2[2] = {1'b0,layer_1_2[535:528]} - {1'b0, layer_0_2[535:528]};
      mid_0[0] = {1'b0,layer_2_0[519:512]} - {1'b0, layer_1_0[519:512]};
      mid_0[1] = {1'b0,layer_2_0[527:520]} - {1'b0, layer_1_0[527:520]};
      mid_0[2] = {1'b0,layer_2_0[535:528]} - {1'b0, layer_1_0[535:528]};
      mid_1[0] = {1'b0,layer_2_1[519:512]} - {1'b0, layer_1_1[519:512]};
      mid_1[1] = {1'b0,layer_2_1[527:520]} - {1'b0, layer_1_1[527:520]};
      mid_1[2] = {1'b0,layer_2_1[535:528]} - {1'b0, layer_1_1[535:528]};
      mid_2[0] = {1'b0,layer_2_2[519:512]} - {1'b0, layer_1_2[519:512]};
      mid_2[1] = {1'b0,layer_2_2[527:520]} - {1'b0, layer_1_2[527:520]};
      mid_2[2] = {1'b0,layer_2_2[535:528]} - {1'b0, layer_1_2[535:528]};
      btm_0[0] = {1'b0,layer_3_0[519:512]} - {1'b0, layer_2_0[519:512]};
      btm_0[1] = {1'b0,layer_3_0[527:520]} - {1'b0, layer_2_0[527:520]};
      btm_0[2] = {1'b0,layer_3_0[535:528]} - {1'b0, layer_2_0[535:528]};
      btm_1[0] = {1'b0,layer_3_1[519:512]} - {1'b0, layer_2_1[519:512]};
      btm_1[1] = {1'b0,layer_3_1[527:520]} - {1'b0, layer_2_1[527:520]};
      btm_1[2] = {1'b0,layer_3_1[535:528]} - {1'b0, layer_2_1[535:528]};
      btm_2[0] = {1'b0,layer_3_2[519:512]} - {1'b0, layer_2_2[519:512]};
      btm_2[1] = {1'b0,layer_3_2[527:520]} - {1'b0, layer_2_2[527:520]};
      btm_2[2] = {1'b0,layer_3_2[535:528]} - {1'b0, layer_2_2[535:528]};
    end
    'd66: begin
      top_0[0] = {1'b0,layer_1_0[527:520]} - {1'b0, layer_0_0[527:520]};
      top_0[1] = {1'b0,layer_1_0[535:528]} - {1'b0, layer_0_0[535:528]};
      top_0[2] = {1'b0,layer_1_0[543:536]} - {1'b0, layer_0_0[543:536]};
      top_1[0] = {1'b0,layer_1_1[527:520]} - {1'b0, layer_0_1[527:520]};
      top_1[1] = {1'b0,layer_1_1[535:528]} - {1'b0, layer_0_1[535:528]};
      top_1[2] = {1'b0,layer_1_1[543:536]} - {1'b0, layer_0_1[543:536]};
      top_2[0] = {1'b0,layer_1_2[527:520]} - {1'b0, layer_0_2[527:520]};
      top_2[1] = {1'b0,layer_1_2[535:528]} - {1'b0, layer_0_2[535:528]};
      top_2[2] = {1'b0,layer_1_2[543:536]} - {1'b0, layer_0_2[543:536]};
      mid_0[0] = {1'b0,layer_2_0[527:520]} - {1'b0, layer_1_0[527:520]};
      mid_0[1] = {1'b0,layer_2_0[535:528]} - {1'b0, layer_1_0[535:528]};
      mid_0[2] = {1'b0,layer_2_0[543:536]} - {1'b0, layer_1_0[543:536]};
      mid_1[0] = {1'b0,layer_2_1[527:520]} - {1'b0, layer_1_1[527:520]};
      mid_1[1] = {1'b0,layer_2_1[535:528]} - {1'b0, layer_1_1[535:528]};
      mid_1[2] = {1'b0,layer_2_1[543:536]} - {1'b0, layer_1_1[543:536]};
      mid_2[0] = {1'b0,layer_2_2[527:520]} - {1'b0, layer_1_2[527:520]};
      mid_2[1] = {1'b0,layer_2_2[535:528]} - {1'b0, layer_1_2[535:528]};
      mid_2[2] = {1'b0,layer_2_2[543:536]} - {1'b0, layer_1_2[543:536]};
      btm_0[0] = {1'b0,layer_3_0[527:520]} - {1'b0, layer_2_0[527:520]};
      btm_0[1] = {1'b0,layer_3_0[535:528]} - {1'b0, layer_2_0[535:528]};
      btm_0[2] = {1'b0,layer_3_0[543:536]} - {1'b0, layer_2_0[543:536]};
      btm_1[0] = {1'b0,layer_3_1[527:520]} - {1'b0, layer_2_1[527:520]};
      btm_1[1] = {1'b0,layer_3_1[535:528]} - {1'b0, layer_2_1[535:528]};
      btm_1[2] = {1'b0,layer_3_1[543:536]} - {1'b0, layer_2_1[543:536]};
      btm_2[0] = {1'b0,layer_3_2[527:520]} - {1'b0, layer_2_2[527:520]};
      btm_2[1] = {1'b0,layer_3_2[535:528]} - {1'b0, layer_2_2[535:528]};
      btm_2[2] = {1'b0,layer_3_2[543:536]} - {1'b0, layer_2_2[543:536]};
    end
    'd67: begin
      top_0[0] = {1'b0,layer_1_0[535:528]} - {1'b0, layer_0_0[535:528]};
      top_0[1] = {1'b0,layer_1_0[543:536]} - {1'b0, layer_0_0[543:536]};
      top_0[2] = {1'b0,layer_1_0[551:544]} - {1'b0, layer_0_0[551:544]};
      top_1[0] = {1'b0,layer_1_1[535:528]} - {1'b0, layer_0_1[535:528]};
      top_1[1] = {1'b0,layer_1_1[543:536]} - {1'b0, layer_0_1[543:536]};
      top_1[2] = {1'b0,layer_1_1[551:544]} - {1'b0, layer_0_1[551:544]};
      top_2[0] = {1'b0,layer_1_2[535:528]} - {1'b0, layer_0_2[535:528]};
      top_2[1] = {1'b0,layer_1_2[543:536]} - {1'b0, layer_0_2[543:536]};
      top_2[2] = {1'b0,layer_1_2[551:544]} - {1'b0, layer_0_2[551:544]};
      mid_0[0] = {1'b0,layer_2_0[535:528]} - {1'b0, layer_1_0[535:528]};
      mid_0[1] = {1'b0,layer_2_0[543:536]} - {1'b0, layer_1_0[543:536]};
      mid_0[2] = {1'b0,layer_2_0[551:544]} - {1'b0, layer_1_0[551:544]};
      mid_1[0] = {1'b0,layer_2_1[535:528]} - {1'b0, layer_1_1[535:528]};
      mid_1[1] = {1'b0,layer_2_1[543:536]} - {1'b0, layer_1_1[543:536]};
      mid_1[2] = {1'b0,layer_2_1[551:544]} - {1'b0, layer_1_1[551:544]};
      mid_2[0] = {1'b0,layer_2_2[535:528]} - {1'b0, layer_1_2[535:528]};
      mid_2[1] = {1'b0,layer_2_2[543:536]} - {1'b0, layer_1_2[543:536]};
      mid_2[2] = {1'b0,layer_2_2[551:544]} - {1'b0, layer_1_2[551:544]};
      btm_0[0] = {1'b0,layer_3_0[535:528]} - {1'b0, layer_2_0[535:528]};
      btm_0[1] = {1'b0,layer_3_0[543:536]} - {1'b0, layer_2_0[543:536]};
      btm_0[2] = {1'b0,layer_3_0[551:544]} - {1'b0, layer_2_0[551:544]};
      btm_1[0] = {1'b0,layer_3_1[535:528]} - {1'b0, layer_2_1[535:528]};
      btm_1[1] = {1'b0,layer_3_1[543:536]} - {1'b0, layer_2_1[543:536]};
      btm_1[2] = {1'b0,layer_3_1[551:544]} - {1'b0, layer_2_1[551:544]};
      btm_2[0] = {1'b0,layer_3_2[535:528]} - {1'b0, layer_2_2[535:528]};
      btm_2[1] = {1'b0,layer_3_2[543:536]} - {1'b0, layer_2_2[543:536]};
      btm_2[2] = {1'b0,layer_3_2[551:544]} - {1'b0, layer_2_2[551:544]};
    end
    'd68: begin
      top_0[0] = {1'b0,layer_1_0[543:536]} - {1'b0, layer_0_0[543:536]};
      top_0[1] = {1'b0,layer_1_0[551:544]} - {1'b0, layer_0_0[551:544]};
      top_0[2] = {1'b0,layer_1_0[559:552]} - {1'b0, layer_0_0[559:552]};
      top_1[0] = {1'b0,layer_1_1[543:536]} - {1'b0, layer_0_1[543:536]};
      top_1[1] = {1'b0,layer_1_1[551:544]} - {1'b0, layer_0_1[551:544]};
      top_1[2] = {1'b0,layer_1_1[559:552]} - {1'b0, layer_0_1[559:552]};
      top_2[0] = {1'b0,layer_1_2[543:536]} - {1'b0, layer_0_2[543:536]};
      top_2[1] = {1'b0,layer_1_2[551:544]} - {1'b0, layer_0_2[551:544]};
      top_2[2] = {1'b0,layer_1_2[559:552]} - {1'b0, layer_0_2[559:552]};
      mid_0[0] = {1'b0,layer_2_0[543:536]} - {1'b0, layer_1_0[543:536]};
      mid_0[1] = {1'b0,layer_2_0[551:544]} - {1'b0, layer_1_0[551:544]};
      mid_0[2] = {1'b0,layer_2_0[559:552]} - {1'b0, layer_1_0[559:552]};
      mid_1[0] = {1'b0,layer_2_1[543:536]} - {1'b0, layer_1_1[543:536]};
      mid_1[1] = {1'b0,layer_2_1[551:544]} - {1'b0, layer_1_1[551:544]};
      mid_1[2] = {1'b0,layer_2_1[559:552]} - {1'b0, layer_1_1[559:552]};
      mid_2[0] = {1'b0,layer_2_2[543:536]} - {1'b0, layer_1_2[543:536]};
      mid_2[1] = {1'b0,layer_2_2[551:544]} - {1'b0, layer_1_2[551:544]};
      mid_2[2] = {1'b0,layer_2_2[559:552]} - {1'b0, layer_1_2[559:552]};
      btm_0[0] = {1'b0,layer_3_0[543:536]} - {1'b0, layer_2_0[543:536]};
      btm_0[1] = {1'b0,layer_3_0[551:544]} - {1'b0, layer_2_0[551:544]};
      btm_0[2] = {1'b0,layer_3_0[559:552]} - {1'b0, layer_2_0[559:552]};
      btm_1[0] = {1'b0,layer_3_1[543:536]} - {1'b0, layer_2_1[543:536]};
      btm_1[1] = {1'b0,layer_3_1[551:544]} - {1'b0, layer_2_1[551:544]};
      btm_1[2] = {1'b0,layer_3_1[559:552]} - {1'b0, layer_2_1[559:552]};
      btm_2[0] = {1'b0,layer_3_2[543:536]} - {1'b0, layer_2_2[543:536]};
      btm_2[1] = {1'b0,layer_3_2[551:544]} - {1'b0, layer_2_2[551:544]};
      btm_2[2] = {1'b0,layer_3_2[559:552]} - {1'b0, layer_2_2[559:552]};
    end
    'd69: begin
      top_0[0] = {1'b0,layer_1_0[551:544]} - {1'b0, layer_0_0[551:544]};
      top_0[1] = {1'b0,layer_1_0[559:552]} - {1'b0, layer_0_0[559:552]};
      top_0[2] = {1'b0,layer_1_0[567:560]} - {1'b0, layer_0_0[567:560]};
      top_1[0] = {1'b0,layer_1_1[551:544]} - {1'b0, layer_0_1[551:544]};
      top_1[1] = {1'b0,layer_1_1[559:552]} - {1'b0, layer_0_1[559:552]};
      top_1[2] = {1'b0,layer_1_1[567:560]} - {1'b0, layer_0_1[567:560]};
      top_2[0] = {1'b0,layer_1_2[551:544]} - {1'b0, layer_0_2[551:544]};
      top_2[1] = {1'b0,layer_1_2[559:552]} - {1'b0, layer_0_2[559:552]};
      top_2[2] = {1'b0,layer_1_2[567:560]} - {1'b0, layer_0_2[567:560]};
      mid_0[0] = {1'b0,layer_2_0[551:544]} - {1'b0, layer_1_0[551:544]};
      mid_0[1] = {1'b0,layer_2_0[559:552]} - {1'b0, layer_1_0[559:552]};
      mid_0[2] = {1'b0,layer_2_0[567:560]} - {1'b0, layer_1_0[567:560]};
      mid_1[0] = {1'b0,layer_2_1[551:544]} - {1'b0, layer_1_1[551:544]};
      mid_1[1] = {1'b0,layer_2_1[559:552]} - {1'b0, layer_1_1[559:552]};
      mid_1[2] = {1'b0,layer_2_1[567:560]} - {1'b0, layer_1_1[567:560]};
      mid_2[0] = {1'b0,layer_2_2[551:544]} - {1'b0, layer_1_2[551:544]};
      mid_2[1] = {1'b0,layer_2_2[559:552]} - {1'b0, layer_1_2[559:552]};
      mid_2[2] = {1'b0,layer_2_2[567:560]} - {1'b0, layer_1_2[567:560]};
      btm_0[0] = {1'b0,layer_3_0[551:544]} - {1'b0, layer_2_0[551:544]};
      btm_0[1] = {1'b0,layer_3_0[559:552]} - {1'b0, layer_2_0[559:552]};
      btm_0[2] = {1'b0,layer_3_0[567:560]} - {1'b0, layer_2_0[567:560]};
      btm_1[0] = {1'b0,layer_3_1[551:544]} - {1'b0, layer_2_1[551:544]};
      btm_1[1] = {1'b0,layer_3_1[559:552]} - {1'b0, layer_2_1[559:552]};
      btm_1[2] = {1'b0,layer_3_1[567:560]} - {1'b0, layer_2_1[567:560]};
      btm_2[0] = {1'b0,layer_3_2[551:544]} - {1'b0, layer_2_2[551:544]};
      btm_2[1] = {1'b0,layer_3_2[559:552]} - {1'b0, layer_2_2[559:552]};
      btm_2[2] = {1'b0,layer_3_2[567:560]} - {1'b0, layer_2_2[567:560]};
    end
    'd70: begin
      top_0[0] = {1'b0,layer_1_0[559:552]} - {1'b0, layer_0_0[559:552]};
      top_0[1] = {1'b0,layer_1_0[567:560]} - {1'b0, layer_0_0[567:560]};
      top_0[2] = {1'b0,layer_1_0[575:568]} - {1'b0, layer_0_0[575:568]};
      top_1[0] = {1'b0,layer_1_1[559:552]} - {1'b0, layer_0_1[559:552]};
      top_1[1] = {1'b0,layer_1_1[567:560]} - {1'b0, layer_0_1[567:560]};
      top_1[2] = {1'b0,layer_1_1[575:568]} - {1'b0, layer_0_1[575:568]};
      top_2[0] = {1'b0,layer_1_2[559:552]} - {1'b0, layer_0_2[559:552]};
      top_2[1] = {1'b0,layer_1_2[567:560]} - {1'b0, layer_0_2[567:560]};
      top_2[2] = {1'b0,layer_1_2[575:568]} - {1'b0, layer_0_2[575:568]};
      mid_0[0] = {1'b0,layer_2_0[559:552]} - {1'b0, layer_1_0[559:552]};
      mid_0[1] = {1'b0,layer_2_0[567:560]} - {1'b0, layer_1_0[567:560]};
      mid_0[2] = {1'b0,layer_2_0[575:568]} - {1'b0, layer_1_0[575:568]};
      mid_1[0] = {1'b0,layer_2_1[559:552]} - {1'b0, layer_1_1[559:552]};
      mid_1[1] = {1'b0,layer_2_1[567:560]} - {1'b0, layer_1_1[567:560]};
      mid_1[2] = {1'b0,layer_2_1[575:568]} - {1'b0, layer_1_1[575:568]};
      mid_2[0] = {1'b0,layer_2_2[559:552]} - {1'b0, layer_1_2[559:552]};
      mid_2[1] = {1'b0,layer_2_2[567:560]} - {1'b0, layer_1_2[567:560]};
      mid_2[2] = {1'b0,layer_2_2[575:568]} - {1'b0, layer_1_2[575:568]};
      btm_0[0] = {1'b0,layer_3_0[559:552]} - {1'b0, layer_2_0[559:552]};
      btm_0[1] = {1'b0,layer_3_0[567:560]} - {1'b0, layer_2_0[567:560]};
      btm_0[2] = {1'b0,layer_3_0[575:568]} - {1'b0, layer_2_0[575:568]};
      btm_1[0] = {1'b0,layer_3_1[559:552]} - {1'b0, layer_2_1[559:552]};
      btm_1[1] = {1'b0,layer_3_1[567:560]} - {1'b0, layer_2_1[567:560]};
      btm_1[2] = {1'b0,layer_3_1[575:568]} - {1'b0, layer_2_1[575:568]};
      btm_2[0] = {1'b0,layer_3_2[559:552]} - {1'b0, layer_2_2[559:552]};
      btm_2[1] = {1'b0,layer_3_2[567:560]} - {1'b0, layer_2_2[567:560]};
      btm_2[2] = {1'b0,layer_3_2[575:568]} - {1'b0, layer_2_2[575:568]};
    end
    'd71: begin
      top_0[0] = {1'b0,layer_1_0[567:560]} - {1'b0, layer_0_0[567:560]};
      top_0[1] = {1'b0,layer_1_0[575:568]} - {1'b0, layer_0_0[575:568]};
      top_0[2] = {1'b0,layer_1_0[583:576]} - {1'b0, layer_0_0[583:576]};
      top_1[0] = {1'b0,layer_1_1[567:560]} - {1'b0, layer_0_1[567:560]};
      top_1[1] = {1'b0,layer_1_1[575:568]} - {1'b0, layer_0_1[575:568]};
      top_1[2] = {1'b0,layer_1_1[583:576]} - {1'b0, layer_0_1[583:576]};
      top_2[0] = {1'b0,layer_1_2[567:560]} - {1'b0, layer_0_2[567:560]};
      top_2[1] = {1'b0,layer_1_2[575:568]} - {1'b0, layer_0_2[575:568]};
      top_2[2] = {1'b0,layer_1_2[583:576]} - {1'b0, layer_0_2[583:576]};
      mid_0[0] = {1'b0,layer_2_0[567:560]} - {1'b0, layer_1_0[567:560]};
      mid_0[1] = {1'b0,layer_2_0[575:568]} - {1'b0, layer_1_0[575:568]};
      mid_0[2] = {1'b0,layer_2_0[583:576]} - {1'b0, layer_1_0[583:576]};
      mid_1[0] = {1'b0,layer_2_1[567:560]} - {1'b0, layer_1_1[567:560]};
      mid_1[1] = {1'b0,layer_2_1[575:568]} - {1'b0, layer_1_1[575:568]};
      mid_1[2] = {1'b0,layer_2_1[583:576]} - {1'b0, layer_1_1[583:576]};
      mid_2[0] = {1'b0,layer_2_2[567:560]} - {1'b0, layer_1_2[567:560]};
      mid_2[1] = {1'b0,layer_2_2[575:568]} - {1'b0, layer_1_2[575:568]};
      mid_2[2] = {1'b0,layer_2_2[583:576]} - {1'b0, layer_1_2[583:576]};
      btm_0[0] = {1'b0,layer_3_0[567:560]} - {1'b0, layer_2_0[567:560]};
      btm_0[1] = {1'b0,layer_3_0[575:568]} - {1'b0, layer_2_0[575:568]};
      btm_0[2] = {1'b0,layer_3_0[583:576]} - {1'b0, layer_2_0[583:576]};
      btm_1[0] = {1'b0,layer_3_1[567:560]} - {1'b0, layer_2_1[567:560]};
      btm_1[1] = {1'b0,layer_3_1[575:568]} - {1'b0, layer_2_1[575:568]};
      btm_1[2] = {1'b0,layer_3_1[583:576]} - {1'b0, layer_2_1[583:576]};
      btm_2[0] = {1'b0,layer_3_2[567:560]} - {1'b0, layer_2_2[567:560]};
      btm_2[1] = {1'b0,layer_3_2[575:568]} - {1'b0, layer_2_2[575:568]};
      btm_2[2] = {1'b0,layer_3_2[583:576]} - {1'b0, layer_2_2[583:576]};
    end
    'd72: begin
      top_0[0] = {1'b0,layer_1_0[575:568]} - {1'b0, layer_0_0[575:568]};
      top_0[1] = {1'b0,layer_1_0[583:576]} - {1'b0, layer_0_0[583:576]};
      top_0[2] = {1'b0,layer_1_0[591:584]} - {1'b0, layer_0_0[591:584]};
      top_1[0] = {1'b0,layer_1_1[575:568]} - {1'b0, layer_0_1[575:568]};
      top_1[1] = {1'b0,layer_1_1[583:576]} - {1'b0, layer_0_1[583:576]};
      top_1[2] = {1'b0,layer_1_1[591:584]} - {1'b0, layer_0_1[591:584]};
      top_2[0] = {1'b0,layer_1_2[575:568]} - {1'b0, layer_0_2[575:568]};
      top_2[1] = {1'b0,layer_1_2[583:576]} - {1'b0, layer_0_2[583:576]};
      top_2[2] = {1'b0,layer_1_2[591:584]} - {1'b0, layer_0_2[591:584]};
      mid_0[0] = {1'b0,layer_2_0[575:568]} - {1'b0, layer_1_0[575:568]};
      mid_0[1] = {1'b0,layer_2_0[583:576]} - {1'b0, layer_1_0[583:576]};
      mid_0[2] = {1'b0,layer_2_0[591:584]} - {1'b0, layer_1_0[591:584]};
      mid_1[0] = {1'b0,layer_2_1[575:568]} - {1'b0, layer_1_1[575:568]};
      mid_1[1] = {1'b0,layer_2_1[583:576]} - {1'b0, layer_1_1[583:576]};
      mid_1[2] = {1'b0,layer_2_1[591:584]} - {1'b0, layer_1_1[591:584]};
      mid_2[0] = {1'b0,layer_2_2[575:568]} - {1'b0, layer_1_2[575:568]};
      mid_2[1] = {1'b0,layer_2_2[583:576]} - {1'b0, layer_1_2[583:576]};
      mid_2[2] = {1'b0,layer_2_2[591:584]} - {1'b0, layer_1_2[591:584]};
      btm_0[0] = {1'b0,layer_3_0[575:568]} - {1'b0, layer_2_0[575:568]};
      btm_0[1] = {1'b0,layer_3_0[583:576]} - {1'b0, layer_2_0[583:576]};
      btm_0[2] = {1'b0,layer_3_0[591:584]} - {1'b0, layer_2_0[591:584]};
      btm_1[0] = {1'b0,layer_3_1[575:568]} - {1'b0, layer_2_1[575:568]};
      btm_1[1] = {1'b0,layer_3_1[583:576]} - {1'b0, layer_2_1[583:576]};
      btm_1[2] = {1'b0,layer_3_1[591:584]} - {1'b0, layer_2_1[591:584]};
      btm_2[0] = {1'b0,layer_3_2[575:568]} - {1'b0, layer_2_2[575:568]};
      btm_2[1] = {1'b0,layer_3_2[583:576]} - {1'b0, layer_2_2[583:576]};
      btm_2[2] = {1'b0,layer_3_2[591:584]} - {1'b0, layer_2_2[591:584]};
    end
    'd73: begin
      top_0[0] = {1'b0,layer_1_0[583:576]} - {1'b0, layer_0_0[583:576]};
      top_0[1] = {1'b0,layer_1_0[591:584]} - {1'b0, layer_0_0[591:584]};
      top_0[2] = {1'b0,layer_1_0[599:592]} - {1'b0, layer_0_0[599:592]};
      top_1[0] = {1'b0,layer_1_1[583:576]} - {1'b0, layer_0_1[583:576]};
      top_1[1] = {1'b0,layer_1_1[591:584]} - {1'b0, layer_0_1[591:584]};
      top_1[2] = {1'b0,layer_1_1[599:592]} - {1'b0, layer_0_1[599:592]};
      top_2[0] = {1'b0,layer_1_2[583:576]} - {1'b0, layer_0_2[583:576]};
      top_2[1] = {1'b0,layer_1_2[591:584]} - {1'b0, layer_0_2[591:584]};
      top_2[2] = {1'b0,layer_1_2[599:592]} - {1'b0, layer_0_2[599:592]};
      mid_0[0] = {1'b0,layer_2_0[583:576]} - {1'b0, layer_1_0[583:576]};
      mid_0[1] = {1'b0,layer_2_0[591:584]} - {1'b0, layer_1_0[591:584]};
      mid_0[2] = {1'b0,layer_2_0[599:592]} - {1'b0, layer_1_0[599:592]};
      mid_1[0] = {1'b0,layer_2_1[583:576]} - {1'b0, layer_1_1[583:576]};
      mid_1[1] = {1'b0,layer_2_1[591:584]} - {1'b0, layer_1_1[591:584]};
      mid_1[2] = {1'b0,layer_2_1[599:592]} - {1'b0, layer_1_1[599:592]};
      mid_2[0] = {1'b0,layer_2_2[583:576]} - {1'b0, layer_1_2[583:576]};
      mid_2[1] = {1'b0,layer_2_2[591:584]} - {1'b0, layer_1_2[591:584]};
      mid_2[2] = {1'b0,layer_2_2[599:592]} - {1'b0, layer_1_2[599:592]};
      btm_0[0] = {1'b0,layer_3_0[583:576]} - {1'b0, layer_2_0[583:576]};
      btm_0[1] = {1'b0,layer_3_0[591:584]} - {1'b0, layer_2_0[591:584]};
      btm_0[2] = {1'b0,layer_3_0[599:592]} - {1'b0, layer_2_0[599:592]};
      btm_1[0] = {1'b0,layer_3_1[583:576]} - {1'b0, layer_2_1[583:576]};
      btm_1[1] = {1'b0,layer_3_1[591:584]} - {1'b0, layer_2_1[591:584]};
      btm_1[2] = {1'b0,layer_3_1[599:592]} - {1'b0, layer_2_1[599:592]};
      btm_2[0] = {1'b0,layer_3_2[583:576]} - {1'b0, layer_2_2[583:576]};
      btm_2[1] = {1'b0,layer_3_2[591:584]} - {1'b0, layer_2_2[591:584]};
      btm_2[2] = {1'b0,layer_3_2[599:592]} - {1'b0, layer_2_2[599:592]};
    end
    'd74: begin
      top_0[0] = {1'b0,layer_1_0[591:584]} - {1'b0, layer_0_0[591:584]};
      top_0[1] = {1'b0,layer_1_0[599:592]} - {1'b0, layer_0_0[599:592]};
      top_0[2] = {1'b0,layer_1_0[607:600]} - {1'b0, layer_0_0[607:600]};
      top_1[0] = {1'b0,layer_1_1[591:584]} - {1'b0, layer_0_1[591:584]};
      top_1[1] = {1'b0,layer_1_1[599:592]} - {1'b0, layer_0_1[599:592]};
      top_1[2] = {1'b0,layer_1_1[607:600]} - {1'b0, layer_0_1[607:600]};
      top_2[0] = {1'b0,layer_1_2[591:584]} - {1'b0, layer_0_2[591:584]};
      top_2[1] = {1'b0,layer_1_2[599:592]} - {1'b0, layer_0_2[599:592]};
      top_2[2] = {1'b0,layer_1_2[607:600]} - {1'b0, layer_0_2[607:600]};
      mid_0[0] = {1'b0,layer_2_0[591:584]} - {1'b0, layer_1_0[591:584]};
      mid_0[1] = {1'b0,layer_2_0[599:592]} - {1'b0, layer_1_0[599:592]};
      mid_0[2] = {1'b0,layer_2_0[607:600]} - {1'b0, layer_1_0[607:600]};
      mid_1[0] = {1'b0,layer_2_1[591:584]} - {1'b0, layer_1_1[591:584]};
      mid_1[1] = {1'b0,layer_2_1[599:592]} - {1'b0, layer_1_1[599:592]};
      mid_1[2] = {1'b0,layer_2_1[607:600]} - {1'b0, layer_1_1[607:600]};
      mid_2[0] = {1'b0,layer_2_2[591:584]} - {1'b0, layer_1_2[591:584]};
      mid_2[1] = {1'b0,layer_2_2[599:592]} - {1'b0, layer_1_2[599:592]};
      mid_2[2] = {1'b0,layer_2_2[607:600]} - {1'b0, layer_1_2[607:600]};
      btm_0[0] = {1'b0,layer_3_0[591:584]} - {1'b0, layer_2_0[591:584]};
      btm_0[1] = {1'b0,layer_3_0[599:592]} - {1'b0, layer_2_0[599:592]};
      btm_0[2] = {1'b0,layer_3_0[607:600]} - {1'b0, layer_2_0[607:600]};
      btm_1[0] = {1'b0,layer_3_1[591:584]} - {1'b0, layer_2_1[591:584]};
      btm_1[1] = {1'b0,layer_3_1[599:592]} - {1'b0, layer_2_1[599:592]};
      btm_1[2] = {1'b0,layer_3_1[607:600]} - {1'b0, layer_2_1[607:600]};
      btm_2[0] = {1'b0,layer_3_2[591:584]} - {1'b0, layer_2_2[591:584]};
      btm_2[1] = {1'b0,layer_3_2[599:592]} - {1'b0, layer_2_2[599:592]};
      btm_2[2] = {1'b0,layer_3_2[607:600]} - {1'b0, layer_2_2[607:600]};
    end
    'd75: begin
      top_0[0] = {1'b0,layer_1_0[599:592]} - {1'b0, layer_0_0[599:592]};
      top_0[1] = {1'b0,layer_1_0[607:600]} - {1'b0, layer_0_0[607:600]};
      top_0[2] = {1'b0,layer_1_0[615:608]} - {1'b0, layer_0_0[615:608]};
      top_1[0] = {1'b0,layer_1_1[599:592]} - {1'b0, layer_0_1[599:592]};
      top_1[1] = {1'b0,layer_1_1[607:600]} - {1'b0, layer_0_1[607:600]};
      top_1[2] = {1'b0,layer_1_1[615:608]} - {1'b0, layer_0_1[615:608]};
      top_2[0] = {1'b0,layer_1_2[599:592]} - {1'b0, layer_0_2[599:592]};
      top_2[1] = {1'b0,layer_1_2[607:600]} - {1'b0, layer_0_2[607:600]};
      top_2[2] = {1'b0,layer_1_2[615:608]} - {1'b0, layer_0_2[615:608]};
      mid_0[0] = {1'b0,layer_2_0[599:592]} - {1'b0, layer_1_0[599:592]};
      mid_0[1] = {1'b0,layer_2_0[607:600]} - {1'b0, layer_1_0[607:600]};
      mid_0[2] = {1'b0,layer_2_0[615:608]} - {1'b0, layer_1_0[615:608]};
      mid_1[0] = {1'b0,layer_2_1[599:592]} - {1'b0, layer_1_1[599:592]};
      mid_1[1] = {1'b0,layer_2_1[607:600]} - {1'b0, layer_1_1[607:600]};
      mid_1[2] = {1'b0,layer_2_1[615:608]} - {1'b0, layer_1_1[615:608]};
      mid_2[0] = {1'b0,layer_2_2[599:592]} - {1'b0, layer_1_2[599:592]};
      mid_2[1] = {1'b0,layer_2_2[607:600]} - {1'b0, layer_1_2[607:600]};
      mid_2[2] = {1'b0,layer_2_2[615:608]} - {1'b0, layer_1_2[615:608]};
      btm_0[0] = {1'b0,layer_3_0[599:592]} - {1'b0, layer_2_0[599:592]};
      btm_0[1] = {1'b0,layer_3_0[607:600]} - {1'b0, layer_2_0[607:600]};
      btm_0[2] = {1'b0,layer_3_0[615:608]} - {1'b0, layer_2_0[615:608]};
      btm_1[0] = {1'b0,layer_3_1[599:592]} - {1'b0, layer_2_1[599:592]};
      btm_1[1] = {1'b0,layer_3_1[607:600]} - {1'b0, layer_2_1[607:600]};
      btm_1[2] = {1'b0,layer_3_1[615:608]} - {1'b0, layer_2_1[615:608]};
      btm_2[0] = {1'b0,layer_3_2[599:592]} - {1'b0, layer_2_2[599:592]};
      btm_2[1] = {1'b0,layer_3_2[607:600]} - {1'b0, layer_2_2[607:600]};
      btm_2[2] = {1'b0,layer_3_2[615:608]} - {1'b0, layer_2_2[615:608]};
    end
    'd76: begin
      top_0[0] = {1'b0,layer_1_0[607:600]} - {1'b0, layer_0_0[607:600]};
      top_0[1] = {1'b0,layer_1_0[615:608]} - {1'b0, layer_0_0[615:608]};
      top_0[2] = {1'b0,layer_1_0[623:616]} - {1'b0, layer_0_0[623:616]};
      top_1[0] = {1'b0,layer_1_1[607:600]} - {1'b0, layer_0_1[607:600]};
      top_1[1] = {1'b0,layer_1_1[615:608]} - {1'b0, layer_0_1[615:608]};
      top_1[2] = {1'b0,layer_1_1[623:616]} - {1'b0, layer_0_1[623:616]};
      top_2[0] = {1'b0,layer_1_2[607:600]} - {1'b0, layer_0_2[607:600]};
      top_2[1] = {1'b0,layer_1_2[615:608]} - {1'b0, layer_0_2[615:608]};
      top_2[2] = {1'b0,layer_1_2[623:616]} - {1'b0, layer_0_2[623:616]};
      mid_0[0] = {1'b0,layer_2_0[607:600]} - {1'b0, layer_1_0[607:600]};
      mid_0[1] = {1'b0,layer_2_0[615:608]} - {1'b0, layer_1_0[615:608]};
      mid_0[2] = {1'b0,layer_2_0[623:616]} - {1'b0, layer_1_0[623:616]};
      mid_1[0] = {1'b0,layer_2_1[607:600]} - {1'b0, layer_1_1[607:600]};
      mid_1[1] = {1'b0,layer_2_1[615:608]} - {1'b0, layer_1_1[615:608]};
      mid_1[2] = {1'b0,layer_2_1[623:616]} - {1'b0, layer_1_1[623:616]};
      mid_2[0] = {1'b0,layer_2_2[607:600]} - {1'b0, layer_1_2[607:600]};
      mid_2[1] = {1'b0,layer_2_2[615:608]} - {1'b0, layer_1_2[615:608]};
      mid_2[2] = {1'b0,layer_2_2[623:616]} - {1'b0, layer_1_2[623:616]};
      btm_0[0] = {1'b0,layer_3_0[607:600]} - {1'b0, layer_2_0[607:600]};
      btm_0[1] = {1'b0,layer_3_0[615:608]} - {1'b0, layer_2_0[615:608]};
      btm_0[2] = {1'b0,layer_3_0[623:616]} - {1'b0, layer_2_0[623:616]};
      btm_1[0] = {1'b0,layer_3_1[607:600]} - {1'b0, layer_2_1[607:600]};
      btm_1[1] = {1'b0,layer_3_1[615:608]} - {1'b0, layer_2_1[615:608]};
      btm_1[2] = {1'b0,layer_3_1[623:616]} - {1'b0, layer_2_1[623:616]};
      btm_2[0] = {1'b0,layer_3_2[607:600]} - {1'b0, layer_2_2[607:600]};
      btm_2[1] = {1'b0,layer_3_2[615:608]} - {1'b0, layer_2_2[615:608]};
      btm_2[2] = {1'b0,layer_3_2[623:616]} - {1'b0, layer_2_2[623:616]};
    end
    'd77: begin
      top_0[0] = {1'b0,layer_1_0[615:608]} - {1'b0, layer_0_0[615:608]};
      top_0[1] = {1'b0,layer_1_0[623:616]} - {1'b0, layer_0_0[623:616]};
      top_0[2] = {1'b0,layer_1_0[631:624]} - {1'b0, layer_0_0[631:624]};
      top_1[0] = {1'b0,layer_1_1[615:608]} - {1'b0, layer_0_1[615:608]};
      top_1[1] = {1'b0,layer_1_1[623:616]} - {1'b0, layer_0_1[623:616]};
      top_1[2] = {1'b0,layer_1_1[631:624]} - {1'b0, layer_0_1[631:624]};
      top_2[0] = {1'b0,layer_1_2[615:608]} - {1'b0, layer_0_2[615:608]};
      top_2[1] = {1'b0,layer_1_2[623:616]} - {1'b0, layer_0_2[623:616]};
      top_2[2] = {1'b0,layer_1_2[631:624]} - {1'b0, layer_0_2[631:624]};
      mid_0[0] = {1'b0,layer_2_0[615:608]} - {1'b0, layer_1_0[615:608]};
      mid_0[1] = {1'b0,layer_2_0[623:616]} - {1'b0, layer_1_0[623:616]};
      mid_0[2] = {1'b0,layer_2_0[631:624]} - {1'b0, layer_1_0[631:624]};
      mid_1[0] = {1'b0,layer_2_1[615:608]} - {1'b0, layer_1_1[615:608]};
      mid_1[1] = {1'b0,layer_2_1[623:616]} - {1'b0, layer_1_1[623:616]};
      mid_1[2] = {1'b0,layer_2_1[631:624]} - {1'b0, layer_1_1[631:624]};
      mid_2[0] = {1'b0,layer_2_2[615:608]} - {1'b0, layer_1_2[615:608]};
      mid_2[1] = {1'b0,layer_2_2[623:616]} - {1'b0, layer_1_2[623:616]};
      mid_2[2] = {1'b0,layer_2_2[631:624]} - {1'b0, layer_1_2[631:624]};
      btm_0[0] = {1'b0,layer_3_0[615:608]} - {1'b0, layer_2_0[615:608]};
      btm_0[1] = {1'b0,layer_3_0[623:616]} - {1'b0, layer_2_0[623:616]};
      btm_0[2] = {1'b0,layer_3_0[631:624]} - {1'b0, layer_2_0[631:624]};
      btm_1[0] = {1'b0,layer_3_1[615:608]} - {1'b0, layer_2_1[615:608]};
      btm_1[1] = {1'b0,layer_3_1[623:616]} - {1'b0, layer_2_1[623:616]};
      btm_1[2] = {1'b0,layer_3_1[631:624]} - {1'b0, layer_2_1[631:624]};
      btm_2[0] = {1'b0,layer_3_2[615:608]} - {1'b0, layer_2_2[615:608]};
      btm_2[1] = {1'b0,layer_3_2[623:616]} - {1'b0, layer_2_2[623:616]};
      btm_2[2] = {1'b0,layer_3_2[631:624]} - {1'b0, layer_2_2[631:624]};
    end
    'd78: begin
      top_0[0] = {1'b0,layer_1_0[623:616]} - {1'b0, layer_0_0[623:616]};
      top_0[1] = {1'b0,layer_1_0[631:624]} - {1'b0, layer_0_0[631:624]};
      top_0[2] = {1'b0,layer_1_0[639:632]} - {1'b0, layer_0_0[639:632]};
      top_1[0] = {1'b0,layer_1_1[623:616]} - {1'b0, layer_0_1[623:616]};
      top_1[1] = {1'b0,layer_1_1[631:624]} - {1'b0, layer_0_1[631:624]};
      top_1[2] = {1'b0,layer_1_1[639:632]} - {1'b0, layer_0_1[639:632]};
      top_2[0] = {1'b0,layer_1_2[623:616]} - {1'b0, layer_0_2[623:616]};
      top_2[1] = {1'b0,layer_1_2[631:624]} - {1'b0, layer_0_2[631:624]};
      top_2[2] = {1'b0,layer_1_2[639:632]} - {1'b0, layer_0_2[639:632]};
      mid_0[0] = {1'b0,layer_2_0[623:616]} - {1'b0, layer_1_0[623:616]};
      mid_0[1] = {1'b0,layer_2_0[631:624]} - {1'b0, layer_1_0[631:624]};
      mid_0[2] = {1'b0,layer_2_0[639:632]} - {1'b0, layer_1_0[639:632]};
      mid_1[0] = {1'b0,layer_2_1[623:616]} - {1'b0, layer_1_1[623:616]};
      mid_1[1] = {1'b0,layer_2_1[631:624]} - {1'b0, layer_1_1[631:624]};
      mid_1[2] = {1'b0,layer_2_1[639:632]} - {1'b0, layer_1_1[639:632]};
      mid_2[0] = {1'b0,layer_2_2[623:616]} - {1'b0, layer_1_2[623:616]};
      mid_2[1] = {1'b0,layer_2_2[631:624]} - {1'b0, layer_1_2[631:624]};
      mid_2[2] = {1'b0,layer_2_2[639:632]} - {1'b0, layer_1_2[639:632]};
      btm_0[0] = {1'b0,layer_3_0[623:616]} - {1'b0, layer_2_0[623:616]};
      btm_0[1] = {1'b0,layer_3_0[631:624]} - {1'b0, layer_2_0[631:624]};
      btm_0[2] = {1'b0,layer_3_0[639:632]} - {1'b0, layer_2_0[639:632]};
      btm_1[0] = {1'b0,layer_3_1[623:616]} - {1'b0, layer_2_1[623:616]};
      btm_1[1] = {1'b0,layer_3_1[631:624]} - {1'b0, layer_2_1[631:624]};
      btm_1[2] = {1'b0,layer_3_1[639:632]} - {1'b0, layer_2_1[639:632]};
      btm_2[0] = {1'b0,layer_3_2[623:616]} - {1'b0, layer_2_2[623:616]};
      btm_2[1] = {1'b0,layer_3_2[631:624]} - {1'b0, layer_2_2[631:624]};
      btm_2[2] = {1'b0,layer_3_2[639:632]} - {1'b0, layer_2_2[639:632]};
    end
    'd79: begin
      top_0[0] = {1'b0,layer_1_0[631:624]} - {1'b0, layer_0_0[631:624]};
      top_0[1] = {1'b0,layer_1_0[639:632]} - {1'b0, layer_0_0[639:632]};
      top_0[2] = {1'b0,layer_1_0[647:640]} - {1'b0, layer_0_0[647:640]};
      top_1[0] = {1'b0,layer_1_1[631:624]} - {1'b0, layer_0_1[631:624]};
      top_1[1] = {1'b0,layer_1_1[639:632]} - {1'b0, layer_0_1[639:632]};
      top_1[2] = {1'b0,layer_1_1[647:640]} - {1'b0, layer_0_1[647:640]};
      top_2[0] = {1'b0,layer_1_2[631:624]} - {1'b0, layer_0_2[631:624]};
      top_2[1] = {1'b0,layer_1_2[639:632]} - {1'b0, layer_0_2[639:632]};
      top_2[2] = {1'b0,layer_1_2[647:640]} - {1'b0, layer_0_2[647:640]};
      mid_0[0] = {1'b0,layer_2_0[631:624]} - {1'b0, layer_1_0[631:624]};
      mid_0[1] = {1'b0,layer_2_0[639:632]} - {1'b0, layer_1_0[639:632]};
      mid_0[2] = {1'b0,layer_2_0[647:640]} - {1'b0, layer_1_0[647:640]};
      mid_1[0] = {1'b0,layer_2_1[631:624]} - {1'b0, layer_1_1[631:624]};
      mid_1[1] = {1'b0,layer_2_1[639:632]} - {1'b0, layer_1_1[639:632]};
      mid_1[2] = {1'b0,layer_2_1[647:640]} - {1'b0, layer_1_1[647:640]};
      mid_2[0] = {1'b0,layer_2_2[631:624]} - {1'b0, layer_1_2[631:624]};
      mid_2[1] = {1'b0,layer_2_2[639:632]} - {1'b0, layer_1_2[639:632]};
      mid_2[2] = {1'b0,layer_2_2[647:640]} - {1'b0, layer_1_2[647:640]};
      btm_0[0] = {1'b0,layer_3_0[631:624]} - {1'b0, layer_2_0[631:624]};
      btm_0[1] = {1'b0,layer_3_0[639:632]} - {1'b0, layer_2_0[639:632]};
      btm_0[2] = {1'b0,layer_3_0[647:640]} - {1'b0, layer_2_0[647:640]};
      btm_1[0] = {1'b0,layer_3_1[631:624]} - {1'b0, layer_2_1[631:624]};
      btm_1[1] = {1'b0,layer_3_1[639:632]} - {1'b0, layer_2_1[639:632]};
      btm_1[2] = {1'b0,layer_3_1[647:640]} - {1'b0, layer_2_1[647:640]};
      btm_2[0] = {1'b0,layer_3_2[631:624]} - {1'b0, layer_2_2[631:624]};
      btm_2[1] = {1'b0,layer_3_2[639:632]} - {1'b0, layer_2_2[639:632]};
      btm_2[2] = {1'b0,layer_3_2[647:640]} - {1'b0, layer_2_2[647:640]};
    end
    'd80: begin
      top_0[0] = {1'b0,layer_1_0[639:632]} - {1'b0, layer_0_0[639:632]};
      top_0[1] = {1'b0,layer_1_0[647:640]} - {1'b0, layer_0_0[647:640]};
      top_0[2] = {1'b0,layer_1_0[655:648]} - {1'b0, layer_0_0[655:648]};
      top_1[0] = {1'b0,layer_1_1[639:632]} - {1'b0, layer_0_1[639:632]};
      top_1[1] = {1'b0,layer_1_1[647:640]} - {1'b0, layer_0_1[647:640]};
      top_1[2] = {1'b0,layer_1_1[655:648]} - {1'b0, layer_0_1[655:648]};
      top_2[0] = {1'b0,layer_1_2[639:632]} - {1'b0, layer_0_2[639:632]};
      top_2[1] = {1'b0,layer_1_2[647:640]} - {1'b0, layer_0_2[647:640]};
      top_2[2] = {1'b0,layer_1_2[655:648]} - {1'b0, layer_0_2[655:648]};
      mid_0[0] = {1'b0,layer_2_0[639:632]} - {1'b0, layer_1_0[639:632]};
      mid_0[1] = {1'b0,layer_2_0[647:640]} - {1'b0, layer_1_0[647:640]};
      mid_0[2] = {1'b0,layer_2_0[655:648]} - {1'b0, layer_1_0[655:648]};
      mid_1[0] = {1'b0,layer_2_1[639:632]} - {1'b0, layer_1_1[639:632]};
      mid_1[1] = {1'b0,layer_2_1[647:640]} - {1'b0, layer_1_1[647:640]};
      mid_1[2] = {1'b0,layer_2_1[655:648]} - {1'b0, layer_1_1[655:648]};
      mid_2[0] = {1'b0,layer_2_2[639:632]} - {1'b0, layer_1_2[639:632]};
      mid_2[1] = {1'b0,layer_2_2[647:640]} - {1'b0, layer_1_2[647:640]};
      mid_2[2] = {1'b0,layer_2_2[655:648]} - {1'b0, layer_1_2[655:648]};
      btm_0[0] = {1'b0,layer_3_0[639:632]} - {1'b0, layer_2_0[639:632]};
      btm_0[1] = {1'b0,layer_3_0[647:640]} - {1'b0, layer_2_0[647:640]};
      btm_0[2] = {1'b0,layer_3_0[655:648]} - {1'b0, layer_2_0[655:648]};
      btm_1[0] = {1'b0,layer_3_1[639:632]} - {1'b0, layer_2_1[639:632]};
      btm_1[1] = {1'b0,layer_3_1[647:640]} - {1'b0, layer_2_1[647:640]};
      btm_1[2] = {1'b0,layer_3_1[655:648]} - {1'b0, layer_2_1[655:648]};
      btm_2[0] = {1'b0,layer_3_2[639:632]} - {1'b0, layer_2_2[639:632]};
      btm_2[1] = {1'b0,layer_3_2[647:640]} - {1'b0, layer_2_2[647:640]};
      btm_2[2] = {1'b0,layer_3_2[655:648]} - {1'b0, layer_2_2[655:648]};
    end
    'd81: begin
      top_0[0] = {1'b0,layer_1_0[647:640]} - {1'b0, layer_0_0[647:640]};
      top_0[1] = {1'b0,layer_1_0[655:648]} - {1'b0, layer_0_0[655:648]};
      top_0[2] = {1'b0,layer_1_0[663:656]} - {1'b0, layer_0_0[663:656]};
      top_1[0] = {1'b0,layer_1_1[647:640]} - {1'b0, layer_0_1[647:640]};
      top_1[1] = {1'b0,layer_1_1[655:648]} - {1'b0, layer_0_1[655:648]};
      top_1[2] = {1'b0,layer_1_1[663:656]} - {1'b0, layer_0_1[663:656]};
      top_2[0] = {1'b0,layer_1_2[647:640]} - {1'b0, layer_0_2[647:640]};
      top_2[1] = {1'b0,layer_1_2[655:648]} - {1'b0, layer_0_2[655:648]};
      top_2[2] = {1'b0,layer_1_2[663:656]} - {1'b0, layer_0_2[663:656]};
      mid_0[0] = {1'b0,layer_2_0[647:640]} - {1'b0, layer_1_0[647:640]};
      mid_0[1] = {1'b0,layer_2_0[655:648]} - {1'b0, layer_1_0[655:648]};
      mid_0[2] = {1'b0,layer_2_0[663:656]} - {1'b0, layer_1_0[663:656]};
      mid_1[0] = {1'b0,layer_2_1[647:640]} - {1'b0, layer_1_1[647:640]};
      mid_1[1] = {1'b0,layer_2_1[655:648]} - {1'b0, layer_1_1[655:648]};
      mid_1[2] = {1'b0,layer_2_1[663:656]} - {1'b0, layer_1_1[663:656]};
      mid_2[0] = {1'b0,layer_2_2[647:640]} - {1'b0, layer_1_2[647:640]};
      mid_2[1] = {1'b0,layer_2_2[655:648]} - {1'b0, layer_1_2[655:648]};
      mid_2[2] = {1'b0,layer_2_2[663:656]} - {1'b0, layer_1_2[663:656]};
      btm_0[0] = {1'b0,layer_3_0[647:640]} - {1'b0, layer_2_0[647:640]};
      btm_0[1] = {1'b0,layer_3_0[655:648]} - {1'b0, layer_2_0[655:648]};
      btm_0[2] = {1'b0,layer_3_0[663:656]} - {1'b0, layer_2_0[663:656]};
      btm_1[0] = {1'b0,layer_3_1[647:640]} - {1'b0, layer_2_1[647:640]};
      btm_1[1] = {1'b0,layer_3_1[655:648]} - {1'b0, layer_2_1[655:648]};
      btm_1[2] = {1'b0,layer_3_1[663:656]} - {1'b0, layer_2_1[663:656]};
      btm_2[0] = {1'b0,layer_3_2[647:640]} - {1'b0, layer_2_2[647:640]};
      btm_2[1] = {1'b0,layer_3_2[655:648]} - {1'b0, layer_2_2[655:648]};
      btm_2[2] = {1'b0,layer_3_2[663:656]} - {1'b0, layer_2_2[663:656]};
    end
    'd82: begin
      top_0[0] = {1'b0,layer_1_0[655:648]} - {1'b0, layer_0_0[655:648]};
      top_0[1] = {1'b0,layer_1_0[663:656]} - {1'b0, layer_0_0[663:656]};
      top_0[2] = {1'b0,layer_1_0[671:664]} - {1'b0, layer_0_0[671:664]};
      top_1[0] = {1'b0,layer_1_1[655:648]} - {1'b0, layer_0_1[655:648]};
      top_1[1] = {1'b0,layer_1_1[663:656]} - {1'b0, layer_0_1[663:656]};
      top_1[2] = {1'b0,layer_1_1[671:664]} - {1'b0, layer_0_1[671:664]};
      top_2[0] = {1'b0,layer_1_2[655:648]} - {1'b0, layer_0_2[655:648]};
      top_2[1] = {1'b0,layer_1_2[663:656]} - {1'b0, layer_0_2[663:656]};
      top_2[2] = {1'b0,layer_1_2[671:664]} - {1'b0, layer_0_2[671:664]};
      mid_0[0] = {1'b0,layer_2_0[655:648]} - {1'b0, layer_1_0[655:648]};
      mid_0[1] = {1'b0,layer_2_0[663:656]} - {1'b0, layer_1_0[663:656]};
      mid_0[2] = {1'b0,layer_2_0[671:664]} - {1'b0, layer_1_0[671:664]};
      mid_1[0] = {1'b0,layer_2_1[655:648]} - {1'b0, layer_1_1[655:648]};
      mid_1[1] = {1'b0,layer_2_1[663:656]} - {1'b0, layer_1_1[663:656]};
      mid_1[2] = {1'b0,layer_2_1[671:664]} - {1'b0, layer_1_1[671:664]};
      mid_2[0] = {1'b0,layer_2_2[655:648]} - {1'b0, layer_1_2[655:648]};
      mid_2[1] = {1'b0,layer_2_2[663:656]} - {1'b0, layer_1_2[663:656]};
      mid_2[2] = {1'b0,layer_2_2[671:664]} - {1'b0, layer_1_2[671:664]};
      btm_0[0] = {1'b0,layer_3_0[655:648]} - {1'b0, layer_2_0[655:648]};
      btm_0[1] = {1'b0,layer_3_0[663:656]} - {1'b0, layer_2_0[663:656]};
      btm_0[2] = {1'b0,layer_3_0[671:664]} - {1'b0, layer_2_0[671:664]};
      btm_1[0] = {1'b0,layer_3_1[655:648]} - {1'b0, layer_2_1[655:648]};
      btm_1[1] = {1'b0,layer_3_1[663:656]} - {1'b0, layer_2_1[663:656]};
      btm_1[2] = {1'b0,layer_3_1[671:664]} - {1'b0, layer_2_1[671:664]};
      btm_2[0] = {1'b0,layer_3_2[655:648]} - {1'b0, layer_2_2[655:648]};
      btm_2[1] = {1'b0,layer_3_2[663:656]} - {1'b0, layer_2_2[663:656]};
      btm_2[2] = {1'b0,layer_3_2[671:664]} - {1'b0, layer_2_2[671:664]};
    end
    'd83: begin
      top_0[0] = {1'b0,layer_1_0[663:656]} - {1'b0, layer_0_0[663:656]};
      top_0[1] = {1'b0,layer_1_0[671:664]} - {1'b0, layer_0_0[671:664]};
      top_0[2] = {1'b0,layer_1_0[679:672]} - {1'b0, layer_0_0[679:672]};
      top_1[0] = {1'b0,layer_1_1[663:656]} - {1'b0, layer_0_1[663:656]};
      top_1[1] = {1'b0,layer_1_1[671:664]} - {1'b0, layer_0_1[671:664]};
      top_1[2] = {1'b0,layer_1_1[679:672]} - {1'b0, layer_0_1[679:672]};
      top_2[0] = {1'b0,layer_1_2[663:656]} - {1'b0, layer_0_2[663:656]};
      top_2[1] = {1'b0,layer_1_2[671:664]} - {1'b0, layer_0_2[671:664]};
      top_2[2] = {1'b0,layer_1_2[679:672]} - {1'b0, layer_0_2[679:672]};
      mid_0[0] = {1'b0,layer_2_0[663:656]} - {1'b0, layer_1_0[663:656]};
      mid_0[1] = {1'b0,layer_2_0[671:664]} - {1'b0, layer_1_0[671:664]};
      mid_0[2] = {1'b0,layer_2_0[679:672]} - {1'b0, layer_1_0[679:672]};
      mid_1[0] = {1'b0,layer_2_1[663:656]} - {1'b0, layer_1_1[663:656]};
      mid_1[1] = {1'b0,layer_2_1[671:664]} - {1'b0, layer_1_1[671:664]};
      mid_1[2] = {1'b0,layer_2_1[679:672]} - {1'b0, layer_1_1[679:672]};
      mid_2[0] = {1'b0,layer_2_2[663:656]} - {1'b0, layer_1_2[663:656]};
      mid_2[1] = {1'b0,layer_2_2[671:664]} - {1'b0, layer_1_2[671:664]};
      mid_2[2] = {1'b0,layer_2_2[679:672]} - {1'b0, layer_1_2[679:672]};
      btm_0[0] = {1'b0,layer_3_0[663:656]} - {1'b0, layer_2_0[663:656]};
      btm_0[1] = {1'b0,layer_3_0[671:664]} - {1'b0, layer_2_0[671:664]};
      btm_0[2] = {1'b0,layer_3_0[679:672]} - {1'b0, layer_2_0[679:672]};
      btm_1[0] = {1'b0,layer_3_1[663:656]} - {1'b0, layer_2_1[663:656]};
      btm_1[1] = {1'b0,layer_3_1[671:664]} - {1'b0, layer_2_1[671:664]};
      btm_1[2] = {1'b0,layer_3_1[679:672]} - {1'b0, layer_2_1[679:672]};
      btm_2[0] = {1'b0,layer_3_2[663:656]} - {1'b0, layer_2_2[663:656]};
      btm_2[1] = {1'b0,layer_3_2[671:664]} - {1'b0, layer_2_2[671:664]};
      btm_2[2] = {1'b0,layer_3_2[679:672]} - {1'b0, layer_2_2[679:672]};
    end
    'd84: begin
      top_0[0] = {1'b0,layer_1_0[671:664]} - {1'b0, layer_0_0[671:664]};
      top_0[1] = {1'b0,layer_1_0[679:672]} - {1'b0, layer_0_0[679:672]};
      top_0[2] = {1'b0,layer_1_0[687:680]} - {1'b0, layer_0_0[687:680]};
      top_1[0] = {1'b0,layer_1_1[671:664]} - {1'b0, layer_0_1[671:664]};
      top_1[1] = {1'b0,layer_1_1[679:672]} - {1'b0, layer_0_1[679:672]};
      top_1[2] = {1'b0,layer_1_1[687:680]} - {1'b0, layer_0_1[687:680]};
      top_2[0] = {1'b0,layer_1_2[671:664]} - {1'b0, layer_0_2[671:664]};
      top_2[1] = {1'b0,layer_1_2[679:672]} - {1'b0, layer_0_2[679:672]};
      top_2[2] = {1'b0,layer_1_2[687:680]} - {1'b0, layer_0_2[687:680]};
      mid_0[0] = {1'b0,layer_2_0[671:664]} - {1'b0, layer_1_0[671:664]};
      mid_0[1] = {1'b0,layer_2_0[679:672]} - {1'b0, layer_1_0[679:672]};
      mid_0[2] = {1'b0,layer_2_0[687:680]} - {1'b0, layer_1_0[687:680]};
      mid_1[0] = {1'b0,layer_2_1[671:664]} - {1'b0, layer_1_1[671:664]};
      mid_1[1] = {1'b0,layer_2_1[679:672]} - {1'b0, layer_1_1[679:672]};
      mid_1[2] = {1'b0,layer_2_1[687:680]} - {1'b0, layer_1_1[687:680]};
      mid_2[0] = {1'b0,layer_2_2[671:664]} - {1'b0, layer_1_2[671:664]};
      mid_2[1] = {1'b0,layer_2_2[679:672]} - {1'b0, layer_1_2[679:672]};
      mid_2[2] = {1'b0,layer_2_2[687:680]} - {1'b0, layer_1_2[687:680]};
      btm_0[0] = {1'b0,layer_3_0[671:664]} - {1'b0, layer_2_0[671:664]};
      btm_0[1] = {1'b0,layer_3_0[679:672]} - {1'b0, layer_2_0[679:672]};
      btm_0[2] = {1'b0,layer_3_0[687:680]} - {1'b0, layer_2_0[687:680]};
      btm_1[0] = {1'b0,layer_3_1[671:664]} - {1'b0, layer_2_1[671:664]};
      btm_1[1] = {1'b0,layer_3_1[679:672]} - {1'b0, layer_2_1[679:672]};
      btm_1[2] = {1'b0,layer_3_1[687:680]} - {1'b0, layer_2_1[687:680]};
      btm_2[0] = {1'b0,layer_3_2[671:664]} - {1'b0, layer_2_2[671:664]};
      btm_2[1] = {1'b0,layer_3_2[679:672]} - {1'b0, layer_2_2[679:672]};
      btm_2[2] = {1'b0,layer_3_2[687:680]} - {1'b0, layer_2_2[687:680]};
    end
    'd85: begin
      top_0[0] = {1'b0,layer_1_0[679:672]} - {1'b0, layer_0_0[679:672]};
      top_0[1] = {1'b0,layer_1_0[687:680]} - {1'b0, layer_0_0[687:680]};
      top_0[2] = {1'b0,layer_1_0[695:688]} - {1'b0, layer_0_0[695:688]};
      top_1[0] = {1'b0,layer_1_1[679:672]} - {1'b0, layer_0_1[679:672]};
      top_1[1] = {1'b0,layer_1_1[687:680]} - {1'b0, layer_0_1[687:680]};
      top_1[2] = {1'b0,layer_1_1[695:688]} - {1'b0, layer_0_1[695:688]};
      top_2[0] = {1'b0,layer_1_2[679:672]} - {1'b0, layer_0_2[679:672]};
      top_2[1] = {1'b0,layer_1_2[687:680]} - {1'b0, layer_0_2[687:680]};
      top_2[2] = {1'b0,layer_1_2[695:688]} - {1'b0, layer_0_2[695:688]};
      mid_0[0] = {1'b0,layer_2_0[679:672]} - {1'b0, layer_1_0[679:672]};
      mid_0[1] = {1'b0,layer_2_0[687:680]} - {1'b0, layer_1_0[687:680]};
      mid_0[2] = {1'b0,layer_2_0[695:688]} - {1'b0, layer_1_0[695:688]};
      mid_1[0] = {1'b0,layer_2_1[679:672]} - {1'b0, layer_1_1[679:672]};
      mid_1[1] = {1'b0,layer_2_1[687:680]} - {1'b0, layer_1_1[687:680]};
      mid_1[2] = {1'b0,layer_2_1[695:688]} - {1'b0, layer_1_1[695:688]};
      mid_2[0] = {1'b0,layer_2_2[679:672]} - {1'b0, layer_1_2[679:672]};
      mid_2[1] = {1'b0,layer_2_2[687:680]} - {1'b0, layer_1_2[687:680]};
      mid_2[2] = {1'b0,layer_2_2[695:688]} - {1'b0, layer_1_2[695:688]};
      btm_0[0] = {1'b0,layer_3_0[679:672]} - {1'b0, layer_2_0[679:672]};
      btm_0[1] = {1'b0,layer_3_0[687:680]} - {1'b0, layer_2_0[687:680]};
      btm_0[2] = {1'b0,layer_3_0[695:688]} - {1'b0, layer_2_0[695:688]};
      btm_1[0] = {1'b0,layer_3_1[679:672]} - {1'b0, layer_2_1[679:672]};
      btm_1[1] = {1'b0,layer_3_1[687:680]} - {1'b0, layer_2_1[687:680]};
      btm_1[2] = {1'b0,layer_3_1[695:688]} - {1'b0, layer_2_1[695:688]};
      btm_2[0] = {1'b0,layer_3_2[679:672]} - {1'b0, layer_2_2[679:672]};
      btm_2[1] = {1'b0,layer_3_2[687:680]} - {1'b0, layer_2_2[687:680]};
      btm_2[2] = {1'b0,layer_3_2[695:688]} - {1'b0, layer_2_2[695:688]};
    end
    'd86: begin
      top_0[0] = {1'b0,layer_1_0[687:680]} - {1'b0, layer_0_0[687:680]};
      top_0[1] = {1'b0,layer_1_0[695:688]} - {1'b0, layer_0_0[695:688]};
      top_0[2] = {1'b0,layer_1_0[703:696]} - {1'b0, layer_0_0[703:696]};
      top_1[0] = {1'b0,layer_1_1[687:680]} - {1'b0, layer_0_1[687:680]};
      top_1[1] = {1'b0,layer_1_1[695:688]} - {1'b0, layer_0_1[695:688]};
      top_1[2] = {1'b0,layer_1_1[703:696]} - {1'b0, layer_0_1[703:696]};
      top_2[0] = {1'b0,layer_1_2[687:680]} - {1'b0, layer_0_2[687:680]};
      top_2[1] = {1'b0,layer_1_2[695:688]} - {1'b0, layer_0_2[695:688]};
      top_2[2] = {1'b0,layer_1_2[703:696]} - {1'b0, layer_0_2[703:696]};
      mid_0[0] = {1'b0,layer_2_0[687:680]} - {1'b0, layer_1_0[687:680]};
      mid_0[1] = {1'b0,layer_2_0[695:688]} - {1'b0, layer_1_0[695:688]};
      mid_0[2] = {1'b0,layer_2_0[703:696]} - {1'b0, layer_1_0[703:696]};
      mid_1[0] = {1'b0,layer_2_1[687:680]} - {1'b0, layer_1_1[687:680]};
      mid_1[1] = {1'b0,layer_2_1[695:688]} - {1'b0, layer_1_1[695:688]};
      mid_1[2] = {1'b0,layer_2_1[703:696]} - {1'b0, layer_1_1[703:696]};
      mid_2[0] = {1'b0,layer_2_2[687:680]} - {1'b0, layer_1_2[687:680]};
      mid_2[1] = {1'b0,layer_2_2[695:688]} - {1'b0, layer_1_2[695:688]};
      mid_2[2] = {1'b0,layer_2_2[703:696]} - {1'b0, layer_1_2[703:696]};
      btm_0[0] = {1'b0,layer_3_0[687:680]} - {1'b0, layer_2_0[687:680]};
      btm_0[1] = {1'b0,layer_3_0[695:688]} - {1'b0, layer_2_0[695:688]};
      btm_0[2] = {1'b0,layer_3_0[703:696]} - {1'b0, layer_2_0[703:696]};
      btm_1[0] = {1'b0,layer_3_1[687:680]} - {1'b0, layer_2_1[687:680]};
      btm_1[1] = {1'b0,layer_3_1[695:688]} - {1'b0, layer_2_1[695:688]};
      btm_1[2] = {1'b0,layer_3_1[703:696]} - {1'b0, layer_2_1[703:696]};
      btm_2[0] = {1'b0,layer_3_2[687:680]} - {1'b0, layer_2_2[687:680]};
      btm_2[1] = {1'b0,layer_3_2[695:688]} - {1'b0, layer_2_2[695:688]};
      btm_2[2] = {1'b0,layer_3_2[703:696]} - {1'b0, layer_2_2[703:696]};
    end
    'd87: begin
      top_0[0] = {1'b0,layer_1_0[695:688]} - {1'b0, layer_0_0[695:688]};
      top_0[1] = {1'b0,layer_1_0[703:696]} - {1'b0, layer_0_0[703:696]};
      top_0[2] = {1'b0,layer_1_0[711:704]} - {1'b0, layer_0_0[711:704]};
      top_1[0] = {1'b0,layer_1_1[695:688]} - {1'b0, layer_0_1[695:688]};
      top_1[1] = {1'b0,layer_1_1[703:696]} - {1'b0, layer_0_1[703:696]};
      top_1[2] = {1'b0,layer_1_1[711:704]} - {1'b0, layer_0_1[711:704]};
      top_2[0] = {1'b0,layer_1_2[695:688]} - {1'b0, layer_0_2[695:688]};
      top_2[1] = {1'b0,layer_1_2[703:696]} - {1'b0, layer_0_2[703:696]};
      top_2[2] = {1'b0,layer_1_2[711:704]} - {1'b0, layer_0_2[711:704]};
      mid_0[0] = {1'b0,layer_2_0[695:688]} - {1'b0, layer_1_0[695:688]};
      mid_0[1] = {1'b0,layer_2_0[703:696]} - {1'b0, layer_1_0[703:696]};
      mid_0[2] = {1'b0,layer_2_0[711:704]} - {1'b0, layer_1_0[711:704]};
      mid_1[0] = {1'b0,layer_2_1[695:688]} - {1'b0, layer_1_1[695:688]};
      mid_1[1] = {1'b0,layer_2_1[703:696]} - {1'b0, layer_1_1[703:696]};
      mid_1[2] = {1'b0,layer_2_1[711:704]} - {1'b0, layer_1_1[711:704]};
      mid_2[0] = {1'b0,layer_2_2[695:688]} - {1'b0, layer_1_2[695:688]};
      mid_2[1] = {1'b0,layer_2_2[703:696]} - {1'b0, layer_1_2[703:696]};
      mid_2[2] = {1'b0,layer_2_2[711:704]} - {1'b0, layer_1_2[711:704]};
      btm_0[0] = {1'b0,layer_3_0[695:688]} - {1'b0, layer_2_0[695:688]};
      btm_0[1] = {1'b0,layer_3_0[703:696]} - {1'b0, layer_2_0[703:696]};
      btm_0[2] = {1'b0,layer_3_0[711:704]} - {1'b0, layer_2_0[711:704]};
      btm_1[0] = {1'b0,layer_3_1[695:688]} - {1'b0, layer_2_1[695:688]};
      btm_1[1] = {1'b0,layer_3_1[703:696]} - {1'b0, layer_2_1[703:696]};
      btm_1[2] = {1'b0,layer_3_1[711:704]} - {1'b0, layer_2_1[711:704]};
      btm_2[0] = {1'b0,layer_3_2[695:688]} - {1'b0, layer_2_2[695:688]};
      btm_2[1] = {1'b0,layer_3_2[703:696]} - {1'b0, layer_2_2[703:696]};
      btm_2[2] = {1'b0,layer_3_2[711:704]} - {1'b0, layer_2_2[711:704]};
    end
    'd88: begin
      top_0[0] = {1'b0,layer_1_0[703:696]} - {1'b0, layer_0_0[703:696]};
      top_0[1] = {1'b0,layer_1_0[711:704]} - {1'b0, layer_0_0[711:704]};
      top_0[2] = {1'b0,layer_1_0[719:712]} - {1'b0, layer_0_0[719:712]};
      top_1[0] = {1'b0,layer_1_1[703:696]} - {1'b0, layer_0_1[703:696]};
      top_1[1] = {1'b0,layer_1_1[711:704]} - {1'b0, layer_0_1[711:704]};
      top_1[2] = {1'b0,layer_1_1[719:712]} - {1'b0, layer_0_1[719:712]};
      top_2[0] = {1'b0,layer_1_2[703:696]} - {1'b0, layer_0_2[703:696]};
      top_2[1] = {1'b0,layer_1_2[711:704]} - {1'b0, layer_0_2[711:704]};
      top_2[2] = {1'b0,layer_1_2[719:712]} - {1'b0, layer_0_2[719:712]};
      mid_0[0] = {1'b0,layer_2_0[703:696]} - {1'b0, layer_1_0[703:696]};
      mid_0[1] = {1'b0,layer_2_0[711:704]} - {1'b0, layer_1_0[711:704]};
      mid_0[2] = {1'b0,layer_2_0[719:712]} - {1'b0, layer_1_0[719:712]};
      mid_1[0] = {1'b0,layer_2_1[703:696]} - {1'b0, layer_1_1[703:696]};
      mid_1[1] = {1'b0,layer_2_1[711:704]} - {1'b0, layer_1_1[711:704]};
      mid_1[2] = {1'b0,layer_2_1[719:712]} - {1'b0, layer_1_1[719:712]};
      mid_2[0] = {1'b0,layer_2_2[703:696]} - {1'b0, layer_1_2[703:696]};
      mid_2[1] = {1'b0,layer_2_2[711:704]} - {1'b0, layer_1_2[711:704]};
      mid_2[2] = {1'b0,layer_2_2[719:712]} - {1'b0, layer_1_2[719:712]};
      btm_0[0] = {1'b0,layer_3_0[703:696]} - {1'b0, layer_2_0[703:696]};
      btm_0[1] = {1'b0,layer_3_0[711:704]} - {1'b0, layer_2_0[711:704]};
      btm_0[2] = {1'b0,layer_3_0[719:712]} - {1'b0, layer_2_0[719:712]};
      btm_1[0] = {1'b0,layer_3_1[703:696]} - {1'b0, layer_2_1[703:696]};
      btm_1[1] = {1'b0,layer_3_1[711:704]} - {1'b0, layer_2_1[711:704]};
      btm_1[2] = {1'b0,layer_3_1[719:712]} - {1'b0, layer_2_1[719:712]};
      btm_2[0] = {1'b0,layer_3_2[703:696]} - {1'b0, layer_2_2[703:696]};
      btm_2[1] = {1'b0,layer_3_2[711:704]} - {1'b0, layer_2_2[711:704]};
      btm_2[2] = {1'b0,layer_3_2[719:712]} - {1'b0, layer_2_2[719:712]};
    end
    'd89: begin
      top_0[0] = {1'b0,layer_1_0[711:704]} - {1'b0, layer_0_0[711:704]};
      top_0[1] = {1'b0,layer_1_0[719:712]} - {1'b0, layer_0_0[719:712]};
      top_0[2] = {1'b0,layer_1_0[727:720]} - {1'b0, layer_0_0[727:720]};
      top_1[0] = {1'b0,layer_1_1[711:704]} - {1'b0, layer_0_1[711:704]};
      top_1[1] = {1'b0,layer_1_1[719:712]} - {1'b0, layer_0_1[719:712]};
      top_1[2] = {1'b0,layer_1_1[727:720]} - {1'b0, layer_0_1[727:720]};
      top_2[0] = {1'b0,layer_1_2[711:704]} - {1'b0, layer_0_2[711:704]};
      top_2[1] = {1'b0,layer_1_2[719:712]} - {1'b0, layer_0_2[719:712]};
      top_2[2] = {1'b0,layer_1_2[727:720]} - {1'b0, layer_0_2[727:720]};
      mid_0[0] = {1'b0,layer_2_0[711:704]} - {1'b0, layer_1_0[711:704]};
      mid_0[1] = {1'b0,layer_2_0[719:712]} - {1'b0, layer_1_0[719:712]};
      mid_0[2] = {1'b0,layer_2_0[727:720]} - {1'b0, layer_1_0[727:720]};
      mid_1[0] = {1'b0,layer_2_1[711:704]} - {1'b0, layer_1_1[711:704]};
      mid_1[1] = {1'b0,layer_2_1[719:712]} - {1'b0, layer_1_1[719:712]};
      mid_1[2] = {1'b0,layer_2_1[727:720]} - {1'b0, layer_1_1[727:720]};
      mid_2[0] = {1'b0,layer_2_2[711:704]} - {1'b0, layer_1_2[711:704]};
      mid_2[1] = {1'b0,layer_2_2[719:712]} - {1'b0, layer_1_2[719:712]};
      mid_2[2] = {1'b0,layer_2_2[727:720]} - {1'b0, layer_1_2[727:720]};
      btm_0[0] = {1'b0,layer_3_0[711:704]} - {1'b0, layer_2_0[711:704]};
      btm_0[1] = {1'b0,layer_3_0[719:712]} - {1'b0, layer_2_0[719:712]};
      btm_0[2] = {1'b0,layer_3_0[727:720]} - {1'b0, layer_2_0[727:720]};
      btm_1[0] = {1'b0,layer_3_1[711:704]} - {1'b0, layer_2_1[711:704]};
      btm_1[1] = {1'b0,layer_3_1[719:712]} - {1'b0, layer_2_1[719:712]};
      btm_1[2] = {1'b0,layer_3_1[727:720]} - {1'b0, layer_2_1[727:720]};
      btm_2[0] = {1'b0,layer_3_2[711:704]} - {1'b0, layer_2_2[711:704]};
      btm_2[1] = {1'b0,layer_3_2[719:712]} - {1'b0, layer_2_2[719:712]};
      btm_2[2] = {1'b0,layer_3_2[727:720]} - {1'b0, layer_2_2[727:720]};
    end
    'd90: begin
      top_0[0] = {1'b0,layer_1_0[719:712]} - {1'b0, layer_0_0[719:712]};
      top_0[1] = {1'b0,layer_1_0[727:720]} - {1'b0, layer_0_0[727:720]};
      top_0[2] = {1'b0,layer_1_0[735:728]} - {1'b0, layer_0_0[735:728]};
      top_1[0] = {1'b0,layer_1_1[719:712]} - {1'b0, layer_0_1[719:712]};
      top_1[1] = {1'b0,layer_1_1[727:720]} - {1'b0, layer_0_1[727:720]};
      top_1[2] = {1'b0,layer_1_1[735:728]} - {1'b0, layer_0_1[735:728]};
      top_2[0] = {1'b0,layer_1_2[719:712]} - {1'b0, layer_0_2[719:712]};
      top_2[1] = {1'b0,layer_1_2[727:720]} - {1'b0, layer_0_2[727:720]};
      top_2[2] = {1'b0,layer_1_2[735:728]} - {1'b0, layer_0_2[735:728]};
      mid_0[0] = {1'b0,layer_2_0[719:712]} - {1'b0, layer_1_0[719:712]};
      mid_0[1] = {1'b0,layer_2_0[727:720]} - {1'b0, layer_1_0[727:720]};
      mid_0[2] = {1'b0,layer_2_0[735:728]} - {1'b0, layer_1_0[735:728]};
      mid_1[0] = {1'b0,layer_2_1[719:712]} - {1'b0, layer_1_1[719:712]};
      mid_1[1] = {1'b0,layer_2_1[727:720]} - {1'b0, layer_1_1[727:720]};
      mid_1[2] = {1'b0,layer_2_1[735:728]} - {1'b0, layer_1_1[735:728]};
      mid_2[0] = {1'b0,layer_2_2[719:712]} - {1'b0, layer_1_2[719:712]};
      mid_2[1] = {1'b0,layer_2_2[727:720]} - {1'b0, layer_1_2[727:720]};
      mid_2[2] = {1'b0,layer_2_2[735:728]} - {1'b0, layer_1_2[735:728]};
      btm_0[0] = {1'b0,layer_3_0[719:712]} - {1'b0, layer_2_0[719:712]};
      btm_0[1] = {1'b0,layer_3_0[727:720]} - {1'b0, layer_2_0[727:720]};
      btm_0[2] = {1'b0,layer_3_0[735:728]} - {1'b0, layer_2_0[735:728]};
      btm_1[0] = {1'b0,layer_3_1[719:712]} - {1'b0, layer_2_1[719:712]};
      btm_1[1] = {1'b0,layer_3_1[727:720]} - {1'b0, layer_2_1[727:720]};
      btm_1[2] = {1'b0,layer_3_1[735:728]} - {1'b0, layer_2_1[735:728]};
      btm_2[0] = {1'b0,layer_3_2[719:712]} - {1'b0, layer_2_2[719:712]};
      btm_2[1] = {1'b0,layer_3_2[727:720]} - {1'b0, layer_2_2[727:720]};
      btm_2[2] = {1'b0,layer_3_2[735:728]} - {1'b0, layer_2_2[735:728]};
    end
    'd91: begin
      top_0[0] = {1'b0,layer_1_0[727:720]} - {1'b0, layer_0_0[727:720]};
      top_0[1] = {1'b0,layer_1_0[735:728]} - {1'b0, layer_0_0[735:728]};
      top_0[2] = {1'b0,layer_1_0[743:736]} - {1'b0, layer_0_0[743:736]};
      top_1[0] = {1'b0,layer_1_1[727:720]} - {1'b0, layer_0_1[727:720]};
      top_1[1] = {1'b0,layer_1_1[735:728]} - {1'b0, layer_0_1[735:728]};
      top_1[2] = {1'b0,layer_1_1[743:736]} - {1'b0, layer_0_1[743:736]};
      top_2[0] = {1'b0,layer_1_2[727:720]} - {1'b0, layer_0_2[727:720]};
      top_2[1] = {1'b0,layer_1_2[735:728]} - {1'b0, layer_0_2[735:728]};
      top_2[2] = {1'b0,layer_1_2[743:736]} - {1'b0, layer_0_2[743:736]};
      mid_0[0] = {1'b0,layer_2_0[727:720]} - {1'b0, layer_1_0[727:720]};
      mid_0[1] = {1'b0,layer_2_0[735:728]} - {1'b0, layer_1_0[735:728]};
      mid_0[2] = {1'b0,layer_2_0[743:736]} - {1'b0, layer_1_0[743:736]};
      mid_1[0] = {1'b0,layer_2_1[727:720]} - {1'b0, layer_1_1[727:720]};
      mid_1[1] = {1'b0,layer_2_1[735:728]} - {1'b0, layer_1_1[735:728]};
      mid_1[2] = {1'b0,layer_2_1[743:736]} - {1'b0, layer_1_1[743:736]};
      mid_2[0] = {1'b0,layer_2_2[727:720]} - {1'b0, layer_1_2[727:720]};
      mid_2[1] = {1'b0,layer_2_2[735:728]} - {1'b0, layer_1_2[735:728]};
      mid_2[2] = {1'b0,layer_2_2[743:736]} - {1'b0, layer_1_2[743:736]};
      btm_0[0] = {1'b0,layer_3_0[727:720]} - {1'b0, layer_2_0[727:720]};
      btm_0[1] = {1'b0,layer_3_0[735:728]} - {1'b0, layer_2_0[735:728]};
      btm_0[2] = {1'b0,layer_3_0[743:736]} - {1'b0, layer_2_0[743:736]};
      btm_1[0] = {1'b0,layer_3_1[727:720]} - {1'b0, layer_2_1[727:720]};
      btm_1[1] = {1'b0,layer_3_1[735:728]} - {1'b0, layer_2_1[735:728]};
      btm_1[2] = {1'b0,layer_3_1[743:736]} - {1'b0, layer_2_1[743:736]};
      btm_2[0] = {1'b0,layer_3_2[727:720]} - {1'b0, layer_2_2[727:720]};
      btm_2[1] = {1'b0,layer_3_2[735:728]} - {1'b0, layer_2_2[735:728]};
      btm_2[2] = {1'b0,layer_3_2[743:736]} - {1'b0, layer_2_2[743:736]};
    end
    'd92: begin
      top_0[0] = {1'b0,layer_1_0[735:728]} - {1'b0, layer_0_0[735:728]};
      top_0[1] = {1'b0,layer_1_0[743:736]} - {1'b0, layer_0_0[743:736]};
      top_0[2] = {1'b0,layer_1_0[751:744]} - {1'b0, layer_0_0[751:744]};
      top_1[0] = {1'b0,layer_1_1[735:728]} - {1'b0, layer_0_1[735:728]};
      top_1[1] = {1'b0,layer_1_1[743:736]} - {1'b0, layer_0_1[743:736]};
      top_1[2] = {1'b0,layer_1_1[751:744]} - {1'b0, layer_0_1[751:744]};
      top_2[0] = {1'b0,layer_1_2[735:728]} - {1'b0, layer_0_2[735:728]};
      top_2[1] = {1'b0,layer_1_2[743:736]} - {1'b0, layer_0_2[743:736]};
      top_2[2] = {1'b0,layer_1_2[751:744]} - {1'b0, layer_0_2[751:744]};
      mid_0[0] = {1'b0,layer_2_0[735:728]} - {1'b0, layer_1_0[735:728]};
      mid_0[1] = {1'b0,layer_2_0[743:736]} - {1'b0, layer_1_0[743:736]};
      mid_0[2] = {1'b0,layer_2_0[751:744]} - {1'b0, layer_1_0[751:744]};
      mid_1[0] = {1'b0,layer_2_1[735:728]} - {1'b0, layer_1_1[735:728]};
      mid_1[1] = {1'b0,layer_2_1[743:736]} - {1'b0, layer_1_1[743:736]};
      mid_1[2] = {1'b0,layer_2_1[751:744]} - {1'b0, layer_1_1[751:744]};
      mid_2[0] = {1'b0,layer_2_2[735:728]} - {1'b0, layer_1_2[735:728]};
      mid_2[1] = {1'b0,layer_2_2[743:736]} - {1'b0, layer_1_2[743:736]};
      mid_2[2] = {1'b0,layer_2_2[751:744]} - {1'b0, layer_1_2[751:744]};
      btm_0[0] = {1'b0,layer_3_0[735:728]} - {1'b0, layer_2_0[735:728]};
      btm_0[1] = {1'b0,layer_3_0[743:736]} - {1'b0, layer_2_0[743:736]};
      btm_0[2] = {1'b0,layer_3_0[751:744]} - {1'b0, layer_2_0[751:744]};
      btm_1[0] = {1'b0,layer_3_1[735:728]} - {1'b0, layer_2_1[735:728]};
      btm_1[1] = {1'b0,layer_3_1[743:736]} - {1'b0, layer_2_1[743:736]};
      btm_1[2] = {1'b0,layer_3_1[751:744]} - {1'b0, layer_2_1[751:744]};
      btm_2[0] = {1'b0,layer_3_2[735:728]} - {1'b0, layer_2_2[735:728]};
      btm_2[1] = {1'b0,layer_3_2[743:736]} - {1'b0, layer_2_2[743:736]};
      btm_2[2] = {1'b0,layer_3_2[751:744]} - {1'b0, layer_2_2[751:744]};
    end
    'd93: begin
      top_0[0] = {1'b0,layer_1_0[743:736]} - {1'b0, layer_0_0[743:736]};
      top_0[1] = {1'b0,layer_1_0[751:744]} - {1'b0, layer_0_0[751:744]};
      top_0[2] = {1'b0,layer_1_0[759:752]} - {1'b0, layer_0_0[759:752]};
      top_1[0] = {1'b0,layer_1_1[743:736]} - {1'b0, layer_0_1[743:736]};
      top_1[1] = {1'b0,layer_1_1[751:744]} - {1'b0, layer_0_1[751:744]};
      top_1[2] = {1'b0,layer_1_1[759:752]} - {1'b0, layer_0_1[759:752]};
      top_2[0] = {1'b0,layer_1_2[743:736]} - {1'b0, layer_0_2[743:736]};
      top_2[1] = {1'b0,layer_1_2[751:744]} - {1'b0, layer_0_2[751:744]};
      top_2[2] = {1'b0,layer_1_2[759:752]} - {1'b0, layer_0_2[759:752]};
      mid_0[0] = {1'b0,layer_2_0[743:736]} - {1'b0, layer_1_0[743:736]};
      mid_0[1] = {1'b0,layer_2_0[751:744]} - {1'b0, layer_1_0[751:744]};
      mid_0[2] = {1'b0,layer_2_0[759:752]} - {1'b0, layer_1_0[759:752]};
      mid_1[0] = {1'b0,layer_2_1[743:736]} - {1'b0, layer_1_1[743:736]};
      mid_1[1] = {1'b0,layer_2_1[751:744]} - {1'b0, layer_1_1[751:744]};
      mid_1[2] = {1'b0,layer_2_1[759:752]} - {1'b0, layer_1_1[759:752]};
      mid_2[0] = {1'b0,layer_2_2[743:736]} - {1'b0, layer_1_2[743:736]};
      mid_2[1] = {1'b0,layer_2_2[751:744]} - {1'b0, layer_1_2[751:744]};
      mid_2[2] = {1'b0,layer_2_2[759:752]} - {1'b0, layer_1_2[759:752]};
      btm_0[0] = {1'b0,layer_3_0[743:736]} - {1'b0, layer_2_0[743:736]};
      btm_0[1] = {1'b0,layer_3_0[751:744]} - {1'b0, layer_2_0[751:744]};
      btm_0[2] = {1'b0,layer_3_0[759:752]} - {1'b0, layer_2_0[759:752]};
      btm_1[0] = {1'b0,layer_3_1[743:736]} - {1'b0, layer_2_1[743:736]};
      btm_1[1] = {1'b0,layer_3_1[751:744]} - {1'b0, layer_2_1[751:744]};
      btm_1[2] = {1'b0,layer_3_1[759:752]} - {1'b0, layer_2_1[759:752]};
      btm_2[0] = {1'b0,layer_3_2[743:736]} - {1'b0, layer_2_2[743:736]};
      btm_2[1] = {1'b0,layer_3_2[751:744]} - {1'b0, layer_2_2[751:744]};
      btm_2[2] = {1'b0,layer_3_2[759:752]} - {1'b0, layer_2_2[759:752]};
    end
    'd94: begin
      top_0[0] = {1'b0,layer_1_0[751:744]} - {1'b0, layer_0_0[751:744]};
      top_0[1] = {1'b0,layer_1_0[759:752]} - {1'b0, layer_0_0[759:752]};
      top_0[2] = {1'b0,layer_1_0[767:760]} - {1'b0, layer_0_0[767:760]};
      top_1[0] = {1'b0,layer_1_1[751:744]} - {1'b0, layer_0_1[751:744]};
      top_1[1] = {1'b0,layer_1_1[759:752]} - {1'b0, layer_0_1[759:752]};
      top_1[2] = {1'b0,layer_1_1[767:760]} - {1'b0, layer_0_1[767:760]};
      top_2[0] = {1'b0,layer_1_2[751:744]} - {1'b0, layer_0_2[751:744]};
      top_2[1] = {1'b0,layer_1_2[759:752]} - {1'b0, layer_0_2[759:752]};
      top_2[2] = {1'b0,layer_1_2[767:760]} - {1'b0, layer_0_2[767:760]};
      mid_0[0] = {1'b0,layer_2_0[751:744]} - {1'b0, layer_1_0[751:744]};
      mid_0[1] = {1'b0,layer_2_0[759:752]} - {1'b0, layer_1_0[759:752]};
      mid_0[2] = {1'b0,layer_2_0[767:760]} - {1'b0, layer_1_0[767:760]};
      mid_1[0] = {1'b0,layer_2_1[751:744]} - {1'b0, layer_1_1[751:744]};
      mid_1[1] = {1'b0,layer_2_1[759:752]} - {1'b0, layer_1_1[759:752]};
      mid_1[2] = {1'b0,layer_2_1[767:760]} - {1'b0, layer_1_1[767:760]};
      mid_2[0] = {1'b0,layer_2_2[751:744]} - {1'b0, layer_1_2[751:744]};
      mid_2[1] = {1'b0,layer_2_2[759:752]} - {1'b0, layer_1_2[759:752]};
      mid_2[2] = {1'b0,layer_2_2[767:760]} - {1'b0, layer_1_2[767:760]};
      btm_0[0] = {1'b0,layer_3_0[751:744]} - {1'b0, layer_2_0[751:744]};
      btm_0[1] = {1'b0,layer_3_0[759:752]} - {1'b0, layer_2_0[759:752]};
      btm_0[2] = {1'b0,layer_3_0[767:760]} - {1'b0, layer_2_0[767:760]};
      btm_1[0] = {1'b0,layer_3_1[751:744]} - {1'b0, layer_2_1[751:744]};
      btm_1[1] = {1'b0,layer_3_1[759:752]} - {1'b0, layer_2_1[759:752]};
      btm_1[2] = {1'b0,layer_3_1[767:760]} - {1'b0, layer_2_1[767:760]};
      btm_2[0] = {1'b0,layer_3_2[751:744]} - {1'b0, layer_2_2[751:744]};
      btm_2[1] = {1'b0,layer_3_2[759:752]} - {1'b0, layer_2_2[759:752]};
      btm_2[2] = {1'b0,layer_3_2[767:760]} - {1'b0, layer_2_2[767:760]};
    end
    'd95: begin
      top_0[0] = {1'b0,layer_1_0[759:752]} - {1'b0, layer_0_0[759:752]};
      top_0[1] = {1'b0,layer_1_0[767:760]} - {1'b0, layer_0_0[767:760]};
      top_0[2] = {1'b0,layer_1_0[775:768]} - {1'b0, layer_0_0[775:768]};
      top_1[0] = {1'b0,layer_1_1[759:752]} - {1'b0, layer_0_1[759:752]};
      top_1[1] = {1'b0,layer_1_1[767:760]} - {1'b0, layer_0_1[767:760]};
      top_1[2] = {1'b0,layer_1_1[775:768]} - {1'b0, layer_0_1[775:768]};
      top_2[0] = {1'b0,layer_1_2[759:752]} - {1'b0, layer_0_2[759:752]};
      top_2[1] = {1'b0,layer_1_2[767:760]} - {1'b0, layer_0_2[767:760]};
      top_2[2] = {1'b0,layer_1_2[775:768]} - {1'b0, layer_0_2[775:768]};
      mid_0[0] = {1'b0,layer_2_0[759:752]} - {1'b0, layer_1_0[759:752]};
      mid_0[1] = {1'b0,layer_2_0[767:760]} - {1'b0, layer_1_0[767:760]};
      mid_0[2] = {1'b0,layer_2_0[775:768]} - {1'b0, layer_1_0[775:768]};
      mid_1[0] = {1'b0,layer_2_1[759:752]} - {1'b0, layer_1_1[759:752]};
      mid_1[1] = {1'b0,layer_2_1[767:760]} - {1'b0, layer_1_1[767:760]};
      mid_1[2] = {1'b0,layer_2_1[775:768]} - {1'b0, layer_1_1[775:768]};
      mid_2[0] = {1'b0,layer_2_2[759:752]} - {1'b0, layer_1_2[759:752]};
      mid_2[1] = {1'b0,layer_2_2[767:760]} - {1'b0, layer_1_2[767:760]};
      mid_2[2] = {1'b0,layer_2_2[775:768]} - {1'b0, layer_1_2[775:768]};
      btm_0[0] = {1'b0,layer_3_0[759:752]} - {1'b0, layer_2_0[759:752]};
      btm_0[1] = {1'b0,layer_3_0[767:760]} - {1'b0, layer_2_0[767:760]};
      btm_0[2] = {1'b0,layer_3_0[775:768]} - {1'b0, layer_2_0[775:768]};
      btm_1[0] = {1'b0,layer_3_1[759:752]} - {1'b0, layer_2_1[759:752]};
      btm_1[1] = {1'b0,layer_3_1[767:760]} - {1'b0, layer_2_1[767:760]};
      btm_1[2] = {1'b0,layer_3_1[775:768]} - {1'b0, layer_2_1[775:768]};
      btm_2[0] = {1'b0,layer_3_2[759:752]} - {1'b0, layer_2_2[759:752]};
      btm_2[1] = {1'b0,layer_3_2[767:760]} - {1'b0, layer_2_2[767:760]};
      btm_2[2] = {1'b0,layer_3_2[775:768]} - {1'b0, layer_2_2[775:768]};
    end
    'd96: begin
      top_0[0] = {1'b0,layer_1_0[767:760]} - {1'b0, layer_0_0[767:760]};
      top_0[1] = {1'b0,layer_1_0[775:768]} - {1'b0, layer_0_0[775:768]};
      top_0[2] = {1'b0,layer_1_0[783:776]} - {1'b0, layer_0_0[783:776]};
      top_1[0] = {1'b0,layer_1_1[767:760]} - {1'b0, layer_0_1[767:760]};
      top_1[1] = {1'b0,layer_1_1[775:768]} - {1'b0, layer_0_1[775:768]};
      top_1[2] = {1'b0,layer_1_1[783:776]} - {1'b0, layer_0_1[783:776]};
      top_2[0] = {1'b0,layer_1_2[767:760]} - {1'b0, layer_0_2[767:760]};
      top_2[1] = {1'b0,layer_1_2[775:768]} - {1'b0, layer_0_2[775:768]};
      top_2[2] = {1'b0,layer_1_2[783:776]} - {1'b0, layer_0_2[783:776]};
      mid_0[0] = {1'b0,layer_2_0[767:760]} - {1'b0, layer_1_0[767:760]};
      mid_0[1] = {1'b0,layer_2_0[775:768]} - {1'b0, layer_1_0[775:768]};
      mid_0[2] = {1'b0,layer_2_0[783:776]} - {1'b0, layer_1_0[783:776]};
      mid_1[0] = {1'b0,layer_2_1[767:760]} - {1'b0, layer_1_1[767:760]};
      mid_1[1] = {1'b0,layer_2_1[775:768]} - {1'b0, layer_1_1[775:768]};
      mid_1[2] = {1'b0,layer_2_1[783:776]} - {1'b0, layer_1_1[783:776]};
      mid_2[0] = {1'b0,layer_2_2[767:760]} - {1'b0, layer_1_2[767:760]};
      mid_2[1] = {1'b0,layer_2_2[775:768]} - {1'b0, layer_1_2[775:768]};
      mid_2[2] = {1'b0,layer_2_2[783:776]} - {1'b0, layer_1_2[783:776]};
      btm_0[0] = {1'b0,layer_3_0[767:760]} - {1'b0, layer_2_0[767:760]};
      btm_0[1] = {1'b0,layer_3_0[775:768]} - {1'b0, layer_2_0[775:768]};
      btm_0[2] = {1'b0,layer_3_0[783:776]} - {1'b0, layer_2_0[783:776]};
      btm_1[0] = {1'b0,layer_3_1[767:760]} - {1'b0, layer_2_1[767:760]};
      btm_1[1] = {1'b0,layer_3_1[775:768]} - {1'b0, layer_2_1[775:768]};
      btm_1[2] = {1'b0,layer_3_1[783:776]} - {1'b0, layer_2_1[783:776]};
      btm_2[0] = {1'b0,layer_3_2[767:760]} - {1'b0, layer_2_2[767:760]};
      btm_2[1] = {1'b0,layer_3_2[775:768]} - {1'b0, layer_2_2[775:768]};
      btm_2[2] = {1'b0,layer_3_2[783:776]} - {1'b0, layer_2_2[783:776]};
    end
    'd97: begin
      top_0[0] = {1'b0,layer_1_0[775:768]} - {1'b0, layer_0_0[775:768]};
      top_0[1] = {1'b0,layer_1_0[783:776]} - {1'b0, layer_0_0[783:776]};
      top_0[2] = {1'b0,layer_1_0[791:784]} - {1'b0, layer_0_0[791:784]};
      top_1[0] = {1'b0,layer_1_1[775:768]} - {1'b0, layer_0_1[775:768]};
      top_1[1] = {1'b0,layer_1_1[783:776]} - {1'b0, layer_0_1[783:776]};
      top_1[2] = {1'b0,layer_1_1[791:784]} - {1'b0, layer_0_1[791:784]};
      top_2[0] = {1'b0,layer_1_2[775:768]} - {1'b0, layer_0_2[775:768]};
      top_2[1] = {1'b0,layer_1_2[783:776]} - {1'b0, layer_0_2[783:776]};
      top_2[2] = {1'b0,layer_1_2[791:784]} - {1'b0, layer_0_2[791:784]};
      mid_0[0] = {1'b0,layer_2_0[775:768]} - {1'b0, layer_1_0[775:768]};
      mid_0[1] = {1'b0,layer_2_0[783:776]} - {1'b0, layer_1_0[783:776]};
      mid_0[2] = {1'b0,layer_2_0[791:784]} - {1'b0, layer_1_0[791:784]};
      mid_1[0] = {1'b0,layer_2_1[775:768]} - {1'b0, layer_1_1[775:768]};
      mid_1[1] = {1'b0,layer_2_1[783:776]} - {1'b0, layer_1_1[783:776]};
      mid_1[2] = {1'b0,layer_2_1[791:784]} - {1'b0, layer_1_1[791:784]};
      mid_2[0] = {1'b0,layer_2_2[775:768]} - {1'b0, layer_1_2[775:768]};
      mid_2[1] = {1'b0,layer_2_2[783:776]} - {1'b0, layer_1_2[783:776]};
      mid_2[2] = {1'b0,layer_2_2[791:784]} - {1'b0, layer_1_2[791:784]};
      btm_0[0] = {1'b0,layer_3_0[775:768]} - {1'b0, layer_2_0[775:768]};
      btm_0[1] = {1'b0,layer_3_0[783:776]} - {1'b0, layer_2_0[783:776]};
      btm_0[2] = {1'b0,layer_3_0[791:784]} - {1'b0, layer_2_0[791:784]};
      btm_1[0] = {1'b0,layer_3_1[775:768]} - {1'b0, layer_2_1[775:768]};
      btm_1[1] = {1'b0,layer_3_1[783:776]} - {1'b0, layer_2_1[783:776]};
      btm_1[2] = {1'b0,layer_3_1[791:784]} - {1'b0, layer_2_1[791:784]};
      btm_2[0] = {1'b0,layer_3_2[775:768]} - {1'b0, layer_2_2[775:768]};
      btm_2[1] = {1'b0,layer_3_2[783:776]} - {1'b0, layer_2_2[783:776]};
      btm_2[2] = {1'b0,layer_3_2[791:784]} - {1'b0, layer_2_2[791:784]};
    end
    'd98: begin
      top_0[0] = {1'b0,layer_1_0[783:776]} - {1'b0, layer_0_0[783:776]};
      top_0[1] = {1'b0,layer_1_0[791:784]} - {1'b0, layer_0_0[791:784]};
      top_0[2] = {1'b0,layer_1_0[799:792]} - {1'b0, layer_0_0[799:792]};
      top_1[0] = {1'b0,layer_1_1[783:776]} - {1'b0, layer_0_1[783:776]};
      top_1[1] = {1'b0,layer_1_1[791:784]} - {1'b0, layer_0_1[791:784]};
      top_1[2] = {1'b0,layer_1_1[799:792]} - {1'b0, layer_0_1[799:792]};
      top_2[0] = {1'b0,layer_1_2[783:776]} - {1'b0, layer_0_2[783:776]};
      top_2[1] = {1'b0,layer_1_2[791:784]} - {1'b0, layer_0_2[791:784]};
      top_2[2] = {1'b0,layer_1_2[799:792]} - {1'b0, layer_0_2[799:792]};
      mid_0[0] = {1'b0,layer_2_0[783:776]} - {1'b0, layer_1_0[783:776]};
      mid_0[1] = {1'b0,layer_2_0[791:784]} - {1'b0, layer_1_0[791:784]};
      mid_0[2] = {1'b0,layer_2_0[799:792]} - {1'b0, layer_1_0[799:792]};
      mid_1[0] = {1'b0,layer_2_1[783:776]} - {1'b0, layer_1_1[783:776]};
      mid_1[1] = {1'b0,layer_2_1[791:784]} - {1'b0, layer_1_1[791:784]};
      mid_1[2] = {1'b0,layer_2_1[799:792]} - {1'b0, layer_1_1[799:792]};
      mid_2[0] = {1'b0,layer_2_2[783:776]} - {1'b0, layer_1_2[783:776]};
      mid_2[1] = {1'b0,layer_2_2[791:784]} - {1'b0, layer_1_2[791:784]};
      mid_2[2] = {1'b0,layer_2_2[799:792]} - {1'b0, layer_1_2[799:792]};
      btm_0[0] = {1'b0,layer_3_0[783:776]} - {1'b0, layer_2_0[783:776]};
      btm_0[1] = {1'b0,layer_3_0[791:784]} - {1'b0, layer_2_0[791:784]};
      btm_0[2] = {1'b0,layer_3_0[799:792]} - {1'b0, layer_2_0[799:792]};
      btm_1[0] = {1'b0,layer_3_1[783:776]} - {1'b0, layer_2_1[783:776]};
      btm_1[1] = {1'b0,layer_3_1[791:784]} - {1'b0, layer_2_1[791:784]};
      btm_1[2] = {1'b0,layer_3_1[799:792]} - {1'b0, layer_2_1[799:792]};
      btm_2[0] = {1'b0,layer_3_2[783:776]} - {1'b0, layer_2_2[783:776]};
      btm_2[1] = {1'b0,layer_3_2[791:784]} - {1'b0, layer_2_2[791:784]};
      btm_2[2] = {1'b0,layer_3_2[799:792]} - {1'b0, layer_2_2[799:792]};
    end
    'd99: begin
      top_0[0] = {1'b0,layer_1_0[791:784]} - {1'b0, layer_0_0[791:784]};
      top_0[1] = {1'b0,layer_1_0[799:792]} - {1'b0, layer_0_0[799:792]};
      top_0[2] = {1'b0,layer_1_0[807:800]} - {1'b0, layer_0_0[807:800]};
      top_1[0] = {1'b0,layer_1_1[791:784]} - {1'b0, layer_0_1[791:784]};
      top_1[1] = {1'b0,layer_1_1[799:792]} - {1'b0, layer_0_1[799:792]};
      top_1[2] = {1'b0,layer_1_1[807:800]} - {1'b0, layer_0_1[807:800]};
      top_2[0] = {1'b0,layer_1_2[791:784]} - {1'b0, layer_0_2[791:784]};
      top_2[1] = {1'b0,layer_1_2[799:792]} - {1'b0, layer_0_2[799:792]};
      top_2[2] = {1'b0,layer_1_2[807:800]} - {1'b0, layer_0_2[807:800]};
      mid_0[0] = {1'b0,layer_2_0[791:784]} - {1'b0, layer_1_0[791:784]};
      mid_0[1] = {1'b0,layer_2_0[799:792]} - {1'b0, layer_1_0[799:792]};
      mid_0[2] = {1'b0,layer_2_0[807:800]} - {1'b0, layer_1_0[807:800]};
      mid_1[0] = {1'b0,layer_2_1[791:784]} - {1'b0, layer_1_1[791:784]};
      mid_1[1] = {1'b0,layer_2_1[799:792]} - {1'b0, layer_1_1[799:792]};
      mid_1[2] = {1'b0,layer_2_1[807:800]} - {1'b0, layer_1_1[807:800]};
      mid_2[0] = {1'b0,layer_2_2[791:784]} - {1'b0, layer_1_2[791:784]};
      mid_2[1] = {1'b0,layer_2_2[799:792]} - {1'b0, layer_1_2[799:792]};
      mid_2[2] = {1'b0,layer_2_2[807:800]} - {1'b0, layer_1_2[807:800]};
      btm_0[0] = {1'b0,layer_3_0[791:784]} - {1'b0, layer_2_0[791:784]};
      btm_0[1] = {1'b0,layer_3_0[799:792]} - {1'b0, layer_2_0[799:792]};
      btm_0[2] = {1'b0,layer_3_0[807:800]} - {1'b0, layer_2_0[807:800]};
      btm_1[0] = {1'b0,layer_3_1[791:784]} - {1'b0, layer_2_1[791:784]};
      btm_1[1] = {1'b0,layer_3_1[799:792]} - {1'b0, layer_2_1[799:792]};
      btm_1[2] = {1'b0,layer_3_1[807:800]} - {1'b0, layer_2_1[807:800]};
      btm_2[0] = {1'b0,layer_3_2[791:784]} - {1'b0, layer_2_2[791:784]};
      btm_2[1] = {1'b0,layer_3_2[799:792]} - {1'b0, layer_2_2[799:792]};
      btm_2[2] = {1'b0,layer_3_2[807:800]} - {1'b0, layer_2_2[807:800]};
    end
    'd100: begin
      top_0[0] = {1'b0,layer_1_0[799:792]} - {1'b0, layer_0_0[799:792]};
      top_0[1] = {1'b0,layer_1_0[807:800]} - {1'b0, layer_0_0[807:800]};
      top_0[2] = {1'b0,layer_1_0[815:808]} - {1'b0, layer_0_0[815:808]};
      top_1[0] = {1'b0,layer_1_1[799:792]} - {1'b0, layer_0_1[799:792]};
      top_1[1] = {1'b0,layer_1_1[807:800]} - {1'b0, layer_0_1[807:800]};
      top_1[2] = {1'b0,layer_1_1[815:808]} - {1'b0, layer_0_1[815:808]};
      top_2[0] = {1'b0,layer_1_2[799:792]} - {1'b0, layer_0_2[799:792]};
      top_2[1] = {1'b0,layer_1_2[807:800]} - {1'b0, layer_0_2[807:800]};
      top_2[2] = {1'b0,layer_1_2[815:808]} - {1'b0, layer_0_2[815:808]};
      mid_0[0] = {1'b0,layer_2_0[799:792]} - {1'b0, layer_1_0[799:792]};
      mid_0[1] = {1'b0,layer_2_0[807:800]} - {1'b0, layer_1_0[807:800]};
      mid_0[2] = {1'b0,layer_2_0[815:808]} - {1'b0, layer_1_0[815:808]};
      mid_1[0] = {1'b0,layer_2_1[799:792]} - {1'b0, layer_1_1[799:792]};
      mid_1[1] = {1'b0,layer_2_1[807:800]} - {1'b0, layer_1_1[807:800]};
      mid_1[2] = {1'b0,layer_2_1[815:808]} - {1'b0, layer_1_1[815:808]};
      mid_2[0] = {1'b0,layer_2_2[799:792]} - {1'b0, layer_1_2[799:792]};
      mid_2[1] = {1'b0,layer_2_2[807:800]} - {1'b0, layer_1_2[807:800]};
      mid_2[2] = {1'b0,layer_2_2[815:808]} - {1'b0, layer_1_2[815:808]};
      btm_0[0] = {1'b0,layer_3_0[799:792]} - {1'b0, layer_2_0[799:792]};
      btm_0[1] = {1'b0,layer_3_0[807:800]} - {1'b0, layer_2_0[807:800]};
      btm_0[2] = {1'b0,layer_3_0[815:808]} - {1'b0, layer_2_0[815:808]};
      btm_1[0] = {1'b0,layer_3_1[799:792]} - {1'b0, layer_2_1[799:792]};
      btm_1[1] = {1'b0,layer_3_1[807:800]} - {1'b0, layer_2_1[807:800]};
      btm_1[2] = {1'b0,layer_3_1[815:808]} - {1'b0, layer_2_1[815:808]};
      btm_2[0] = {1'b0,layer_3_2[799:792]} - {1'b0, layer_2_2[799:792]};
      btm_2[1] = {1'b0,layer_3_2[807:800]} - {1'b0, layer_2_2[807:800]};
      btm_2[2] = {1'b0,layer_3_2[815:808]} - {1'b0, layer_2_2[815:808]};
    end
    'd101: begin
      top_0[0] = {1'b0,layer_1_0[807:800]} - {1'b0, layer_0_0[807:800]};
      top_0[1] = {1'b0,layer_1_0[815:808]} - {1'b0, layer_0_0[815:808]};
      top_0[2] = {1'b0,layer_1_0[823:816]} - {1'b0, layer_0_0[823:816]};
      top_1[0] = {1'b0,layer_1_1[807:800]} - {1'b0, layer_0_1[807:800]};
      top_1[1] = {1'b0,layer_1_1[815:808]} - {1'b0, layer_0_1[815:808]};
      top_1[2] = {1'b0,layer_1_1[823:816]} - {1'b0, layer_0_1[823:816]};
      top_2[0] = {1'b0,layer_1_2[807:800]} - {1'b0, layer_0_2[807:800]};
      top_2[1] = {1'b0,layer_1_2[815:808]} - {1'b0, layer_0_2[815:808]};
      top_2[2] = {1'b0,layer_1_2[823:816]} - {1'b0, layer_0_2[823:816]};
      mid_0[0] = {1'b0,layer_2_0[807:800]} - {1'b0, layer_1_0[807:800]};
      mid_0[1] = {1'b0,layer_2_0[815:808]} - {1'b0, layer_1_0[815:808]};
      mid_0[2] = {1'b0,layer_2_0[823:816]} - {1'b0, layer_1_0[823:816]};
      mid_1[0] = {1'b0,layer_2_1[807:800]} - {1'b0, layer_1_1[807:800]};
      mid_1[1] = {1'b0,layer_2_1[815:808]} - {1'b0, layer_1_1[815:808]};
      mid_1[2] = {1'b0,layer_2_1[823:816]} - {1'b0, layer_1_1[823:816]};
      mid_2[0] = {1'b0,layer_2_2[807:800]} - {1'b0, layer_1_2[807:800]};
      mid_2[1] = {1'b0,layer_2_2[815:808]} - {1'b0, layer_1_2[815:808]};
      mid_2[2] = {1'b0,layer_2_2[823:816]} - {1'b0, layer_1_2[823:816]};
      btm_0[0] = {1'b0,layer_3_0[807:800]} - {1'b0, layer_2_0[807:800]};
      btm_0[1] = {1'b0,layer_3_0[815:808]} - {1'b0, layer_2_0[815:808]};
      btm_0[2] = {1'b0,layer_3_0[823:816]} - {1'b0, layer_2_0[823:816]};
      btm_1[0] = {1'b0,layer_3_1[807:800]} - {1'b0, layer_2_1[807:800]};
      btm_1[1] = {1'b0,layer_3_1[815:808]} - {1'b0, layer_2_1[815:808]};
      btm_1[2] = {1'b0,layer_3_1[823:816]} - {1'b0, layer_2_1[823:816]};
      btm_2[0] = {1'b0,layer_3_2[807:800]} - {1'b0, layer_2_2[807:800]};
      btm_2[1] = {1'b0,layer_3_2[815:808]} - {1'b0, layer_2_2[815:808]};
      btm_2[2] = {1'b0,layer_3_2[823:816]} - {1'b0, layer_2_2[823:816]};
    end
    'd102: begin
      top_0[0] = {1'b0,layer_1_0[815:808]} - {1'b0, layer_0_0[815:808]};
      top_0[1] = {1'b0,layer_1_0[823:816]} - {1'b0, layer_0_0[823:816]};
      top_0[2] = {1'b0,layer_1_0[831:824]} - {1'b0, layer_0_0[831:824]};
      top_1[0] = {1'b0,layer_1_1[815:808]} - {1'b0, layer_0_1[815:808]};
      top_1[1] = {1'b0,layer_1_1[823:816]} - {1'b0, layer_0_1[823:816]};
      top_1[2] = {1'b0,layer_1_1[831:824]} - {1'b0, layer_0_1[831:824]};
      top_2[0] = {1'b0,layer_1_2[815:808]} - {1'b0, layer_0_2[815:808]};
      top_2[1] = {1'b0,layer_1_2[823:816]} - {1'b0, layer_0_2[823:816]};
      top_2[2] = {1'b0,layer_1_2[831:824]} - {1'b0, layer_0_2[831:824]};
      mid_0[0] = {1'b0,layer_2_0[815:808]} - {1'b0, layer_1_0[815:808]};
      mid_0[1] = {1'b0,layer_2_0[823:816]} - {1'b0, layer_1_0[823:816]};
      mid_0[2] = {1'b0,layer_2_0[831:824]} - {1'b0, layer_1_0[831:824]};
      mid_1[0] = {1'b0,layer_2_1[815:808]} - {1'b0, layer_1_1[815:808]};
      mid_1[1] = {1'b0,layer_2_1[823:816]} - {1'b0, layer_1_1[823:816]};
      mid_1[2] = {1'b0,layer_2_1[831:824]} - {1'b0, layer_1_1[831:824]};
      mid_2[0] = {1'b0,layer_2_2[815:808]} - {1'b0, layer_1_2[815:808]};
      mid_2[1] = {1'b0,layer_2_2[823:816]} - {1'b0, layer_1_2[823:816]};
      mid_2[2] = {1'b0,layer_2_2[831:824]} - {1'b0, layer_1_2[831:824]};
      btm_0[0] = {1'b0,layer_3_0[815:808]} - {1'b0, layer_2_0[815:808]};
      btm_0[1] = {1'b0,layer_3_0[823:816]} - {1'b0, layer_2_0[823:816]};
      btm_0[2] = {1'b0,layer_3_0[831:824]} - {1'b0, layer_2_0[831:824]};
      btm_1[0] = {1'b0,layer_3_1[815:808]} - {1'b0, layer_2_1[815:808]};
      btm_1[1] = {1'b0,layer_3_1[823:816]} - {1'b0, layer_2_1[823:816]};
      btm_1[2] = {1'b0,layer_3_1[831:824]} - {1'b0, layer_2_1[831:824]};
      btm_2[0] = {1'b0,layer_3_2[815:808]} - {1'b0, layer_2_2[815:808]};
      btm_2[1] = {1'b0,layer_3_2[823:816]} - {1'b0, layer_2_2[823:816]};
      btm_2[2] = {1'b0,layer_3_2[831:824]} - {1'b0, layer_2_2[831:824]};
    end
    'd103: begin
      top_0[0] = {1'b0,layer_1_0[823:816]} - {1'b0, layer_0_0[823:816]};
      top_0[1] = {1'b0,layer_1_0[831:824]} - {1'b0, layer_0_0[831:824]};
      top_0[2] = {1'b0,layer_1_0[839:832]} - {1'b0, layer_0_0[839:832]};
      top_1[0] = {1'b0,layer_1_1[823:816]} - {1'b0, layer_0_1[823:816]};
      top_1[1] = {1'b0,layer_1_1[831:824]} - {1'b0, layer_0_1[831:824]};
      top_1[2] = {1'b0,layer_1_1[839:832]} - {1'b0, layer_0_1[839:832]};
      top_2[0] = {1'b0,layer_1_2[823:816]} - {1'b0, layer_0_2[823:816]};
      top_2[1] = {1'b0,layer_1_2[831:824]} - {1'b0, layer_0_2[831:824]};
      top_2[2] = {1'b0,layer_1_2[839:832]} - {1'b0, layer_0_2[839:832]};
      mid_0[0] = {1'b0,layer_2_0[823:816]} - {1'b0, layer_1_0[823:816]};
      mid_0[1] = {1'b0,layer_2_0[831:824]} - {1'b0, layer_1_0[831:824]};
      mid_0[2] = {1'b0,layer_2_0[839:832]} - {1'b0, layer_1_0[839:832]};
      mid_1[0] = {1'b0,layer_2_1[823:816]} - {1'b0, layer_1_1[823:816]};
      mid_1[1] = {1'b0,layer_2_1[831:824]} - {1'b0, layer_1_1[831:824]};
      mid_1[2] = {1'b0,layer_2_1[839:832]} - {1'b0, layer_1_1[839:832]};
      mid_2[0] = {1'b0,layer_2_2[823:816]} - {1'b0, layer_1_2[823:816]};
      mid_2[1] = {1'b0,layer_2_2[831:824]} - {1'b0, layer_1_2[831:824]};
      mid_2[2] = {1'b0,layer_2_2[839:832]} - {1'b0, layer_1_2[839:832]};
      btm_0[0] = {1'b0,layer_3_0[823:816]} - {1'b0, layer_2_0[823:816]};
      btm_0[1] = {1'b0,layer_3_0[831:824]} - {1'b0, layer_2_0[831:824]};
      btm_0[2] = {1'b0,layer_3_0[839:832]} - {1'b0, layer_2_0[839:832]};
      btm_1[0] = {1'b0,layer_3_1[823:816]} - {1'b0, layer_2_1[823:816]};
      btm_1[1] = {1'b0,layer_3_1[831:824]} - {1'b0, layer_2_1[831:824]};
      btm_1[2] = {1'b0,layer_3_1[839:832]} - {1'b0, layer_2_1[839:832]};
      btm_2[0] = {1'b0,layer_3_2[823:816]} - {1'b0, layer_2_2[823:816]};
      btm_2[1] = {1'b0,layer_3_2[831:824]} - {1'b0, layer_2_2[831:824]};
      btm_2[2] = {1'b0,layer_3_2[839:832]} - {1'b0, layer_2_2[839:832]};
    end
    'd104: begin
      top_0[0] = {1'b0,layer_1_0[831:824]} - {1'b0, layer_0_0[831:824]};
      top_0[1] = {1'b0,layer_1_0[839:832]} - {1'b0, layer_0_0[839:832]};
      top_0[2] = {1'b0,layer_1_0[847:840]} - {1'b0, layer_0_0[847:840]};
      top_1[0] = {1'b0,layer_1_1[831:824]} - {1'b0, layer_0_1[831:824]};
      top_1[1] = {1'b0,layer_1_1[839:832]} - {1'b0, layer_0_1[839:832]};
      top_1[2] = {1'b0,layer_1_1[847:840]} - {1'b0, layer_0_1[847:840]};
      top_2[0] = {1'b0,layer_1_2[831:824]} - {1'b0, layer_0_2[831:824]};
      top_2[1] = {1'b0,layer_1_2[839:832]} - {1'b0, layer_0_2[839:832]};
      top_2[2] = {1'b0,layer_1_2[847:840]} - {1'b0, layer_0_2[847:840]};
      mid_0[0] = {1'b0,layer_2_0[831:824]} - {1'b0, layer_1_0[831:824]};
      mid_0[1] = {1'b0,layer_2_0[839:832]} - {1'b0, layer_1_0[839:832]};
      mid_0[2] = {1'b0,layer_2_0[847:840]} - {1'b0, layer_1_0[847:840]};
      mid_1[0] = {1'b0,layer_2_1[831:824]} - {1'b0, layer_1_1[831:824]};
      mid_1[1] = {1'b0,layer_2_1[839:832]} - {1'b0, layer_1_1[839:832]};
      mid_1[2] = {1'b0,layer_2_1[847:840]} - {1'b0, layer_1_1[847:840]};
      mid_2[0] = {1'b0,layer_2_2[831:824]} - {1'b0, layer_1_2[831:824]};
      mid_2[1] = {1'b0,layer_2_2[839:832]} - {1'b0, layer_1_2[839:832]};
      mid_2[2] = {1'b0,layer_2_2[847:840]} - {1'b0, layer_1_2[847:840]};
      btm_0[0] = {1'b0,layer_3_0[831:824]} - {1'b0, layer_2_0[831:824]};
      btm_0[1] = {1'b0,layer_3_0[839:832]} - {1'b0, layer_2_0[839:832]};
      btm_0[2] = {1'b0,layer_3_0[847:840]} - {1'b0, layer_2_0[847:840]};
      btm_1[0] = {1'b0,layer_3_1[831:824]} - {1'b0, layer_2_1[831:824]};
      btm_1[1] = {1'b0,layer_3_1[839:832]} - {1'b0, layer_2_1[839:832]};
      btm_1[2] = {1'b0,layer_3_1[847:840]} - {1'b0, layer_2_1[847:840]};
      btm_2[0] = {1'b0,layer_3_2[831:824]} - {1'b0, layer_2_2[831:824]};
      btm_2[1] = {1'b0,layer_3_2[839:832]} - {1'b0, layer_2_2[839:832]};
      btm_2[2] = {1'b0,layer_3_2[847:840]} - {1'b0, layer_2_2[847:840]};
    end
    'd105: begin
      top_0[0] = {1'b0,layer_1_0[839:832]} - {1'b0, layer_0_0[839:832]};
      top_0[1] = {1'b0,layer_1_0[847:840]} - {1'b0, layer_0_0[847:840]};
      top_0[2] = {1'b0,layer_1_0[855:848]} - {1'b0, layer_0_0[855:848]};
      top_1[0] = {1'b0,layer_1_1[839:832]} - {1'b0, layer_0_1[839:832]};
      top_1[1] = {1'b0,layer_1_1[847:840]} - {1'b0, layer_0_1[847:840]};
      top_1[2] = {1'b0,layer_1_1[855:848]} - {1'b0, layer_0_1[855:848]};
      top_2[0] = {1'b0,layer_1_2[839:832]} - {1'b0, layer_0_2[839:832]};
      top_2[1] = {1'b0,layer_1_2[847:840]} - {1'b0, layer_0_2[847:840]};
      top_2[2] = {1'b0,layer_1_2[855:848]} - {1'b0, layer_0_2[855:848]};
      mid_0[0] = {1'b0,layer_2_0[839:832]} - {1'b0, layer_1_0[839:832]};
      mid_0[1] = {1'b0,layer_2_0[847:840]} - {1'b0, layer_1_0[847:840]};
      mid_0[2] = {1'b0,layer_2_0[855:848]} - {1'b0, layer_1_0[855:848]};
      mid_1[0] = {1'b0,layer_2_1[839:832]} - {1'b0, layer_1_1[839:832]};
      mid_1[1] = {1'b0,layer_2_1[847:840]} - {1'b0, layer_1_1[847:840]};
      mid_1[2] = {1'b0,layer_2_1[855:848]} - {1'b0, layer_1_1[855:848]};
      mid_2[0] = {1'b0,layer_2_2[839:832]} - {1'b0, layer_1_2[839:832]};
      mid_2[1] = {1'b0,layer_2_2[847:840]} - {1'b0, layer_1_2[847:840]};
      mid_2[2] = {1'b0,layer_2_2[855:848]} - {1'b0, layer_1_2[855:848]};
      btm_0[0] = {1'b0,layer_3_0[839:832]} - {1'b0, layer_2_0[839:832]};
      btm_0[1] = {1'b0,layer_3_0[847:840]} - {1'b0, layer_2_0[847:840]};
      btm_0[2] = {1'b0,layer_3_0[855:848]} - {1'b0, layer_2_0[855:848]};
      btm_1[0] = {1'b0,layer_3_1[839:832]} - {1'b0, layer_2_1[839:832]};
      btm_1[1] = {1'b0,layer_3_1[847:840]} - {1'b0, layer_2_1[847:840]};
      btm_1[2] = {1'b0,layer_3_1[855:848]} - {1'b0, layer_2_1[855:848]};
      btm_2[0] = {1'b0,layer_3_2[839:832]} - {1'b0, layer_2_2[839:832]};
      btm_2[1] = {1'b0,layer_3_2[847:840]} - {1'b0, layer_2_2[847:840]};
      btm_2[2] = {1'b0,layer_3_2[855:848]} - {1'b0, layer_2_2[855:848]};
    end
    'd106: begin
      top_0[0] = {1'b0,layer_1_0[847:840]} - {1'b0, layer_0_0[847:840]};
      top_0[1] = {1'b0,layer_1_0[855:848]} - {1'b0, layer_0_0[855:848]};
      top_0[2] = {1'b0,layer_1_0[863:856]} - {1'b0, layer_0_0[863:856]};
      top_1[0] = {1'b0,layer_1_1[847:840]} - {1'b0, layer_0_1[847:840]};
      top_1[1] = {1'b0,layer_1_1[855:848]} - {1'b0, layer_0_1[855:848]};
      top_1[2] = {1'b0,layer_1_1[863:856]} - {1'b0, layer_0_1[863:856]};
      top_2[0] = {1'b0,layer_1_2[847:840]} - {1'b0, layer_0_2[847:840]};
      top_2[1] = {1'b0,layer_1_2[855:848]} - {1'b0, layer_0_2[855:848]};
      top_2[2] = {1'b0,layer_1_2[863:856]} - {1'b0, layer_0_2[863:856]};
      mid_0[0] = {1'b0,layer_2_0[847:840]} - {1'b0, layer_1_0[847:840]};
      mid_0[1] = {1'b0,layer_2_0[855:848]} - {1'b0, layer_1_0[855:848]};
      mid_0[2] = {1'b0,layer_2_0[863:856]} - {1'b0, layer_1_0[863:856]};
      mid_1[0] = {1'b0,layer_2_1[847:840]} - {1'b0, layer_1_1[847:840]};
      mid_1[1] = {1'b0,layer_2_1[855:848]} - {1'b0, layer_1_1[855:848]};
      mid_1[2] = {1'b0,layer_2_1[863:856]} - {1'b0, layer_1_1[863:856]};
      mid_2[0] = {1'b0,layer_2_2[847:840]} - {1'b0, layer_1_2[847:840]};
      mid_2[1] = {1'b0,layer_2_2[855:848]} - {1'b0, layer_1_2[855:848]};
      mid_2[2] = {1'b0,layer_2_2[863:856]} - {1'b0, layer_1_2[863:856]};
      btm_0[0] = {1'b0,layer_3_0[847:840]} - {1'b0, layer_2_0[847:840]};
      btm_0[1] = {1'b0,layer_3_0[855:848]} - {1'b0, layer_2_0[855:848]};
      btm_0[2] = {1'b0,layer_3_0[863:856]} - {1'b0, layer_2_0[863:856]};
      btm_1[0] = {1'b0,layer_3_1[847:840]} - {1'b0, layer_2_1[847:840]};
      btm_1[1] = {1'b0,layer_3_1[855:848]} - {1'b0, layer_2_1[855:848]};
      btm_1[2] = {1'b0,layer_3_1[863:856]} - {1'b0, layer_2_1[863:856]};
      btm_2[0] = {1'b0,layer_3_2[847:840]} - {1'b0, layer_2_2[847:840]};
      btm_2[1] = {1'b0,layer_3_2[855:848]} - {1'b0, layer_2_2[855:848]};
      btm_2[2] = {1'b0,layer_3_2[863:856]} - {1'b0, layer_2_2[863:856]};
    end
    'd107: begin
      top_0[0] = {1'b0,layer_1_0[855:848]} - {1'b0, layer_0_0[855:848]};
      top_0[1] = {1'b0,layer_1_0[863:856]} - {1'b0, layer_0_0[863:856]};
      top_0[2] = {1'b0,layer_1_0[871:864]} - {1'b0, layer_0_0[871:864]};
      top_1[0] = {1'b0,layer_1_1[855:848]} - {1'b0, layer_0_1[855:848]};
      top_1[1] = {1'b0,layer_1_1[863:856]} - {1'b0, layer_0_1[863:856]};
      top_1[2] = {1'b0,layer_1_1[871:864]} - {1'b0, layer_0_1[871:864]};
      top_2[0] = {1'b0,layer_1_2[855:848]} - {1'b0, layer_0_2[855:848]};
      top_2[1] = {1'b0,layer_1_2[863:856]} - {1'b0, layer_0_2[863:856]};
      top_2[2] = {1'b0,layer_1_2[871:864]} - {1'b0, layer_0_2[871:864]};
      mid_0[0] = {1'b0,layer_2_0[855:848]} - {1'b0, layer_1_0[855:848]};
      mid_0[1] = {1'b0,layer_2_0[863:856]} - {1'b0, layer_1_0[863:856]};
      mid_0[2] = {1'b0,layer_2_0[871:864]} - {1'b0, layer_1_0[871:864]};
      mid_1[0] = {1'b0,layer_2_1[855:848]} - {1'b0, layer_1_1[855:848]};
      mid_1[1] = {1'b0,layer_2_1[863:856]} - {1'b0, layer_1_1[863:856]};
      mid_1[2] = {1'b0,layer_2_1[871:864]} - {1'b0, layer_1_1[871:864]};
      mid_2[0] = {1'b0,layer_2_2[855:848]} - {1'b0, layer_1_2[855:848]};
      mid_2[1] = {1'b0,layer_2_2[863:856]} - {1'b0, layer_1_2[863:856]};
      mid_2[2] = {1'b0,layer_2_2[871:864]} - {1'b0, layer_1_2[871:864]};
      btm_0[0] = {1'b0,layer_3_0[855:848]} - {1'b0, layer_2_0[855:848]};
      btm_0[1] = {1'b0,layer_3_0[863:856]} - {1'b0, layer_2_0[863:856]};
      btm_0[2] = {1'b0,layer_3_0[871:864]} - {1'b0, layer_2_0[871:864]};
      btm_1[0] = {1'b0,layer_3_1[855:848]} - {1'b0, layer_2_1[855:848]};
      btm_1[1] = {1'b0,layer_3_1[863:856]} - {1'b0, layer_2_1[863:856]};
      btm_1[2] = {1'b0,layer_3_1[871:864]} - {1'b0, layer_2_1[871:864]};
      btm_2[0] = {1'b0,layer_3_2[855:848]} - {1'b0, layer_2_2[855:848]};
      btm_2[1] = {1'b0,layer_3_2[863:856]} - {1'b0, layer_2_2[863:856]};
      btm_2[2] = {1'b0,layer_3_2[871:864]} - {1'b0, layer_2_2[871:864]};
    end
    'd108: begin
      top_0[0] = {1'b0,layer_1_0[863:856]} - {1'b0, layer_0_0[863:856]};
      top_0[1] = {1'b0,layer_1_0[871:864]} - {1'b0, layer_0_0[871:864]};
      top_0[2] = {1'b0,layer_1_0[879:872]} - {1'b0, layer_0_0[879:872]};
      top_1[0] = {1'b0,layer_1_1[863:856]} - {1'b0, layer_0_1[863:856]};
      top_1[1] = {1'b0,layer_1_1[871:864]} - {1'b0, layer_0_1[871:864]};
      top_1[2] = {1'b0,layer_1_1[879:872]} - {1'b0, layer_0_1[879:872]};
      top_2[0] = {1'b0,layer_1_2[863:856]} - {1'b0, layer_0_2[863:856]};
      top_2[1] = {1'b0,layer_1_2[871:864]} - {1'b0, layer_0_2[871:864]};
      top_2[2] = {1'b0,layer_1_2[879:872]} - {1'b0, layer_0_2[879:872]};
      mid_0[0] = {1'b0,layer_2_0[863:856]} - {1'b0, layer_1_0[863:856]};
      mid_0[1] = {1'b0,layer_2_0[871:864]} - {1'b0, layer_1_0[871:864]};
      mid_0[2] = {1'b0,layer_2_0[879:872]} - {1'b0, layer_1_0[879:872]};
      mid_1[0] = {1'b0,layer_2_1[863:856]} - {1'b0, layer_1_1[863:856]};
      mid_1[1] = {1'b0,layer_2_1[871:864]} - {1'b0, layer_1_1[871:864]};
      mid_1[2] = {1'b0,layer_2_1[879:872]} - {1'b0, layer_1_1[879:872]};
      mid_2[0] = {1'b0,layer_2_2[863:856]} - {1'b0, layer_1_2[863:856]};
      mid_2[1] = {1'b0,layer_2_2[871:864]} - {1'b0, layer_1_2[871:864]};
      mid_2[2] = {1'b0,layer_2_2[879:872]} - {1'b0, layer_1_2[879:872]};
      btm_0[0] = {1'b0,layer_3_0[863:856]} - {1'b0, layer_2_0[863:856]};
      btm_0[1] = {1'b0,layer_3_0[871:864]} - {1'b0, layer_2_0[871:864]};
      btm_0[2] = {1'b0,layer_3_0[879:872]} - {1'b0, layer_2_0[879:872]};
      btm_1[0] = {1'b0,layer_3_1[863:856]} - {1'b0, layer_2_1[863:856]};
      btm_1[1] = {1'b0,layer_3_1[871:864]} - {1'b0, layer_2_1[871:864]};
      btm_1[2] = {1'b0,layer_3_1[879:872]} - {1'b0, layer_2_1[879:872]};
      btm_2[0] = {1'b0,layer_3_2[863:856]} - {1'b0, layer_2_2[863:856]};
      btm_2[1] = {1'b0,layer_3_2[871:864]} - {1'b0, layer_2_2[871:864]};
      btm_2[2] = {1'b0,layer_3_2[879:872]} - {1'b0, layer_2_2[879:872]};
    end
    'd109: begin
      top_0[0] = {1'b0,layer_1_0[871:864]} - {1'b0, layer_0_0[871:864]};
      top_0[1] = {1'b0,layer_1_0[879:872]} - {1'b0, layer_0_0[879:872]};
      top_0[2] = {1'b0,layer_1_0[887:880]} - {1'b0, layer_0_0[887:880]};
      top_1[0] = {1'b0,layer_1_1[871:864]} - {1'b0, layer_0_1[871:864]};
      top_1[1] = {1'b0,layer_1_1[879:872]} - {1'b0, layer_0_1[879:872]};
      top_1[2] = {1'b0,layer_1_1[887:880]} - {1'b0, layer_0_1[887:880]};
      top_2[0] = {1'b0,layer_1_2[871:864]} - {1'b0, layer_0_2[871:864]};
      top_2[1] = {1'b0,layer_1_2[879:872]} - {1'b0, layer_0_2[879:872]};
      top_2[2] = {1'b0,layer_1_2[887:880]} - {1'b0, layer_0_2[887:880]};
      mid_0[0] = {1'b0,layer_2_0[871:864]} - {1'b0, layer_1_0[871:864]};
      mid_0[1] = {1'b0,layer_2_0[879:872]} - {1'b0, layer_1_0[879:872]};
      mid_0[2] = {1'b0,layer_2_0[887:880]} - {1'b0, layer_1_0[887:880]};
      mid_1[0] = {1'b0,layer_2_1[871:864]} - {1'b0, layer_1_1[871:864]};
      mid_1[1] = {1'b0,layer_2_1[879:872]} - {1'b0, layer_1_1[879:872]};
      mid_1[2] = {1'b0,layer_2_1[887:880]} - {1'b0, layer_1_1[887:880]};
      mid_2[0] = {1'b0,layer_2_2[871:864]} - {1'b0, layer_1_2[871:864]};
      mid_2[1] = {1'b0,layer_2_2[879:872]} - {1'b0, layer_1_2[879:872]};
      mid_2[2] = {1'b0,layer_2_2[887:880]} - {1'b0, layer_1_2[887:880]};
      btm_0[0] = {1'b0,layer_3_0[871:864]} - {1'b0, layer_2_0[871:864]};
      btm_0[1] = {1'b0,layer_3_0[879:872]} - {1'b0, layer_2_0[879:872]};
      btm_0[2] = {1'b0,layer_3_0[887:880]} - {1'b0, layer_2_0[887:880]};
      btm_1[0] = {1'b0,layer_3_1[871:864]} - {1'b0, layer_2_1[871:864]};
      btm_1[1] = {1'b0,layer_3_1[879:872]} - {1'b0, layer_2_1[879:872]};
      btm_1[2] = {1'b0,layer_3_1[887:880]} - {1'b0, layer_2_1[887:880]};
      btm_2[0] = {1'b0,layer_3_2[871:864]} - {1'b0, layer_2_2[871:864]};
      btm_2[1] = {1'b0,layer_3_2[879:872]} - {1'b0, layer_2_2[879:872]};
      btm_2[2] = {1'b0,layer_3_2[887:880]} - {1'b0, layer_2_2[887:880]};
    end
    'd110: begin
      top_0[0] = {1'b0,layer_1_0[879:872]} - {1'b0, layer_0_0[879:872]};
      top_0[1] = {1'b0,layer_1_0[887:880]} - {1'b0, layer_0_0[887:880]};
      top_0[2] = {1'b0,layer_1_0[895:888]} - {1'b0, layer_0_0[895:888]};
      top_1[0] = {1'b0,layer_1_1[879:872]} - {1'b0, layer_0_1[879:872]};
      top_1[1] = {1'b0,layer_1_1[887:880]} - {1'b0, layer_0_1[887:880]};
      top_1[2] = {1'b0,layer_1_1[895:888]} - {1'b0, layer_0_1[895:888]};
      top_2[0] = {1'b0,layer_1_2[879:872]} - {1'b0, layer_0_2[879:872]};
      top_2[1] = {1'b0,layer_1_2[887:880]} - {1'b0, layer_0_2[887:880]};
      top_2[2] = {1'b0,layer_1_2[895:888]} - {1'b0, layer_0_2[895:888]};
      mid_0[0] = {1'b0,layer_2_0[879:872]} - {1'b0, layer_1_0[879:872]};
      mid_0[1] = {1'b0,layer_2_0[887:880]} - {1'b0, layer_1_0[887:880]};
      mid_0[2] = {1'b0,layer_2_0[895:888]} - {1'b0, layer_1_0[895:888]};
      mid_1[0] = {1'b0,layer_2_1[879:872]} - {1'b0, layer_1_1[879:872]};
      mid_1[1] = {1'b0,layer_2_1[887:880]} - {1'b0, layer_1_1[887:880]};
      mid_1[2] = {1'b0,layer_2_1[895:888]} - {1'b0, layer_1_1[895:888]};
      mid_2[0] = {1'b0,layer_2_2[879:872]} - {1'b0, layer_1_2[879:872]};
      mid_2[1] = {1'b0,layer_2_2[887:880]} - {1'b0, layer_1_2[887:880]};
      mid_2[2] = {1'b0,layer_2_2[895:888]} - {1'b0, layer_1_2[895:888]};
      btm_0[0] = {1'b0,layer_3_0[879:872]} - {1'b0, layer_2_0[879:872]};
      btm_0[1] = {1'b0,layer_3_0[887:880]} - {1'b0, layer_2_0[887:880]};
      btm_0[2] = {1'b0,layer_3_0[895:888]} - {1'b0, layer_2_0[895:888]};
      btm_1[0] = {1'b0,layer_3_1[879:872]} - {1'b0, layer_2_1[879:872]};
      btm_1[1] = {1'b0,layer_3_1[887:880]} - {1'b0, layer_2_1[887:880]};
      btm_1[2] = {1'b0,layer_3_1[895:888]} - {1'b0, layer_2_1[895:888]};
      btm_2[0] = {1'b0,layer_3_2[879:872]} - {1'b0, layer_2_2[879:872]};
      btm_2[1] = {1'b0,layer_3_2[887:880]} - {1'b0, layer_2_2[887:880]};
      btm_2[2] = {1'b0,layer_3_2[895:888]} - {1'b0, layer_2_2[895:888]};
    end
    'd111: begin
      top_0[0] = {1'b0,layer_1_0[887:880]} - {1'b0, layer_0_0[887:880]};
      top_0[1] = {1'b0,layer_1_0[895:888]} - {1'b0, layer_0_0[895:888]};
      top_0[2] = {1'b0,layer_1_0[903:896]} - {1'b0, layer_0_0[903:896]};
      top_1[0] = {1'b0,layer_1_1[887:880]} - {1'b0, layer_0_1[887:880]};
      top_1[1] = {1'b0,layer_1_1[895:888]} - {1'b0, layer_0_1[895:888]};
      top_1[2] = {1'b0,layer_1_1[903:896]} - {1'b0, layer_0_1[903:896]};
      top_2[0] = {1'b0,layer_1_2[887:880]} - {1'b0, layer_0_2[887:880]};
      top_2[1] = {1'b0,layer_1_2[895:888]} - {1'b0, layer_0_2[895:888]};
      top_2[2] = {1'b0,layer_1_2[903:896]} - {1'b0, layer_0_2[903:896]};
      mid_0[0] = {1'b0,layer_2_0[887:880]} - {1'b0, layer_1_0[887:880]};
      mid_0[1] = {1'b0,layer_2_0[895:888]} - {1'b0, layer_1_0[895:888]};
      mid_0[2] = {1'b0,layer_2_0[903:896]} - {1'b0, layer_1_0[903:896]};
      mid_1[0] = {1'b0,layer_2_1[887:880]} - {1'b0, layer_1_1[887:880]};
      mid_1[1] = {1'b0,layer_2_1[895:888]} - {1'b0, layer_1_1[895:888]};
      mid_1[2] = {1'b0,layer_2_1[903:896]} - {1'b0, layer_1_1[903:896]};
      mid_2[0] = {1'b0,layer_2_2[887:880]} - {1'b0, layer_1_2[887:880]};
      mid_2[1] = {1'b0,layer_2_2[895:888]} - {1'b0, layer_1_2[895:888]};
      mid_2[2] = {1'b0,layer_2_2[903:896]} - {1'b0, layer_1_2[903:896]};
      btm_0[0] = {1'b0,layer_3_0[887:880]} - {1'b0, layer_2_0[887:880]};
      btm_0[1] = {1'b0,layer_3_0[895:888]} - {1'b0, layer_2_0[895:888]};
      btm_0[2] = {1'b0,layer_3_0[903:896]} - {1'b0, layer_2_0[903:896]};
      btm_1[0] = {1'b0,layer_3_1[887:880]} - {1'b0, layer_2_1[887:880]};
      btm_1[1] = {1'b0,layer_3_1[895:888]} - {1'b0, layer_2_1[895:888]};
      btm_1[2] = {1'b0,layer_3_1[903:896]} - {1'b0, layer_2_1[903:896]};
      btm_2[0] = {1'b0,layer_3_2[887:880]} - {1'b0, layer_2_2[887:880]};
      btm_2[1] = {1'b0,layer_3_2[895:888]} - {1'b0, layer_2_2[895:888]};
      btm_2[2] = {1'b0,layer_3_2[903:896]} - {1'b0, layer_2_2[903:896]};
    end
    'd112: begin
      top_0[0] = {1'b0,layer_1_0[895:888]} - {1'b0, layer_0_0[895:888]};
      top_0[1] = {1'b0,layer_1_0[903:896]} - {1'b0, layer_0_0[903:896]};
      top_0[2] = {1'b0,layer_1_0[911:904]} - {1'b0, layer_0_0[911:904]};
      top_1[0] = {1'b0,layer_1_1[895:888]} - {1'b0, layer_0_1[895:888]};
      top_1[1] = {1'b0,layer_1_1[903:896]} - {1'b0, layer_0_1[903:896]};
      top_1[2] = {1'b0,layer_1_1[911:904]} - {1'b0, layer_0_1[911:904]};
      top_2[0] = {1'b0,layer_1_2[895:888]} - {1'b0, layer_0_2[895:888]};
      top_2[1] = {1'b0,layer_1_2[903:896]} - {1'b0, layer_0_2[903:896]};
      top_2[2] = {1'b0,layer_1_2[911:904]} - {1'b0, layer_0_2[911:904]};
      mid_0[0] = {1'b0,layer_2_0[895:888]} - {1'b0, layer_1_0[895:888]};
      mid_0[1] = {1'b0,layer_2_0[903:896]} - {1'b0, layer_1_0[903:896]};
      mid_0[2] = {1'b0,layer_2_0[911:904]} - {1'b0, layer_1_0[911:904]};
      mid_1[0] = {1'b0,layer_2_1[895:888]} - {1'b0, layer_1_1[895:888]};
      mid_1[1] = {1'b0,layer_2_1[903:896]} - {1'b0, layer_1_1[903:896]};
      mid_1[2] = {1'b0,layer_2_1[911:904]} - {1'b0, layer_1_1[911:904]};
      mid_2[0] = {1'b0,layer_2_2[895:888]} - {1'b0, layer_1_2[895:888]};
      mid_2[1] = {1'b0,layer_2_2[903:896]} - {1'b0, layer_1_2[903:896]};
      mid_2[2] = {1'b0,layer_2_2[911:904]} - {1'b0, layer_1_2[911:904]};
      btm_0[0] = {1'b0,layer_3_0[895:888]} - {1'b0, layer_2_0[895:888]};
      btm_0[1] = {1'b0,layer_3_0[903:896]} - {1'b0, layer_2_0[903:896]};
      btm_0[2] = {1'b0,layer_3_0[911:904]} - {1'b0, layer_2_0[911:904]};
      btm_1[0] = {1'b0,layer_3_1[895:888]} - {1'b0, layer_2_1[895:888]};
      btm_1[1] = {1'b0,layer_3_1[903:896]} - {1'b0, layer_2_1[903:896]};
      btm_1[2] = {1'b0,layer_3_1[911:904]} - {1'b0, layer_2_1[911:904]};
      btm_2[0] = {1'b0,layer_3_2[895:888]} - {1'b0, layer_2_2[895:888]};
      btm_2[1] = {1'b0,layer_3_2[903:896]} - {1'b0, layer_2_2[903:896]};
      btm_2[2] = {1'b0,layer_3_2[911:904]} - {1'b0, layer_2_2[911:904]};
    end
    'd113: begin
      top_0[0] = {1'b0,layer_1_0[903:896]} - {1'b0, layer_0_0[903:896]};
      top_0[1] = {1'b0,layer_1_0[911:904]} - {1'b0, layer_0_0[911:904]};
      top_0[2] = {1'b0,layer_1_0[919:912]} - {1'b0, layer_0_0[919:912]};
      top_1[0] = {1'b0,layer_1_1[903:896]} - {1'b0, layer_0_1[903:896]};
      top_1[1] = {1'b0,layer_1_1[911:904]} - {1'b0, layer_0_1[911:904]};
      top_1[2] = {1'b0,layer_1_1[919:912]} - {1'b0, layer_0_1[919:912]};
      top_2[0] = {1'b0,layer_1_2[903:896]} - {1'b0, layer_0_2[903:896]};
      top_2[1] = {1'b0,layer_1_2[911:904]} - {1'b0, layer_0_2[911:904]};
      top_2[2] = {1'b0,layer_1_2[919:912]} - {1'b0, layer_0_2[919:912]};
      mid_0[0] = {1'b0,layer_2_0[903:896]} - {1'b0, layer_1_0[903:896]};
      mid_0[1] = {1'b0,layer_2_0[911:904]} - {1'b0, layer_1_0[911:904]};
      mid_0[2] = {1'b0,layer_2_0[919:912]} - {1'b0, layer_1_0[919:912]};
      mid_1[0] = {1'b0,layer_2_1[903:896]} - {1'b0, layer_1_1[903:896]};
      mid_1[1] = {1'b0,layer_2_1[911:904]} - {1'b0, layer_1_1[911:904]};
      mid_1[2] = {1'b0,layer_2_1[919:912]} - {1'b0, layer_1_1[919:912]};
      mid_2[0] = {1'b0,layer_2_2[903:896]} - {1'b0, layer_1_2[903:896]};
      mid_2[1] = {1'b0,layer_2_2[911:904]} - {1'b0, layer_1_2[911:904]};
      mid_2[2] = {1'b0,layer_2_2[919:912]} - {1'b0, layer_1_2[919:912]};
      btm_0[0] = {1'b0,layer_3_0[903:896]} - {1'b0, layer_2_0[903:896]};
      btm_0[1] = {1'b0,layer_3_0[911:904]} - {1'b0, layer_2_0[911:904]};
      btm_0[2] = {1'b0,layer_3_0[919:912]} - {1'b0, layer_2_0[919:912]};
      btm_1[0] = {1'b0,layer_3_1[903:896]} - {1'b0, layer_2_1[903:896]};
      btm_1[1] = {1'b0,layer_3_1[911:904]} - {1'b0, layer_2_1[911:904]};
      btm_1[2] = {1'b0,layer_3_1[919:912]} - {1'b0, layer_2_1[919:912]};
      btm_2[0] = {1'b0,layer_3_2[903:896]} - {1'b0, layer_2_2[903:896]};
      btm_2[1] = {1'b0,layer_3_2[911:904]} - {1'b0, layer_2_2[911:904]};
      btm_2[2] = {1'b0,layer_3_2[919:912]} - {1'b0, layer_2_2[919:912]};
    end
    'd114: begin
      top_0[0] = {1'b0,layer_1_0[911:904]} - {1'b0, layer_0_0[911:904]};
      top_0[1] = {1'b0,layer_1_0[919:912]} - {1'b0, layer_0_0[919:912]};
      top_0[2] = {1'b0,layer_1_0[927:920]} - {1'b0, layer_0_0[927:920]};
      top_1[0] = {1'b0,layer_1_1[911:904]} - {1'b0, layer_0_1[911:904]};
      top_1[1] = {1'b0,layer_1_1[919:912]} - {1'b0, layer_0_1[919:912]};
      top_1[2] = {1'b0,layer_1_1[927:920]} - {1'b0, layer_0_1[927:920]};
      top_2[0] = {1'b0,layer_1_2[911:904]} - {1'b0, layer_0_2[911:904]};
      top_2[1] = {1'b0,layer_1_2[919:912]} - {1'b0, layer_0_2[919:912]};
      top_2[2] = {1'b0,layer_1_2[927:920]} - {1'b0, layer_0_2[927:920]};
      mid_0[0] = {1'b0,layer_2_0[911:904]} - {1'b0, layer_1_0[911:904]};
      mid_0[1] = {1'b0,layer_2_0[919:912]} - {1'b0, layer_1_0[919:912]};
      mid_0[2] = {1'b0,layer_2_0[927:920]} - {1'b0, layer_1_0[927:920]};
      mid_1[0] = {1'b0,layer_2_1[911:904]} - {1'b0, layer_1_1[911:904]};
      mid_1[1] = {1'b0,layer_2_1[919:912]} - {1'b0, layer_1_1[919:912]};
      mid_1[2] = {1'b0,layer_2_1[927:920]} - {1'b0, layer_1_1[927:920]};
      mid_2[0] = {1'b0,layer_2_2[911:904]} - {1'b0, layer_1_2[911:904]};
      mid_2[1] = {1'b0,layer_2_2[919:912]} - {1'b0, layer_1_2[919:912]};
      mid_2[2] = {1'b0,layer_2_2[927:920]} - {1'b0, layer_1_2[927:920]};
      btm_0[0] = {1'b0,layer_3_0[911:904]} - {1'b0, layer_2_0[911:904]};
      btm_0[1] = {1'b0,layer_3_0[919:912]} - {1'b0, layer_2_0[919:912]};
      btm_0[2] = {1'b0,layer_3_0[927:920]} - {1'b0, layer_2_0[927:920]};
      btm_1[0] = {1'b0,layer_3_1[911:904]} - {1'b0, layer_2_1[911:904]};
      btm_1[1] = {1'b0,layer_3_1[919:912]} - {1'b0, layer_2_1[919:912]};
      btm_1[2] = {1'b0,layer_3_1[927:920]} - {1'b0, layer_2_1[927:920]};
      btm_2[0] = {1'b0,layer_3_2[911:904]} - {1'b0, layer_2_2[911:904]};
      btm_2[1] = {1'b0,layer_3_2[919:912]} - {1'b0, layer_2_2[919:912]};
      btm_2[2] = {1'b0,layer_3_2[927:920]} - {1'b0, layer_2_2[927:920]};
    end
    'd115: begin
      top_0[0] = {1'b0,layer_1_0[919:912]} - {1'b0, layer_0_0[919:912]};
      top_0[1] = {1'b0,layer_1_0[927:920]} - {1'b0, layer_0_0[927:920]};
      top_0[2] = {1'b0,layer_1_0[935:928]} - {1'b0, layer_0_0[935:928]};
      top_1[0] = {1'b0,layer_1_1[919:912]} - {1'b0, layer_0_1[919:912]};
      top_1[1] = {1'b0,layer_1_1[927:920]} - {1'b0, layer_0_1[927:920]};
      top_1[2] = {1'b0,layer_1_1[935:928]} - {1'b0, layer_0_1[935:928]};
      top_2[0] = {1'b0,layer_1_2[919:912]} - {1'b0, layer_0_2[919:912]};
      top_2[1] = {1'b0,layer_1_2[927:920]} - {1'b0, layer_0_2[927:920]};
      top_2[2] = {1'b0,layer_1_2[935:928]} - {1'b0, layer_0_2[935:928]};
      mid_0[0] = {1'b0,layer_2_0[919:912]} - {1'b0, layer_1_0[919:912]};
      mid_0[1] = {1'b0,layer_2_0[927:920]} - {1'b0, layer_1_0[927:920]};
      mid_0[2] = {1'b0,layer_2_0[935:928]} - {1'b0, layer_1_0[935:928]};
      mid_1[0] = {1'b0,layer_2_1[919:912]} - {1'b0, layer_1_1[919:912]};
      mid_1[1] = {1'b0,layer_2_1[927:920]} - {1'b0, layer_1_1[927:920]};
      mid_1[2] = {1'b0,layer_2_1[935:928]} - {1'b0, layer_1_1[935:928]};
      mid_2[0] = {1'b0,layer_2_2[919:912]} - {1'b0, layer_1_2[919:912]};
      mid_2[1] = {1'b0,layer_2_2[927:920]} - {1'b0, layer_1_2[927:920]};
      mid_2[2] = {1'b0,layer_2_2[935:928]} - {1'b0, layer_1_2[935:928]};
      btm_0[0] = {1'b0,layer_3_0[919:912]} - {1'b0, layer_2_0[919:912]};
      btm_0[1] = {1'b0,layer_3_0[927:920]} - {1'b0, layer_2_0[927:920]};
      btm_0[2] = {1'b0,layer_3_0[935:928]} - {1'b0, layer_2_0[935:928]};
      btm_1[0] = {1'b0,layer_3_1[919:912]} - {1'b0, layer_2_1[919:912]};
      btm_1[1] = {1'b0,layer_3_1[927:920]} - {1'b0, layer_2_1[927:920]};
      btm_1[2] = {1'b0,layer_3_1[935:928]} - {1'b0, layer_2_1[935:928]};
      btm_2[0] = {1'b0,layer_3_2[919:912]} - {1'b0, layer_2_2[919:912]};
      btm_2[1] = {1'b0,layer_3_2[927:920]} - {1'b0, layer_2_2[927:920]};
      btm_2[2] = {1'b0,layer_3_2[935:928]} - {1'b0, layer_2_2[935:928]};
    end
    'd116: begin
      top_0[0] = {1'b0,layer_1_0[927:920]} - {1'b0, layer_0_0[927:920]};
      top_0[1] = {1'b0,layer_1_0[935:928]} - {1'b0, layer_0_0[935:928]};
      top_0[2] = {1'b0,layer_1_0[943:936]} - {1'b0, layer_0_0[943:936]};
      top_1[0] = {1'b0,layer_1_1[927:920]} - {1'b0, layer_0_1[927:920]};
      top_1[1] = {1'b0,layer_1_1[935:928]} - {1'b0, layer_0_1[935:928]};
      top_1[2] = {1'b0,layer_1_1[943:936]} - {1'b0, layer_0_1[943:936]};
      top_2[0] = {1'b0,layer_1_2[927:920]} - {1'b0, layer_0_2[927:920]};
      top_2[1] = {1'b0,layer_1_2[935:928]} - {1'b0, layer_0_2[935:928]};
      top_2[2] = {1'b0,layer_1_2[943:936]} - {1'b0, layer_0_2[943:936]};
      mid_0[0] = {1'b0,layer_2_0[927:920]} - {1'b0, layer_1_0[927:920]};
      mid_0[1] = {1'b0,layer_2_0[935:928]} - {1'b0, layer_1_0[935:928]};
      mid_0[2] = {1'b0,layer_2_0[943:936]} - {1'b0, layer_1_0[943:936]};
      mid_1[0] = {1'b0,layer_2_1[927:920]} - {1'b0, layer_1_1[927:920]};
      mid_1[1] = {1'b0,layer_2_1[935:928]} - {1'b0, layer_1_1[935:928]};
      mid_1[2] = {1'b0,layer_2_1[943:936]} - {1'b0, layer_1_1[943:936]};
      mid_2[0] = {1'b0,layer_2_2[927:920]} - {1'b0, layer_1_2[927:920]};
      mid_2[1] = {1'b0,layer_2_2[935:928]} - {1'b0, layer_1_2[935:928]};
      mid_2[2] = {1'b0,layer_2_2[943:936]} - {1'b0, layer_1_2[943:936]};
      btm_0[0] = {1'b0,layer_3_0[927:920]} - {1'b0, layer_2_0[927:920]};
      btm_0[1] = {1'b0,layer_3_0[935:928]} - {1'b0, layer_2_0[935:928]};
      btm_0[2] = {1'b0,layer_3_0[943:936]} - {1'b0, layer_2_0[943:936]};
      btm_1[0] = {1'b0,layer_3_1[927:920]} - {1'b0, layer_2_1[927:920]};
      btm_1[1] = {1'b0,layer_3_1[935:928]} - {1'b0, layer_2_1[935:928]};
      btm_1[2] = {1'b0,layer_3_1[943:936]} - {1'b0, layer_2_1[943:936]};
      btm_2[0] = {1'b0,layer_3_2[927:920]} - {1'b0, layer_2_2[927:920]};
      btm_2[1] = {1'b0,layer_3_2[935:928]} - {1'b0, layer_2_2[935:928]};
      btm_2[2] = {1'b0,layer_3_2[943:936]} - {1'b0, layer_2_2[943:936]};
    end
    'd117: begin
      top_0[0] = {1'b0,layer_1_0[935:928]} - {1'b0, layer_0_0[935:928]};
      top_0[1] = {1'b0,layer_1_0[943:936]} - {1'b0, layer_0_0[943:936]};
      top_0[2] = {1'b0,layer_1_0[951:944]} - {1'b0, layer_0_0[951:944]};
      top_1[0] = {1'b0,layer_1_1[935:928]} - {1'b0, layer_0_1[935:928]};
      top_1[1] = {1'b0,layer_1_1[943:936]} - {1'b0, layer_0_1[943:936]};
      top_1[2] = {1'b0,layer_1_1[951:944]} - {1'b0, layer_0_1[951:944]};
      top_2[0] = {1'b0,layer_1_2[935:928]} - {1'b0, layer_0_2[935:928]};
      top_2[1] = {1'b0,layer_1_2[943:936]} - {1'b0, layer_0_2[943:936]};
      top_2[2] = {1'b0,layer_1_2[951:944]} - {1'b0, layer_0_2[951:944]};
      mid_0[0] = {1'b0,layer_2_0[935:928]} - {1'b0, layer_1_0[935:928]};
      mid_0[1] = {1'b0,layer_2_0[943:936]} - {1'b0, layer_1_0[943:936]};
      mid_0[2] = {1'b0,layer_2_0[951:944]} - {1'b0, layer_1_0[951:944]};
      mid_1[0] = {1'b0,layer_2_1[935:928]} - {1'b0, layer_1_1[935:928]};
      mid_1[1] = {1'b0,layer_2_1[943:936]} - {1'b0, layer_1_1[943:936]};
      mid_1[2] = {1'b0,layer_2_1[951:944]} - {1'b0, layer_1_1[951:944]};
      mid_2[0] = {1'b0,layer_2_2[935:928]} - {1'b0, layer_1_2[935:928]};
      mid_2[1] = {1'b0,layer_2_2[943:936]} - {1'b0, layer_1_2[943:936]};
      mid_2[2] = {1'b0,layer_2_2[951:944]} - {1'b0, layer_1_2[951:944]};
      btm_0[0] = {1'b0,layer_3_0[935:928]} - {1'b0, layer_2_0[935:928]};
      btm_0[1] = {1'b0,layer_3_0[943:936]} - {1'b0, layer_2_0[943:936]};
      btm_0[2] = {1'b0,layer_3_0[951:944]} - {1'b0, layer_2_0[951:944]};
      btm_1[0] = {1'b0,layer_3_1[935:928]} - {1'b0, layer_2_1[935:928]};
      btm_1[1] = {1'b0,layer_3_1[943:936]} - {1'b0, layer_2_1[943:936]};
      btm_1[2] = {1'b0,layer_3_1[951:944]} - {1'b0, layer_2_1[951:944]};
      btm_2[0] = {1'b0,layer_3_2[935:928]} - {1'b0, layer_2_2[935:928]};
      btm_2[1] = {1'b0,layer_3_2[943:936]} - {1'b0, layer_2_2[943:936]};
      btm_2[2] = {1'b0,layer_3_2[951:944]} - {1'b0, layer_2_2[951:944]};
    end
    'd118: begin
      top_0[0] = {1'b0,layer_1_0[943:936]} - {1'b0, layer_0_0[943:936]};
      top_0[1] = {1'b0,layer_1_0[951:944]} - {1'b0, layer_0_0[951:944]};
      top_0[2] = {1'b0,layer_1_0[959:952]} - {1'b0, layer_0_0[959:952]};
      top_1[0] = {1'b0,layer_1_1[943:936]} - {1'b0, layer_0_1[943:936]};
      top_1[1] = {1'b0,layer_1_1[951:944]} - {1'b0, layer_0_1[951:944]};
      top_1[2] = {1'b0,layer_1_1[959:952]} - {1'b0, layer_0_1[959:952]};
      top_2[0] = {1'b0,layer_1_2[943:936]} - {1'b0, layer_0_2[943:936]};
      top_2[1] = {1'b0,layer_1_2[951:944]} - {1'b0, layer_0_2[951:944]};
      top_2[2] = {1'b0,layer_1_2[959:952]} - {1'b0, layer_0_2[959:952]};
      mid_0[0] = {1'b0,layer_2_0[943:936]} - {1'b0, layer_1_0[943:936]};
      mid_0[1] = {1'b0,layer_2_0[951:944]} - {1'b0, layer_1_0[951:944]};
      mid_0[2] = {1'b0,layer_2_0[959:952]} - {1'b0, layer_1_0[959:952]};
      mid_1[0] = {1'b0,layer_2_1[943:936]} - {1'b0, layer_1_1[943:936]};
      mid_1[1] = {1'b0,layer_2_1[951:944]} - {1'b0, layer_1_1[951:944]};
      mid_1[2] = {1'b0,layer_2_1[959:952]} - {1'b0, layer_1_1[959:952]};
      mid_2[0] = {1'b0,layer_2_2[943:936]} - {1'b0, layer_1_2[943:936]};
      mid_2[1] = {1'b0,layer_2_2[951:944]} - {1'b0, layer_1_2[951:944]};
      mid_2[2] = {1'b0,layer_2_2[959:952]} - {1'b0, layer_1_2[959:952]};
      btm_0[0] = {1'b0,layer_3_0[943:936]} - {1'b0, layer_2_0[943:936]};
      btm_0[1] = {1'b0,layer_3_0[951:944]} - {1'b0, layer_2_0[951:944]};
      btm_0[2] = {1'b0,layer_3_0[959:952]} - {1'b0, layer_2_0[959:952]};
      btm_1[0] = {1'b0,layer_3_1[943:936]} - {1'b0, layer_2_1[943:936]};
      btm_1[1] = {1'b0,layer_3_1[951:944]} - {1'b0, layer_2_1[951:944]};
      btm_1[2] = {1'b0,layer_3_1[959:952]} - {1'b0, layer_2_1[959:952]};
      btm_2[0] = {1'b0,layer_3_2[943:936]} - {1'b0, layer_2_2[943:936]};
      btm_2[1] = {1'b0,layer_3_2[951:944]} - {1'b0, layer_2_2[951:944]};
      btm_2[2] = {1'b0,layer_3_2[959:952]} - {1'b0, layer_2_2[959:952]};
    end
    'd119: begin
      top_0[0] = {1'b0,layer_1_0[951:944]} - {1'b0, layer_0_0[951:944]};
      top_0[1] = {1'b0,layer_1_0[959:952]} - {1'b0, layer_0_0[959:952]};
      top_0[2] = {1'b0,layer_1_0[967:960]} - {1'b0, layer_0_0[967:960]};
      top_1[0] = {1'b0,layer_1_1[951:944]} - {1'b0, layer_0_1[951:944]};
      top_1[1] = {1'b0,layer_1_1[959:952]} - {1'b0, layer_0_1[959:952]};
      top_1[2] = {1'b0,layer_1_1[967:960]} - {1'b0, layer_0_1[967:960]};
      top_2[0] = {1'b0,layer_1_2[951:944]} - {1'b0, layer_0_2[951:944]};
      top_2[1] = {1'b0,layer_1_2[959:952]} - {1'b0, layer_0_2[959:952]};
      top_2[2] = {1'b0,layer_1_2[967:960]} - {1'b0, layer_0_2[967:960]};
      mid_0[0] = {1'b0,layer_2_0[951:944]} - {1'b0, layer_1_0[951:944]};
      mid_0[1] = {1'b0,layer_2_0[959:952]} - {1'b0, layer_1_0[959:952]};
      mid_0[2] = {1'b0,layer_2_0[967:960]} - {1'b0, layer_1_0[967:960]};
      mid_1[0] = {1'b0,layer_2_1[951:944]} - {1'b0, layer_1_1[951:944]};
      mid_1[1] = {1'b0,layer_2_1[959:952]} - {1'b0, layer_1_1[959:952]};
      mid_1[2] = {1'b0,layer_2_1[967:960]} - {1'b0, layer_1_1[967:960]};
      mid_2[0] = {1'b0,layer_2_2[951:944]} - {1'b0, layer_1_2[951:944]};
      mid_2[1] = {1'b0,layer_2_2[959:952]} - {1'b0, layer_1_2[959:952]};
      mid_2[2] = {1'b0,layer_2_2[967:960]} - {1'b0, layer_1_2[967:960]};
      btm_0[0] = {1'b0,layer_3_0[951:944]} - {1'b0, layer_2_0[951:944]};
      btm_0[1] = {1'b0,layer_3_0[959:952]} - {1'b0, layer_2_0[959:952]};
      btm_0[2] = {1'b0,layer_3_0[967:960]} - {1'b0, layer_2_0[967:960]};
      btm_1[0] = {1'b0,layer_3_1[951:944]} - {1'b0, layer_2_1[951:944]};
      btm_1[1] = {1'b0,layer_3_1[959:952]} - {1'b0, layer_2_1[959:952]};
      btm_1[2] = {1'b0,layer_3_1[967:960]} - {1'b0, layer_2_1[967:960]};
      btm_2[0] = {1'b0,layer_3_2[951:944]} - {1'b0, layer_2_2[951:944]};
      btm_2[1] = {1'b0,layer_3_2[959:952]} - {1'b0, layer_2_2[959:952]};
      btm_2[2] = {1'b0,layer_3_2[967:960]} - {1'b0, layer_2_2[967:960]};
    end
    'd120: begin
      top_0[0] = {1'b0,layer_1_0[959:952]} - {1'b0, layer_0_0[959:952]};
      top_0[1] = {1'b0,layer_1_0[967:960]} - {1'b0, layer_0_0[967:960]};
      top_0[2] = {1'b0,layer_1_0[975:968]} - {1'b0, layer_0_0[975:968]};
      top_1[0] = {1'b0,layer_1_1[959:952]} - {1'b0, layer_0_1[959:952]};
      top_1[1] = {1'b0,layer_1_1[967:960]} - {1'b0, layer_0_1[967:960]};
      top_1[2] = {1'b0,layer_1_1[975:968]} - {1'b0, layer_0_1[975:968]};
      top_2[0] = {1'b0,layer_1_2[959:952]} - {1'b0, layer_0_2[959:952]};
      top_2[1] = {1'b0,layer_1_2[967:960]} - {1'b0, layer_0_2[967:960]};
      top_2[2] = {1'b0,layer_1_2[975:968]} - {1'b0, layer_0_2[975:968]};
      mid_0[0] = {1'b0,layer_2_0[959:952]} - {1'b0, layer_1_0[959:952]};
      mid_0[1] = {1'b0,layer_2_0[967:960]} - {1'b0, layer_1_0[967:960]};
      mid_0[2] = {1'b0,layer_2_0[975:968]} - {1'b0, layer_1_0[975:968]};
      mid_1[0] = {1'b0,layer_2_1[959:952]} - {1'b0, layer_1_1[959:952]};
      mid_1[1] = {1'b0,layer_2_1[967:960]} - {1'b0, layer_1_1[967:960]};
      mid_1[2] = {1'b0,layer_2_1[975:968]} - {1'b0, layer_1_1[975:968]};
      mid_2[0] = {1'b0,layer_2_2[959:952]} - {1'b0, layer_1_2[959:952]};
      mid_2[1] = {1'b0,layer_2_2[967:960]} - {1'b0, layer_1_2[967:960]};
      mid_2[2] = {1'b0,layer_2_2[975:968]} - {1'b0, layer_1_2[975:968]};
      btm_0[0] = {1'b0,layer_3_0[959:952]} - {1'b0, layer_2_0[959:952]};
      btm_0[1] = {1'b0,layer_3_0[967:960]} - {1'b0, layer_2_0[967:960]};
      btm_0[2] = {1'b0,layer_3_0[975:968]} - {1'b0, layer_2_0[975:968]};
      btm_1[0] = {1'b0,layer_3_1[959:952]} - {1'b0, layer_2_1[959:952]};
      btm_1[1] = {1'b0,layer_3_1[967:960]} - {1'b0, layer_2_1[967:960]};
      btm_1[2] = {1'b0,layer_3_1[975:968]} - {1'b0, layer_2_1[975:968]};
      btm_2[0] = {1'b0,layer_3_2[959:952]} - {1'b0, layer_2_2[959:952]};
      btm_2[1] = {1'b0,layer_3_2[967:960]} - {1'b0, layer_2_2[967:960]};
      btm_2[2] = {1'b0,layer_3_2[975:968]} - {1'b0, layer_2_2[975:968]};
    end
    'd121: begin
      top_0[0] = {1'b0,layer_1_0[967:960]} - {1'b0, layer_0_0[967:960]};
      top_0[1] = {1'b0,layer_1_0[975:968]} - {1'b0, layer_0_0[975:968]};
      top_0[2] = {1'b0,layer_1_0[983:976]} - {1'b0, layer_0_0[983:976]};
      top_1[0] = {1'b0,layer_1_1[967:960]} - {1'b0, layer_0_1[967:960]};
      top_1[1] = {1'b0,layer_1_1[975:968]} - {1'b0, layer_0_1[975:968]};
      top_1[2] = {1'b0,layer_1_1[983:976]} - {1'b0, layer_0_1[983:976]};
      top_2[0] = {1'b0,layer_1_2[967:960]} - {1'b0, layer_0_2[967:960]};
      top_2[1] = {1'b0,layer_1_2[975:968]} - {1'b0, layer_0_2[975:968]};
      top_2[2] = {1'b0,layer_1_2[983:976]} - {1'b0, layer_0_2[983:976]};
      mid_0[0] = {1'b0,layer_2_0[967:960]} - {1'b0, layer_1_0[967:960]};
      mid_0[1] = {1'b0,layer_2_0[975:968]} - {1'b0, layer_1_0[975:968]};
      mid_0[2] = {1'b0,layer_2_0[983:976]} - {1'b0, layer_1_0[983:976]};
      mid_1[0] = {1'b0,layer_2_1[967:960]} - {1'b0, layer_1_1[967:960]};
      mid_1[1] = {1'b0,layer_2_1[975:968]} - {1'b0, layer_1_1[975:968]};
      mid_1[2] = {1'b0,layer_2_1[983:976]} - {1'b0, layer_1_1[983:976]};
      mid_2[0] = {1'b0,layer_2_2[967:960]} - {1'b0, layer_1_2[967:960]};
      mid_2[1] = {1'b0,layer_2_2[975:968]} - {1'b0, layer_1_2[975:968]};
      mid_2[2] = {1'b0,layer_2_2[983:976]} - {1'b0, layer_1_2[983:976]};
      btm_0[0] = {1'b0,layer_3_0[967:960]} - {1'b0, layer_2_0[967:960]};
      btm_0[1] = {1'b0,layer_3_0[975:968]} - {1'b0, layer_2_0[975:968]};
      btm_0[2] = {1'b0,layer_3_0[983:976]} - {1'b0, layer_2_0[983:976]};
      btm_1[0] = {1'b0,layer_3_1[967:960]} - {1'b0, layer_2_1[967:960]};
      btm_1[1] = {1'b0,layer_3_1[975:968]} - {1'b0, layer_2_1[975:968]};
      btm_1[2] = {1'b0,layer_3_1[983:976]} - {1'b0, layer_2_1[983:976]};
      btm_2[0] = {1'b0,layer_3_2[967:960]} - {1'b0, layer_2_2[967:960]};
      btm_2[1] = {1'b0,layer_3_2[975:968]} - {1'b0, layer_2_2[975:968]};
      btm_2[2] = {1'b0,layer_3_2[983:976]} - {1'b0, layer_2_2[983:976]};
    end
    'd122: begin
      top_0[0] = {1'b0,layer_1_0[975:968]} - {1'b0, layer_0_0[975:968]};
      top_0[1] = {1'b0,layer_1_0[983:976]} - {1'b0, layer_0_0[983:976]};
      top_0[2] = {1'b0,layer_1_0[991:984]} - {1'b0, layer_0_0[991:984]};
      top_1[0] = {1'b0,layer_1_1[975:968]} - {1'b0, layer_0_1[975:968]};
      top_1[1] = {1'b0,layer_1_1[983:976]} - {1'b0, layer_0_1[983:976]};
      top_1[2] = {1'b0,layer_1_1[991:984]} - {1'b0, layer_0_1[991:984]};
      top_2[0] = {1'b0,layer_1_2[975:968]} - {1'b0, layer_0_2[975:968]};
      top_2[1] = {1'b0,layer_1_2[983:976]} - {1'b0, layer_0_2[983:976]};
      top_2[2] = {1'b0,layer_1_2[991:984]} - {1'b0, layer_0_2[991:984]};
      mid_0[0] = {1'b0,layer_2_0[975:968]} - {1'b0, layer_1_0[975:968]};
      mid_0[1] = {1'b0,layer_2_0[983:976]} - {1'b0, layer_1_0[983:976]};
      mid_0[2] = {1'b0,layer_2_0[991:984]} - {1'b0, layer_1_0[991:984]};
      mid_1[0] = {1'b0,layer_2_1[975:968]} - {1'b0, layer_1_1[975:968]};
      mid_1[1] = {1'b0,layer_2_1[983:976]} - {1'b0, layer_1_1[983:976]};
      mid_1[2] = {1'b0,layer_2_1[991:984]} - {1'b0, layer_1_1[991:984]};
      mid_2[0] = {1'b0,layer_2_2[975:968]} - {1'b0, layer_1_2[975:968]};
      mid_2[1] = {1'b0,layer_2_2[983:976]} - {1'b0, layer_1_2[983:976]};
      mid_2[2] = {1'b0,layer_2_2[991:984]} - {1'b0, layer_1_2[991:984]};
      btm_0[0] = {1'b0,layer_3_0[975:968]} - {1'b0, layer_2_0[975:968]};
      btm_0[1] = {1'b0,layer_3_0[983:976]} - {1'b0, layer_2_0[983:976]};
      btm_0[2] = {1'b0,layer_3_0[991:984]} - {1'b0, layer_2_0[991:984]};
      btm_1[0] = {1'b0,layer_3_1[975:968]} - {1'b0, layer_2_1[975:968]};
      btm_1[1] = {1'b0,layer_3_1[983:976]} - {1'b0, layer_2_1[983:976]};
      btm_1[2] = {1'b0,layer_3_1[991:984]} - {1'b0, layer_2_1[991:984]};
      btm_2[0] = {1'b0,layer_3_2[975:968]} - {1'b0, layer_2_2[975:968]};
      btm_2[1] = {1'b0,layer_3_2[983:976]} - {1'b0, layer_2_2[983:976]};
      btm_2[2] = {1'b0,layer_3_2[991:984]} - {1'b0, layer_2_2[991:984]};
    end
    'd123: begin
      top_0[0] = {1'b0,layer_1_0[983:976]} - {1'b0, layer_0_0[983:976]};
      top_0[1] = {1'b0,layer_1_0[991:984]} - {1'b0, layer_0_0[991:984]};
      top_0[2] = {1'b0,layer_1_0[999:992]} - {1'b0, layer_0_0[999:992]};
      top_1[0] = {1'b0,layer_1_1[983:976]} - {1'b0, layer_0_1[983:976]};
      top_1[1] = {1'b0,layer_1_1[991:984]} - {1'b0, layer_0_1[991:984]};
      top_1[2] = {1'b0,layer_1_1[999:992]} - {1'b0, layer_0_1[999:992]};
      top_2[0] = {1'b0,layer_1_2[983:976]} - {1'b0, layer_0_2[983:976]};
      top_2[1] = {1'b0,layer_1_2[991:984]} - {1'b0, layer_0_2[991:984]};
      top_2[2] = {1'b0,layer_1_2[999:992]} - {1'b0, layer_0_2[999:992]};
      mid_0[0] = {1'b0,layer_2_0[983:976]} - {1'b0, layer_1_0[983:976]};
      mid_0[1] = {1'b0,layer_2_0[991:984]} - {1'b0, layer_1_0[991:984]};
      mid_0[2] = {1'b0,layer_2_0[999:992]} - {1'b0, layer_1_0[999:992]};
      mid_1[0] = {1'b0,layer_2_1[983:976]} - {1'b0, layer_1_1[983:976]};
      mid_1[1] = {1'b0,layer_2_1[991:984]} - {1'b0, layer_1_1[991:984]};
      mid_1[2] = {1'b0,layer_2_1[999:992]} - {1'b0, layer_1_1[999:992]};
      mid_2[0] = {1'b0,layer_2_2[983:976]} - {1'b0, layer_1_2[983:976]};
      mid_2[1] = {1'b0,layer_2_2[991:984]} - {1'b0, layer_1_2[991:984]};
      mid_2[2] = {1'b0,layer_2_2[999:992]} - {1'b0, layer_1_2[999:992]};
      btm_0[0] = {1'b0,layer_3_0[983:976]} - {1'b0, layer_2_0[983:976]};
      btm_0[1] = {1'b0,layer_3_0[991:984]} - {1'b0, layer_2_0[991:984]};
      btm_0[2] = {1'b0,layer_3_0[999:992]} - {1'b0, layer_2_0[999:992]};
      btm_1[0] = {1'b0,layer_3_1[983:976]} - {1'b0, layer_2_1[983:976]};
      btm_1[1] = {1'b0,layer_3_1[991:984]} - {1'b0, layer_2_1[991:984]};
      btm_1[2] = {1'b0,layer_3_1[999:992]} - {1'b0, layer_2_1[999:992]};
      btm_2[0] = {1'b0,layer_3_2[983:976]} - {1'b0, layer_2_2[983:976]};
      btm_2[1] = {1'b0,layer_3_2[991:984]} - {1'b0, layer_2_2[991:984]};
      btm_2[2] = {1'b0,layer_3_2[999:992]} - {1'b0, layer_2_2[999:992]};
    end
    'd124: begin
      top_0[0] = {1'b0,layer_1_0[991:984]} - {1'b0, layer_0_0[991:984]};
      top_0[1] = {1'b0,layer_1_0[999:992]} - {1'b0, layer_0_0[999:992]};
      top_0[2] = {1'b0,layer_1_0[1007:1000]} - {1'b0, layer_0_0[1007:1000]};
      top_1[0] = {1'b0,layer_1_1[991:984]} - {1'b0, layer_0_1[991:984]};
      top_1[1] = {1'b0,layer_1_1[999:992]} - {1'b0, layer_0_1[999:992]};
      top_1[2] = {1'b0,layer_1_1[1007:1000]} - {1'b0, layer_0_1[1007:1000]};
      top_2[0] = {1'b0,layer_1_2[991:984]} - {1'b0, layer_0_2[991:984]};
      top_2[1] = {1'b0,layer_1_2[999:992]} - {1'b0, layer_0_2[999:992]};
      top_2[2] = {1'b0,layer_1_2[1007:1000]} - {1'b0, layer_0_2[1007:1000]};
      mid_0[0] = {1'b0,layer_2_0[991:984]} - {1'b0, layer_1_0[991:984]};
      mid_0[1] = {1'b0,layer_2_0[999:992]} - {1'b0, layer_1_0[999:992]};
      mid_0[2] = {1'b0,layer_2_0[1007:1000]} - {1'b0, layer_1_0[1007:1000]};
      mid_1[0] = {1'b0,layer_2_1[991:984]} - {1'b0, layer_1_1[991:984]};
      mid_1[1] = {1'b0,layer_2_1[999:992]} - {1'b0, layer_1_1[999:992]};
      mid_1[2] = {1'b0,layer_2_1[1007:1000]} - {1'b0, layer_1_1[1007:1000]};
      mid_2[0] = {1'b0,layer_2_2[991:984]} - {1'b0, layer_1_2[991:984]};
      mid_2[1] = {1'b0,layer_2_2[999:992]} - {1'b0, layer_1_2[999:992]};
      mid_2[2] = {1'b0,layer_2_2[1007:1000]} - {1'b0, layer_1_2[1007:1000]};
      btm_0[0] = {1'b0,layer_3_0[991:984]} - {1'b0, layer_2_0[991:984]};
      btm_0[1] = {1'b0,layer_3_0[999:992]} - {1'b0, layer_2_0[999:992]};
      btm_0[2] = {1'b0,layer_3_0[1007:1000]} - {1'b0, layer_2_0[1007:1000]};
      btm_1[0] = {1'b0,layer_3_1[991:984]} - {1'b0, layer_2_1[991:984]};
      btm_1[1] = {1'b0,layer_3_1[999:992]} - {1'b0, layer_2_1[999:992]};
      btm_1[2] = {1'b0,layer_3_1[1007:1000]} - {1'b0, layer_2_1[1007:1000]};
      btm_2[0] = {1'b0,layer_3_2[991:984]} - {1'b0, layer_2_2[991:984]};
      btm_2[1] = {1'b0,layer_3_2[999:992]} - {1'b0, layer_2_2[999:992]};
      btm_2[2] = {1'b0,layer_3_2[1007:1000]} - {1'b0, layer_2_2[1007:1000]};
    end
    'd125: begin
      top_0[0] = {1'b0,layer_1_0[999:992]} - {1'b0, layer_0_0[999:992]};
      top_0[1] = {1'b0,layer_1_0[1007:1000]} - {1'b0, layer_0_0[1007:1000]};
      top_0[2] = {1'b0,layer_1_0[1015:1008]} - {1'b0, layer_0_0[1015:1008]};
      top_1[0] = {1'b0,layer_1_1[999:992]} - {1'b0, layer_0_1[999:992]};
      top_1[1] = {1'b0,layer_1_1[1007:1000]} - {1'b0, layer_0_1[1007:1000]};
      top_1[2] = {1'b0,layer_1_1[1015:1008]} - {1'b0, layer_0_1[1015:1008]};
      top_2[0] = {1'b0,layer_1_2[999:992]} - {1'b0, layer_0_2[999:992]};
      top_2[1] = {1'b0,layer_1_2[1007:1000]} - {1'b0, layer_0_2[1007:1000]};
      top_2[2] = {1'b0,layer_1_2[1015:1008]} - {1'b0, layer_0_2[1015:1008]};
      mid_0[0] = {1'b0,layer_2_0[999:992]} - {1'b0, layer_1_0[999:992]};
      mid_0[1] = {1'b0,layer_2_0[1007:1000]} - {1'b0, layer_1_0[1007:1000]};
      mid_0[2] = {1'b0,layer_2_0[1015:1008]} - {1'b0, layer_1_0[1015:1008]};
      mid_1[0] = {1'b0,layer_2_1[999:992]} - {1'b0, layer_1_1[999:992]};
      mid_1[1] = {1'b0,layer_2_1[1007:1000]} - {1'b0, layer_1_1[1007:1000]};
      mid_1[2] = {1'b0,layer_2_1[1015:1008]} - {1'b0, layer_1_1[1015:1008]};
      mid_2[0] = {1'b0,layer_2_2[999:992]} - {1'b0, layer_1_2[999:992]};
      mid_2[1] = {1'b0,layer_2_2[1007:1000]} - {1'b0, layer_1_2[1007:1000]};
      mid_2[2] = {1'b0,layer_2_2[1015:1008]} - {1'b0, layer_1_2[1015:1008]};
      btm_0[0] = {1'b0,layer_3_0[999:992]} - {1'b0, layer_2_0[999:992]};
      btm_0[1] = {1'b0,layer_3_0[1007:1000]} - {1'b0, layer_2_0[1007:1000]};
      btm_0[2] = {1'b0,layer_3_0[1015:1008]} - {1'b0, layer_2_0[1015:1008]};
      btm_1[0] = {1'b0,layer_3_1[999:992]} - {1'b0, layer_2_1[999:992]};
      btm_1[1] = {1'b0,layer_3_1[1007:1000]} - {1'b0, layer_2_1[1007:1000]};
      btm_1[2] = {1'b0,layer_3_1[1015:1008]} - {1'b0, layer_2_1[1015:1008]};
      btm_2[0] = {1'b0,layer_3_2[999:992]} - {1'b0, layer_2_2[999:992]};
      btm_2[1] = {1'b0,layer_3_2[1007:1000]} - {1'b0, layer_2_2[1007:1000]};
      btm_2[2] = {1'b0,layer_3_2[1015:1008]} - {1'b0, layer_2_2[1015:1008]};
    end
    'd126: begin
      top_0[0] = {1'b0,layer_1_0[1007:1000]} - {1'b0, layer_0_0[1007:1000]};
      top_0[1] = {1'b0,layer_1_0[1015:1008]} - {1'b0, layer_0_0[1015:1008]};
      top_0[2] = {1'b0,layer_1_0[1023:1016]} - {1'b0, layer_0_0[1023:1016]};
      top_1[0] = {1'b0,layer_1_1[1007:1000]} - {1'b0, layer_0_1[1007:1000]};
      top_1[1] = {1'b0,layer_1_1[1015:1008]} - {1'b0, layer_0_1[1015:1008]};
      top_1[2] = {1'b0,layer_1_1[1023:1016]} - {1'b0, layer_0_1[1023:1016]};
      top_2[0] = {1'b0,layer_1_2[1007:1000]} - {1'b0, layer_0_2[1007:1000]};
      top_2[1] = {1'b0,layer_1_2[1015:1008]} - {1'b0, layer_0_2[1015:1008]};
      top_2[2] = {1'b0,layer_1_2[1023:1016]} - {1'b0, layer_0_2[1023:1016]};
      mid_0[0] = {1'b0,layer_2_0[1007:1000]} - {1'b0, layer_1_0[1007:1000]};
      mid_0[1] = {1'b0,layer_2_0[1015:1008]} - {1'b0, layer_1_0[1015:1008]};
      mid_0[2] = {1'b0,layer_2_0[1023:1016]} - {1'b0, layer_1_0[1023:1016]};
      mid_1[0] = {1'b0,layer_2_1[1007:1000]} - {1'b0, layer_1_1[1007:1000]};
      mid_1[1] = {1'b0,layer_2_1[1015:1008]} - {1'b0, layer_1_1[1015:1008]};
      mid_1[2] = {1'b0,layer_2_1[1023:1016]} - {1'b0, layer_1_1[1023:1016]};
      mid_2[0] = {1'b0,layer_2_2[1007:1000]} - {1'b0, layer_1_2[1007:1000]};
      mid_2[1] = {1'b0,layer_2_2[1015:1008]} - {1'b0, layer_1_2[1015:1008]};
      mid_2[2] = {1'b0,layer_2_2[1023:1016]} - {1'b0, layer_1_2[1023:1016]};
      btm_0[0] = {1'b0,layer_3_0[1007:1000]} - {1'b0, layer_2_0[1007:1000]};
      btm_0[1] = {1'b0,layer_3_0[1015:1008]} - {1'b0, layer_2_0[1015:1008]};
      btm_0[2] = {1'b0,layer_3_0[1023:1016]} - {1'b0, layer_2_0[1023:1016]};
      btm_1[0] = {1'b0,layer_3_1[1007:1000]} - {1'b0, layer_2_1[1007:1000]};
      btm_1[1] = {1'b0,layer_3_1[1015:1008]} - {1'b0, layer_2_1[1015:1008]};
      btm_1[2] = {1'b0,layer_3_1[1023:1016]} - {1'b0, layer_2_1[1023:1016]};
      btm_2[0] = {1'b0,layer_3_2[1007:1000]} - {1'b0, layer_2_2[1007:1000]};
      btm_2[1] = {1'b0,layer_3_2[1015:1008]} - {1'b0, layer_2_2[1015:1008]};
      btm_2[2] = {1'b0,layer_3_2[1023:1016]} - {1'b0, layer_2_2[1023:1016]};
    end
    'd127: begin
      top_0[0] = {1'b0,layer_1_0[1015:1008]} - {1'b0, layer_0_0[1015:1008]};
      top_0[1] = {1'b0,layer_1_0[1023:1016]} - {1'b0, layer_0_0[1023:1016]};
      top_0[2] = {1'b0,layer_1_0[1031:1024]} - {1'b0, layer_0_0[1031:1024]};
      top_1[0] = {1'b0,layer_1_1[1015:1008]} - {1'b0, layer_0_1[1015:1008]};
      top_1[1] = {1'b0,layer_1_1[1023:1016]} - {1'b0, layer_0_1[1023:1016]};
      top_1[2] = {1'b0,layer_1_1[1031:1024]} - {1'b0, layer_0_1[1031:1024]};
      top_2[0] = {1'b0,layer_1_2[1015:1008]} - {1'b0, layer_0_2[1015:1008]};
      top_2[1] = {1'b0,layer_1_2[1023:1016]} - {1'b0, layer_0_2[1023:1016]};
      top_2[2] = {1'b0,layer_1_2[1031:1024]} - {1'b0, layer_0_2[1031:1024]};
      mid_0[0] = {1'b0,layer_2_0[1015:1008]} - {1'b0, layer_1_0[1015:1008]};
      mid_0[1] = {1'b0,layer_2_0[1023:1016]} - {1'b0, layer_1_0[1023:1016]};
      mid_0[2] = {1'b0,layer_2_0[1031:1024]} - {1'b0, layer_1_0[1031:1024]};
      mid_1[0] = {1'b0,layer_2_1[1015:1008]} - {1'b0, layer_1_1[1015:1008]};
      mid_1[1] = {1'b0,layer_2_1[1023:1016]} - {1'b0, layer_1_1[1023:1016]};
      mid_1[2] = {1'b0,layer_2_1[1031:1024]} - {1'b0, layer_1_1[1031:1024]};
      mid_2[0] = {1'b0,layer_2_2[1015:1008]} - {1'b0, layer_1_2[1015:1008]};
      mid_2[1] = {1'b0,layer_2_2[1023:1016]} - {1'b0, layer_1_2[1023:1016]};
      mid_2[2] = {1'b0,layer_2_2[1031:1024]} - {1'b0, layer_1_2[1031:1024]};
      btm_0[0] = {1'b0,layer_3_0[1015:1008]} - {1'b0, layer_2_0[1015:1008]};
      btm_0[1] = {1'b0,layer_3_0[1023:1016]} - {1'b0, layer_2_0[1023:1016]};
      btm_0[2] = {1'b0,layer_3_0[1031:1024]} - {1'b0, layer_2_0[1031:1024]};
      btm_1[0] = {1'b0,layer_3_1[1015:1008]} - {1'b0, layer_2_1[1015:1008]};
      btm_1[1] = {1'b0,layer_3_1[1023:1016]} - {1'b0, layer_2_1[1023:1016]};
      btm_1[2] = {1'b0,layer_3_1[1031:1024]} - {1'b0, layer_2_1[1031:1024]};
      btm_2[0] = {1'b0,layer_3_2[1015:1008]} - {1'b0, layer_2_2[1015:1008]};
      btm_2[1] = {1'b0,layer_3_2[1023:1016]} - {1'b0, layer_2_2[1023:1016]};
      btm_2[2] = {1'b0,layer_3_2[1031:1024]} - {1'b0, layer_2_2[1031:1024]};
    end
    'd128: begin
      top_0[0] = {1'b0,layer_1_0[1023:1016]} - {1'b0, layer_0_0[1023:1016]};
      top_0[1] = {1'b0,layer_1_0[1031:1024]} - {1'b0, layer_0_0[1031:1024]};
      top_0[2] = {1'b0,layer_1_0[1039:1032]} - {1'b0, layer_0_0[1039:1032]};
      top_1[0] = {1'b0,layer_1_1[1023:1016]} - {1'b0, layer_0_1[1023:1016]};
      top_1[1] = {1'b0,layer_1_1[1031:1024]} - {1'b0, layer_0_1[1031:1024]};
      top_1[2] = {1'b0,layer_1_1[1039:1032]} - {1'b0, layer_0_1[1039:1032]};
      top_2[0] = {1'b0,layer_1_2[1023:1016]} - {1'b0, layer_0_2[1023:1016]};
      top_2[1] = {1'b0,layer_1_2[1031:1024]} - {1'b0, layer_0_2[1031:1024]};
      top_2[2] = {1'b0,layer_1_2[1039:1032]} - {1'b0, layer_0_2[1039:1032]};
      mid_0[0] = {1'b0,layer_2_0[1023:1016]} - {1'b0, layer_1_0[1023:1016]};
      mid_0[1] = {1'b0,layer_2_0[1031:1024]} - {1'b0, layer_1_0[1031:1024]};
      mid_0[2] = {1'b0,layer_2_0[1039:1032]} - {1'b0, layer_1_0[1039:1032]};
      mid_1[0] = {1'b0,layer_2_1[1023:1016]} - {1'b0, layer_1_1[1023:1016]};
      mid_1[1] = {1'b0,layer_2_1[1031:1024]} - {1'b0, layer_1_1[1031:1024]};
      mid_1[2] = {1'b0,layer_2_1[1039:1032]} - {1'b0, layer_1_1[1039:1032]};
      mid_2[0] = {1'b0,layer_2_2[1023:1016]} - {1'b0, layer_1_2[1023:1016]};
      mid_2[1] = {1'b0,layer_2_2[1031:1024]} - {1'b0, layer_1_2[1031:1024]};
      mid_2[2] = {1'b0,layer_2_2[1039:1032]} - {1'b0, layer_1_2[1039:1032]};
      btm_0[0] = {1'b0,layer_3_0[1023:1016]} - {1'b0, layer_2_0[1023:1016]};
      btm_0[1] = {1'b0,layer_3_0[1031:1024]} - {1'b0, layer_2_0[1031:1024]};
      btm_0[2] = {1'b0,layer_3_0[1039:1032]} - {1'b0, layer_2_0[1039:1032]};
      btm_1[0] = {1'b0,layer_3_1[1023:1016]} - {1'b0, layer_2_1[1023:1016]};
      btm_1[1] = {1'b0,layer_3_1[1031:1024]} - {1'b0, layer_2_1[1031:1024]};
      btm_1[2] = {1'b0,layer_3_1[1039:1032]} - {1'b0, layer_2_1[1039:1032]};
      btm_2[0] = {1'b0,layer_3_2[1023:1016]} - {1'b0, layer_2_2[1023:1016]};
      btm_2[1] = {1'b0,layer_3_2[1031:1024]} - {1'b0, layer_2_2[1031:1024]};
      btm_2[2] = {1'b0,layer_3_2[1039:1032]} - {1'b0, layer_2_2[1039:1032]};
    end
    'd129: begin
      top_0[0] = {1'b0,layer_1_0[1031:1024]} - {1'b0, layer_0_0[1031:1024]};
      top_0[1] = {1'b0,layer_1_0[1039:1032]} - {1'b0, layer_0_0[1039:1032]};
      top_0[2] = {1'b0,layer_1_0[1047:1040]} - {1'b0, layer_0_0[1047:1040]};
      top_1[0] = {1'b0,layer_1_1[1031:1024]} - {1'b0, layer_0_1[1031:1024]};
      top_1[1] = {1'b0,layer_1_1[1039:1032]} - {1'b0, layer_0_1[1039:1032]};
      top_1[2] = {1'b0,layer_1_1[1047:1040]} - {1'b0, layer_0_1[1047:1040]};
      top_2[0] = {1'b0,layer_1_2[1031:1024]} - {1'b0, layer_0_2[1031:1024]};
      top_2[1] = {1'b0,layer_1_2[1039:1032]} - {1'b0, layer_0_2[1039:1032]};
      top_2[2] = {1'b0,layer_1_2[1047:1040]} - {1'b0, layer_0_2[1047:1040]};
      mid_0[0] = {1'b0,layer_2_0[1031:1024]} - {1'b0, layer_1_0[1031:1024]};
      mid_0[1] = {1'b0,layer_2_0[1039:1032]} - {1'b0, layer_1_0[1039:1032]};
      mid_0[2] = {1'b0,layer_2_0[1047:1040]} - {1'b0, layer_1_0[1047:1040]};
      mid_1[0] = {1'b0,layer_2_1[1031:1024]} - {1'b0, layer_1_1[1031:1024]};
      mid_1[1] = {1'b0,layer_2_1[1039:1032]} - {1'b0, layer_1_1[1039:1032]};
      mid_1[2] = {1'b0,layer_2_1[1047:1040]} - {1'b0, layer_1_1[1047:1040]};
      mid_2[0] = {1'b0,layer_2_2[1031:1024]} - {1'b0, layer_1_2[1031:1024]};
      mid_2[1] = {1'b0,layer_2_2[1039:1032]} - {1'b0, layer_1_2[1039:1032]};
      mid_2[2] = {1'b0,layer_2_2[1047:1040]} - {1'b0, layer_1_2[1047:1040]};
      btm_0[0] = {1'b0,layer_3_0[1031:1024]} - {1'b0, layer_2_0[1031:1024]};
      btm_0[1] = {1'b0,layer_3_0[1039:1032]} - {1'b0, layer_2_0[1039:1032]};
      btm_0[2] = {1'b0,layer_3_0[1047:1040]} - {1'b0, layer_2_0[1047:1040]};
      btm_1[0] = {1'b0,layer_3_1[1031:1024]} - {1'b0, layer_2_1[1031:1024]};
      btm_1[1] = {1'b0,layer_3_1[1039:1032]} - {1'b0, layer_2_1[1039:1032]};
      btm_1[2] = {1'b0,layer_3_1[1047:1040]} - {1'b0, layer_2_1[1047:1040]};
      btm_2[0] = {1'b0,layer_3_2[1031:1024]} - {1'b0, layer_2_2[1031:1024]};
      btm_2[1] = {1'b0,layer_3_2[1039:1032]} - {1'b0, layer_2_2[1039:1032]};
      btm_2[2] = {1'b0,layer_3_2[1047:1040]} - {1'b0, layer_2_2[1047:1040]};
    end
    'd130: begin
      top_0[0] = {1'b0,layer_1_0[1039:1032]} - {1'b0, layer_0_0[1039:1032]};
      top_0[1] = {1'b0,layer_1_0[1047:1040]} - {1'b0, layer_0_0[1047:1040]};
      top_0[2] = {1'b0,layer_1_0[1055:1048]} - {1'b0, layer_0_0[1055:1048]};
      top_1[0] = {1'b0,layer_1_1[1039:1032]} - {1'b0, layer_0_1[1039:1032]};
      top_1[1] = {1'b0,layer_1_1[1047:1040]} - {1'b0, layer_0_1[1047:1040]};
      top_1[2] = {1'b0,layer_1_1[1055:1048]} - {1'b0, layer_0_1[1055:1048]};
      top_2[0] = {1'b0,layer_1_2[1039:1032]} - {1'b0, layer_0_2[1039:1032]};
      top_2[1] = {1'b0,layer_1_2[1047:1040]} - {1'b0, layer_0_2[1047:1040]};
      top_2[2] = {1'b0,layer_1_2[1055:1048]} - {1'b0, layer_0_2[1055:1048]};
      mid_0[0] = {1'b0,layer_2_0[1039:1032]} - {1'b0, layer_1_0[1039:1032]};
      mid_0[1] = {1'b0,layer_2_0[1047:1040]} - {1'b0, layer_1_0[1047:1040]};
      mid_0[2] = {1'b0,layer_2_0[1055:1048]} - {1'b0, layer_1_0[1055:1048]};
      mid_1[0] = {1'b0,layer_2_1[1039:1032]} - {1'b0, layer_1_1[1039:1032]};
      mid_1[1] = {1'b0,layer_2_1[1047:1040]} - {1'b0, layer_1_1[1047:1040]};
      mid_1[2] = {1'b0,layer_2_1[1055:1048]} - {1'b0, layer_1_1[1055:1048]};
      mid_2[0] = {1'b0,layer_2_2[1039:1032]} - {1'b0, layer_1_2[1039:1032]};
      mid_2[1] = {1'b0,layer_2_2[1047:1040]} - {1'b0, layer_1_2[1047:1040]};
      mid_2[2] = {1'b0,layer_2_2[1055:1048]} - {1'b0, layer_1_2[1055:1048]};
      btm_0[0] = {1'b0,layer_3_0[1039:1032]} - {1'b0, layer_2_0[1039:1032]};
      btm_0[1] = {1'b0,layer_3_0[1047:1040]} - {1'b0, layer_2_0[1047:1040]};
      btm_0[2] = {1'b0,layer_3_0[1055:1048]} - {1'b0, layer_2_0[1055:1048]};
      btm_1[0] = {1'b0,layer_3_1[1039:1032]} - {1'b0, layer_2_1[1039:1032]};
      btm_1[1] = {1'b0,layer_3_1[1047:1040]} - {1'b0, layer_2_1[1047:1040]};
      btm_1[2] = {1'b0,layer_3_1[1055:1048]} - {1'b0, layer_2_1[1055:1048]};
      btm_2[0] = {1'b0,layer_3_2[1039:1032]} - {1'b0, layer_2_2[1039:1032]};
      btm_2[1] = {1'b0,layer_3_2[1047:1040]} - {1'b0, layer_2_2[1047:1040]};
      btm_2[2] = {1'b0,layer_3_2[1055:1048]} - {1'b0, layer_2_2[1055:1048]};
    end
    'd131: begin
      top_0[0] = {1'b0,layer_1_0[1047:1040]} - {1'b0, layer_0_0[1047:1040]};
      top_0[1] = {1'b0,layer_1_0[1055:1048]} - {1'b0, layer_0_0[1055:1048]};
      top_0[2] = {1'b0,layer_1_0[1063:1056]} - {1'b0, layer_0_0[1063:1056]};
      top_1[0] = {1'b0,layer_1_1[1047:1040]} - {1'b0, layer_0_1[1047:1040]};
      top_1[1] = {1'b0,layer_1_1[1055:1048]} - {1'b0, layer_0_1[1055:1048]};
      top_1[2] = {1'b0,layer_1_1[1063:1056]} - {1'b0, layer_0_1[1063:1056]};
      top_2[0] = {1'b0,layer_1_2[1047:1040]} - {1'b0, layer_0_2[1047:1040]};
      top_2[1] = {1'b0,layer_1_2[1055:1048]} - {1'b0, layer_0_2[1055:1048]};
      top_2[2] = {1'b0,layer_1_2[1063:1056]} - {1'b0, layer_0_2[1063:1056]};
      mid_0[0] = {1'b0,layer_2_0[1047:1040]} - {1'b0, layer_1_0[1047:1040]};
      mid_0[1] = {1'b0,layer_2_0[1055:1048]} - {1'b0, layer_1_0[1055:1048]};
      mid_0[2] = {1'b0,layer_2_0[1063:1056]} - {1'b0, layer_1_0[1063:1056]};
      mid_1[0] = {1'b0,layer_2_1[1047:1040]} - {1'b0, layer_1_1[1047:1040]};
      mid_1[1] = {1'b0,layer_2_1[1055:1048]} - {1'b0, layer_1_1[1055:1048]};
      mid_1[2] = {1'b0,layer_2_1[1063:1056]} - {1'b0, layer_1_1[1063:1056]};
      mid_2[0] = {1'b0,layer_2_2[1047:1040]} - {1'b0, layer_1_2[1047:1040]};
      mid_2[1] = {1'b0,layer_2_2[1055:1048]} - {1'b0, layer_1_2[1055:1048]};
      mid_2[2] = {1'b0,layer_2_2[1063:1056]} - {1'b0, layer_1_2[1063:1056]};
      btm_0[0] = {1'b0,layer_3_0[1047:1040]} - {1'b0, layer_2_0[1047:1040]};
      btm_0[1] = {1'b0,layer_3_0[1055:1048]} - {1'b0, layer_2_0[1055:1048]};
      btm_0[2] = {1'b0,layer_3_0[1063:1056]} - {1'b0, layer_2_0[1063:1056]};
      btm_1[0] = {1'b0,layer_3_1[1047:1040]} - {1'b0, layer_2_1[1047:1040]};
      btm_1[1] = {1'b0,layer_3_1[1055:1048]} - {1'b0, layer_2_1[1055:1048]};
      btm_1[2] = {1'b0,layer_3_1[1063:1056]} - {1'b0, layer_2_1[1063:1056]};
      btm_2[0] = {1'b0,layer_3_2[1047:1040]} - {1'b0, layer_2_2[1047:1040]};
      btm_2[1] = {1'b0,layer_3_2[1055:1048]} - {1'b0, layer_2_2[1055:1048]};
      btm_2[2] = {1'b0,layer_3_2[1063:1056]} - {1'b0, layer_2_2[1063:1056]};
    end
    'd132: begin
      top_0[0] = {1'b0,layer_1_0[1055:1048]} - {1'b0, layer_0_0[1055:1048]};
      top_0[1] = {1'b0,layer_1_0[1063:1056]} - {1'b0, layer_0_0[1063:1056]};
      top_0[2] = {1'b0,layer_1_0[1071:1064]} - {1'b0, layer_0_0[1071:1064]};
      top_1[0] = {1'b0,layer_1_1[1055:1048]} - {1'b0, layer_0_1[1055:1048]};
      top_1[1] = {1'b0,layer_1_1[1063:1056]} - {1'b0, layer_0_1[1063:1056]};
      top_1[2] = {1'b0,layer_1_1[1071:1064]} - {1'b0, layer_0_1[1071:1064]};
      top_2[0] = {1'b0,layer_1_2[1055:1048]} - {1'b0, layer_0_2[1055:1048]};
      top_2[1] = {1'b0,layer_1_2[1063:1056]} - {1'b0, layer_0_2[1063:1056]};
      top_2[2] = {1'b0,layer_1_2[1071:1064]} - {1'b0, layer_0_2[1071:1064]};
      mid_0[0] = {1'b0,layer_2_0[1055:1048]} - {1'b0, layer_1_0[1055:1048]};
      mid_0[1] = {1'b0,layer_2_0[1063:1056]} - {1'b0, layer_1_0[1063:1056]};
      mid_0[2] = {1'b0,layer_2_0[1071:1064]} - {1'b0, layer_1_0[1071:1064]};
      mid_1[0] = {1'b0,layer_2_1[1055:1048]} - {1'b0, layer_1_1[1055:1048]};
      mid_1[1] = {1'b0,layer_2_1[1063:1056]} - {1'b0, layer_1_1[1063:1056]};
      mid_1[2] = {1'b0,layer_2_1[1071:1064]} - {1'b0, layer_1_1[1071:1064]};
      mid_2[0] = {1'b0,layer_2_2[1055:1048]} - {1'b0, layer_1_2[1055:1048]};
      mid_2[1] = {1'b0,layer_2_2[1063:1056]} - {1'b0, layer_1_2[1063:1056]};
      mid_2[2] = {1'b0,layer_2_2[1071:1064]} - {1'b0, layer_1_2[1071:1064]};
      btm_0[0] = {1'b0,layer_3_0[1055:1048]} - {1'b0, layer_2_0[1055:1048]};
      btm_0[1] = {1'b0,layer_3_0[1063:1056]} - {1'b0, layer_2_0[1063:1056]};
      btm_0[2] = {1'b0,layer_3_0[1071:1064]} - {1'b0, layer_2_0[1071:1064]};
      btm_1[0] = {1'b0,layer_3_1[1055:1048]} - {1'b0, layer_2_1[1055:1048]};
      btm_1[1] = {1'b0,layer_3_1[1063:1056]} - {1'b0, layer_2_1[1063:1056]};
      btm_1[2] = {1'b0,layer_3_1[1071:1064]} - {1'b0, layer_2_1[1071:1064]};
      btm_2[0] = {1'b0,layer_3_2[1055:1048]} - {1'b0, layer_2_2[1055:1048]};
      btm_2[1] = {1'b0,layer_3_2[1063:1056]} - {1'b0, layer_2_2[1063:1056]};
      btm_2[2] = {1'b0,layer_3_2[1071:1064]} - {1'b0, layer_2_2[1071:1064]};
    end
    'd133: begin
      top_0[0] = {1'b0,layer_1_0[1063:1056]} - {1'b0, layer_0_0[1063:1056]};
      top_0[1] = {1'b0,layer_1_0[1071:1064]} - {1'b0, layer_0_0[1071:1064]};
      top_0[2] = {1'b0,layer_1_0[1079:1072]} - {1'b0, layer_0_0[1079:1072]};
      top_1[0] = {1'b0,layer_1_1[1063:1056]} - {1'b0, layer_0_1[1063:1056]};
      top_1[1] = {1'b0,layer_1_1[1071:1064]} - {1'b0, layer_0_1[1071:1064]};
      top_1[2] = {1'b0,layer_1_1[1079:1072]} - {1'b0, layer_0_1[1079:1072]};
      top_2[0] = {1'b0,layer_1_2[1063:1056]} - {1'b0, layer_0_2[1063:1056]};
      top_2[1] = {1'b0,layer_1_2[1071:1064]} - {1'b0, layer_0_2[1071:1064]};
      top_2[2] = {1'b0,layer_1_2[1079:1072]} - {1'b0, layer_0_2[1079:1072]};
      mid_0[0] = {1'b0,layer_2_0[1063:1056]} - {1'b0, layer_1_0[1063:1056]};
      mid_0[1] = {1'b0,layer_2_0[1071:1064]} - {1'b0, layer_1_0[1071:1064]};
      mid_0[2] = {1'b0,layer_2_0[1079:1072]} - {1'b0, layer_1_0[1079:1072]};
      mid_1[0] = {1'b0,layer_2_1[1063:1056]} - {1'b0, layer_1_1[1063:1056]};
      mid_1[1] = {1'b0,layer_2_1[1071:1064]} - {1'b0, layer_1_1[1071:1064]};
      mid_1[2] = {1'b0,layer_2_1[1079:1072]} - {1'b0, layer_1_1[1079:1072]};
      mid_2[0] = {1'b0,layer_2_2[1063:1056]} - {1'b0, layer_1_2[1063:1056]};
      mid_2[1] = {1'b0,layer_2_2[1071:1064]} - {1'b0, layer_1_2[1071:1064]};
      mid_2[2] = {1'b0,layer_2_2[1079:1072]} - {1'b0, layer_1_2[1079:1072]};
      btm_0[0] = {1'b0,layer_3_0[1063:1056]} - {1'b0, layer_2_0[1063:1056]};
      btm_0[1] = {1'b0,layer_3_0[1071:1064]} - {1'b0, layer_2_0[1071:1064]};
      btm_0[2] = {1'b0,layer_3_0[1079:1072]} - {1'b0, layer_2_0[1079:1072]};
      btm_1[0] = {1'b0,layer_3_1[1063:1056]} - {1'b0, layer_2_1[1063:1056]};
      btm_1[1] = {1'b0,layer_3_1[1071:1064]} - {1'b0, layer_2_1[1071:1064]};
      btm_1[2] = {1'b0,layer_3_1[1079:1072]} - {1'b0, layer_2_1[1079:1072]};
      btm_2[0] = {1'b0,layer_3_2[1063:1056]} - {1'b0, layer_2_2[1063:1056]};
      btm_2[1] = {1'b0,layer_3_2[1071:1064]} - {1'b0, layer_2_2[1071:1064]};
      btm_2[2] = {1'b0,layer_3_2[1079:1072]} - {1'b0, layer_2_2[1079:1072]};
    end
    'd134: begin
      top_0[0] = {1'b0,layer_1_0[1071:1064]} - {1'b0, layer_0_0[1071:1064]};
      top_0[1] = {1'b0,layer_1_0[1079:1072]} - {1'b0, layer_0_0[1079:1072]};
      top_0[2] = {1'b0,layer_1_0[1087:1080]} - {1'b0, layer_0_0[1087:1080]};
      top_1[0] = {1'b0,layer_1_1[1071:1064]} - {1'b0, layer_0_1[1071:1064]};
      top_1[1] = {1'b0,layer_1_1[1079:1072]} - {1'b0, layer_0_1[1079:1072]};
      top_1[2] = {1'b0,layer_1_1[1087:1080]} - {1'b0, layer_0_1[1087:1080]};
      top_2[0] = {1'b0,layer_1_2[1071:1064]} - {1'b0, layer_0_2[1071:1064]};
      top_2[1] = {1'b0,layer_1_2[1079:1072]} - {1'b0, layer_0_2[1079:1072]};
      top_2[2] = {1'b0,layer_1_2[1087:1080]} - {1'b0, layer_0_2[1087:1080]};
      mid_0[0] = {1'b0,layer_2_0[1071:1064]} - {1'b0, layer_1_0[1071:1064]};
      mid_0[1] = {1'b0,layer_2_0[1079:1072]} - {1'b0, layer_1_0[1079:1072]};
      mid_0[2] = {1'b0,layer_2_0[1087:1080]} - {1'b0, layer_1_0[1087:1080]};
      mid_1[0] = {1'b0,layer_2_1[1071:1064]} - {1'b0, layer_1_1[1071:1064]};
      mid_1[1] = {1'b0,layer_2_1[1079:1072]} - {1'b0, layer_1_1[1079:1072]};
      mid_1[2] = {1'b0,layer_2_1[1087:1080]} - {1'b0, layer_1_1[1087:1080]};
      mid_2[0] = {1'b0,layer_2_2[1071:1064]} - {1'b0, layer_1_2[1071:1064]};
      mid_2[1] = {1'b0,layer_2_2[1079:1072]} - {1'b0, layer_1_2[1079:1072]};
      mid_2[2] = {1'b0,layer_2_2[1087:1080]} - {1'b0, layer_1_2[1087:1080]};
      btm_0[0] = {1'b0,layer_3_0[1071:1064]} - {1'b0, layer_2_0[1071:1064]};
      btm_0[1] = {1'b0,layer_3_0[1079:1072]} - {1'b0, layer_2_0[1079:1072]};
      btm_0[2] = {1'b0,layer_3_0[1087:1080]} - {1'b0, layer_2_0[1087:1080]};
      btm_1[0] = {1'b0,layer_3_1[1071:1064]} - {1'b0, layer_2_1[1071:1064]};
      btm_1[1] = {1'b0,layer_3_1[1079:1072]} - {1'b0, layer_2_1[1079:1072]};
      btm_1[2] = {1'b0,layer_3_1[1087:1080]} - {1'b0, layer_2_1[1087:1080]};
      btm_2[0] = {1'b0,layer_3_2[1071:1064]} - {1'b0, layer_2_2[1071:1064]};
      btm_2[1] = {1'b0,layer_3_2[1079:1072]} - {1'b0, layer_2_2[1079:1072]};
      btm_2[2] = {1'b0,layer_3_2[1087:1080]} - {1'b0, layer_2_2[1087:1080]};
    end
    'd135: begin
      top_0[0] = {1'b0,layer_1_0[1079:1072]} - {1'b0, layer_0_0[1079:1072]};
      top_0[1] = {1'b0,layer_1_0[1087:1080]} - {1'b0, layer_0_0[1087:1080]};
      top_0[2] = {1'b0,layer_1_0[1095:1088]} - {1'b0, layer_0_0[1095:1088]};
      top_1[0] = {1'b0,layer_1_1[1079:1072]} - {1'b0, layer_0_1[1079:1072]};
      top_1[1] = {1'b0,layer_1_1[1087:1080]} - {1'b0, layer_0_1[1087:1080]};
      top_1[2] = {1'b0,layer_1_1[1095:1088]} - {1'b0, layer_0_1[1095:1088]};
      top_2[0] = {1'b0,layer_1_2[1079:1072]} - {1'b0, layer_0_2[1079:1072]};
      top_2[1] = {1'b0,layer_1_2[1087:1080]} - {1'b0, layer_0_2[1087:1080]};
      top_2[2] = {1'b0,layer_1_2[1095:1088]} - {1'b0, layer_0_2[1095:1088]};
      mid_0[0] = {1'b0,layer_2_0[1079:1072]} - {1'b0, layer_1_0[1079:1072]};
      mid_0[1] = {1'b0,layer_2_0[1087:1080]} - {1'b0, layer_1_0[1087:1080]};
      mid_0[2] = {1'b0,layer_2_0[1095:1088]} - {1'b0, layer_1_0[1095:1088]};
      mid_1[0] = {1'b0,layer_2_1[1079:1072]} - {1'b0, layer_1_1[1079:1072]};
      mid_1[1] = {1'b0,layer_2_1[1087:1080]} - {1'b0, layer_1_1[1087:1080]};
      mid_1[2] = {1'b0,layer_2_1[1095:1088]} - {1'b0, layer_1_1[1095:1088]};
      mid_2[0] = {1'b0,layer_2_2[1079:1072]} - {1'b0, layer_1_2[1079:1072]};
      mid_2[1] = {1'b0,layer_2_2[1087:1080]} - {1'b0, layer_1_2[1087:1080]};
      mid_2[2] = {1'b0,layer_2_2[1095:1088]} - {1'b0, layer_1_2[1095:1088]};
      btm_0[0] = {1'b0,layer_3_0[1079:1072]} - {1'b0, layer_2_0[1079:1072]};
      btm_0[1] = {1'b0,layer_3_0[1087:1080]} - {1'b0, layer_2_0[1087:1080]};
      btm_0[2] = {1'b0,layer_3_0[1095:1088]} - {1'b0, layer_2_0[1095:1088]};
      btm_1[0] = {1'b0,layer_3_1[1079:1072]} - {1'b0, layer_2_1[1079:1072]};
      btm_1[1] = {1'b0,layer_3_1[1087:1080]} - {1'b0, layer_2_1[1087:1080]};
      btm_1[2] = {1'b0,layer_3_1[1095:1088]} - {1'b0, layer_2_1[1095:1088]};
      btm_2[0] = {1'b0,layer_3_2[1079:1072]} - {1'b0, layer_2_2[1079:1072]};
      btm_2[1] = {1'b0,layer_3_2[1087:1080]} - {1'b0, layer_2_2[1087:1080]};
      btm_2[2] = {1'b0,layer_3_2[1095:1088]} - {1'b0, layer_2_2[1095:1088]};
    end
    'd136: begin
      top_0[0] = {1'b0,layer_1_0[1087:1080]} - {1'b0, layer_0_0[1087:1080]};
      top_0[1] = {1'b0,layer_1_0[1095:1088]} - {1'b0, layer_0_0[1095:1088]};
      top_0[2] = {1'b0,layer_1_0[1103:1096]} - {1'b0, layer_0_0[1103:1096]};
      top_1[0] = {1'b0,layer_1_1[1087:1080]} - {1'b0, layer_0_1[1087:1080]};
      top_1[1] = {1'b0,layer_1_1[1095:1088]} - {1'b0, layer_0_1[1095:1088]};
      top_1[2] = {1'b0,layer_1_1[1103:1096]} - {1'b0, layer_0_1[1103:1096]};
      top_2[0] = {1'b0,layer_1_2[1087:1080]} - {1'b0, layer_0_2[1087:1080]};
      top_2[1] = {1'b0,layer_1_2[1095:1088]} - {1'b0, layer_0_2[1095:1088]};
      top_2[2] = {1'b0,layer_1_2[1103:1096]} - {1'b0, layer_0_2[1103:1096]};
      mid_0[0] = {1'b0,layer_2_0[1087:1080]} - {1'b0, layer_1_0[1087:1080]};
      mid_0[1] = {1'b0,layer_2_0[1095:1088]} - {1'b0, layer_1_0[1095:1088]};
      mid_0[2] = {1'b0,layer_2_0[1103:1096]} - {1'b0, layer_1_0[1103:1096]};
      mid_1[0] = {1'b0,layer_2_1[1087:1080]} - {1'b0, layer_1_1[1087:1080]};
      mid_1[1] = {1'b0,layer_2_1[1095:1088]} - {1'b0, layer_1_1[1095:1088]};
      mid_1[2] = {1'b0,layer_2_1[1103:1096]} - {1'b0, layer_1_1[1103:1096]};
      mid_2[0] = {1'b0,layer_2_2[1087:1080]} - {1'b0, layer_1_2[1087:1080]};
      mid_2[1] = {1'b0,layer_2_2[1095:1088]} - {1'b0, layer_1_2[1095:1088]};
      mid_2[2] = {1'b0,layer_2_2[1103:1096]} - {1'b0, layer_1_2[1103:1096]};
      btm_0[0] = {1'b0,layer_3_0[1087:1080]} - {1'b0, layer_2_0[1087:1080]};
      btm_0[1] = {1'b0,layer_3_0[1095:1088]} - {1'b0, layer_2_0[1095:1088]};
      btm_0[2] = {1'b0,layer_3_0[1103:1096]} - {1'b0, layer_2_0[1103:1096]};
      btm_1[0] = {1'b0,layer_3_1[1087:1080]} - {1'b0, layer_2_1[1087:1080]};
      btm_1[1] = {1'b0,layer_3_1[1095:1088]} - {1'b0, layer_2_1[1095:1088]};
      btm_1[2] = {1'b0,layer_3_1[1103:1096]} - {1'b0, layer_2_1[1103:1096]};
      btm_2[0] = {1'b0,layer_3_2[1087:1080]} - {1'b0, layer_2_2[1087:1080]};
      btm_2[1] = {1'b0,layer_3_2[1095:1088]} - {1'b0, layer_2_2[1095:1088]};
      btm_2[2] = {1'b0,layer_3_2[1103:1096]} - {1'b0, layer_2_2[1103:1096]};
    end
    'd137: begin
      top_0[0] = {1'b0,layer_1_0[1095:1088]} - {1'b0, layer_0_0[1095:1088]};
      top_0[1] = {1'b0,layer_1_0[1103:1096]} - {1'b0, layer_0_0[1103:1096]};
      top_0[2] = {1'b0,layer_1_0[1111:1104]} - {1'b0, layer_0_0[1111:1104]};
      top_1[0] = {1'b0,layer_1_1[1095:1088]} - {1'b0, layer_0_1[1095:1088]};
      top_1[1] = {1'b0,layer_1_1[1103:1096]} - {1'b0, layer_0_1[1103:1096]};
      top_1[2] = {1'b0,layer_1_1[1111:1104]} - {1'b0, layer_0_1[1111:1104]};
      top_2[0] = {1'b0,layer_1_2[1095:1088]} - {1'b0, layer_0_2[1095:1088]};
      top_2[1] = {1'b0,layer_1_2[1103:1096]} - {1'b0, layer_0_2[1103:1096]};
      top_2[2] = {1'b0,layer_1_2[1111:1104]} - {1'b0, layer_0_2[1111:1104]};
      mid_0[0] = {1'b0,layer_2_0[1095:1088]} - {1'b0, layer_1_0[1095:1088]};
      mid_0[1] = {1'b0,layer_2_0[1103:1096]} - {1'b0, layer_1_0[1103:1096]};
      mid_0[2] = {1'b0,layer_2_0[1111:1104]} - {1'b0, layer_1_0[1111:1104]};
      mid_1[0] = {1'b0,layer_2_1[1095:1088]} - {1'b0, layer_1_1[1095:1088]};
      mid_1[1] = {1'b0,layer_2_1[1103:1096]} - {1'b0, layer_1_1[1103:1096]};
      mid_1[2] = {1'b0,layer_2_1[1111:1104]} - {1'b0, layer_1_1[1111:1104]};
      mid_2[0] = {1'b0,layer_2_2[1095:1088]} - {1'b0, layer_1_2[1095:1088]};
      mid_2[1] = {1'b0,layer_2_2[1103:1096]} - {1'b0, layer_1_2[1103:1096]};
      mid_2[2] = {1'b0,layer_2_2[1111:1104]} - {1'b0, layer_1_2[1111:1104]};
      btm_0[0] = {1'b0,layer_3_0[1095:1088]} - {1'b0, layer_2_0[1095:1088]};
      btm_0[1] = {1'b0,layer_3_0[1103:1096]} - {1'b0, layer_2_0[1103:1096]};
      btm_0[2] = {1'b0,layer_3_0[1111:1104]} - {1'b0, layer_2_0[1111:1104]};
      btm_1[0] = {1'b0,layer_3_1[1095:1088]} - {1'b0, layer_2_1[1095:1088]};
      btm_1[1] = {1'b0,layer_3_1[1103:1096]} - {1'b0, layer_2_1[1103:1096]};
      btm_1[2] = {1'b0,layer_3_1[1111:1104]} - {1'b0, layer_2_1[1111:1104]};
      btm_2[0] = {1'b0,layer_3_2[1095:1088]} - {1'b0, layer_2_2[1095:1088]};
      btm_2[1] = {1'b0,layer_3_2[1103:1096]} - {1'b0, layer_2_2[1103:1096]};
      btm_2[2] = {1'b0,layer_3_2[1111:1104]} - {1'b0, layer_2_2[1111:1104]};
    end
    'd138: begin
      top_0[0] = {1'b0,layer_1_0[1103:1096]} - {1'b0, layer_0_0[1103:1096]};
      top_0[1] = {1'b0,layer_1_0[1111:1104]} - {1'b0, layer_0_0[1111:1104]};
      top_0[2] = {1'b0,layer_1_0[1119:1112]} - {1'b0, layer_0_0[1119:1112]};
      top_1[0] = {1'b0,layer_1_1[1103:1096]} - {1'b0, layer_0_1[1103:1096]};
      top_1[1] = {1'b0,layer_1_1[1111:1104]} - {1'b0, layer_0_1[1111:1104]};
      top_1[2] = {1'b0,layer_1_1[1119:1112]} - {1'b0, layer_0_1[1119:1112]};
      top_2[0] = {1'b0,layer_1_2[1103:1096]} - {1'b0, layer_0_2[1103:1096]};
      top_2[1] = {1'b0,layer_1_2[1111:1104]} - {1'b0, layer_0_2[1111:1104]};
      top_2[2] = {1'b0,layer_1_2[1119:1112]} - {1'b0, layer_0_2[1119:1112]};
      mid_0[0] = {1'b0,layer_2_0[1103:1096]} - {1'b0, layer_1_0[1103:1096]};
      mid_0[1] = {1'b0,layer_2_0[1111:1104]} - {1'b0, layer_1_0[1111:1104]};
      mid_0[2] = {1'b0,layer_2_0[1119:1112]} - {1'b0, layer_1_0[1119:1112]};
      mid_1[0] = {1'b0,layer_2_1[1103:1096]} - {1'b0, layer_1_1[1103:1096]};
      mid_1[1] = {1'b0,layer_2_1[1111:1104]} - {1'b0, layer_1_1[1111:1104]};
      mid_1[2] = {1'b0,layer_2_1[1119:1112]} - {1'b0, layer_1_1[1119:1112]};
      mid_2[0] = {1'b0,layer_2_2[1103:1096]} - {1'b0, layer_1_2[1103:1096]};
      mid_2[1] = {1'b0,layer_2_2[1111:1104]} - {1'b0, layer_1_2[1111:1104]};
      mid_2[2] = {1'b0,layer_2_2[1119:1112]} - {1'b0, layer_1_2[1119:1112]};
      btm_0[0] = {1'b0,layer_3_0[1103:1096]} - {1'b0, layer_2_0[1103:1096]};
      btm_0[1] = {1'b0,layer_3_0[1111:1104]} - {1'b0, layer_2_0[1111:1104]};
      btm_0[2] = {1'b0,layer_3_0[1119:1112]} - {1'b0, layer_2_0[1119:1112]};
      btm_1[0] = {1'b0,layer_3_1[1103:1096]} - {1'b0, layer_2_1[1103:1096]};
      btm_1[1] = {1'b0,layer_3_1[1111:1104]} - {1'b0, layer_2_1[1111:1104]};
      btm_1[2] = {1'b0,layer_3_1[1119:1112]} - {1'b0, layer_2_1[1119:1112]};
      btm_2[0] = {1'b0,layer_3_2[1103:1096]} - {1'b0, layer_2_2[1103:1096]};
      btm_2[1] = {1'b0,layer_3_2[1111:1104]} - {1'b0, layer_2_2[1111:1104]};
      btm_2[2] = {1'b0,layer_3_2[1119:1112]} - {1'b0, layer_2_2[1119:1112]};
    end
    'd139: begin
      top_0[0] = {1'b0,layer_1_0[1111:1104]} - {1'b0, layer_0_0[1111:1104]};
      top_0[1] = {1'b0,layer_1_0[1119:1112]} - {1'b0, layer_0_0[1119:1112]};
      top_0[2] = {1'b0,layer_1_0[1127:1120]} - {1'b0, layer_0_0[1127:1120]};
      top_1[0] = {1'b0,layer_1_1[1111:1104]} - {1'b0, layer_0_1[1111:1104]};
      top_1[1] = {1'b0,layer_1_1[1119:1112]} - {1'b0, layer_0_1[1119:1112]};
      top_1[2] = {1'b0,layer_1_1[1127:1120]} - {1'b0, layer_0_1[1127:1120]};
      top_2[0] = {1'b0,layer_1_2[1111:1104]} - {1'b0, layer_0_2[1111:1104]};
      top_2[1] = {1'b0,layer_1_2[1119:1112]} - {1'b0, layer_0_2[1119:1112]};
      top_2[2] = {1'b0,layer_1_2[1127:1120]} - {1'b0, layer_0_2[1127:1120]};
      mid_0[0] = {1'b0,layer_2_0[1111:1104]} - {1'b0, layer_1_0[1111:1104]};
      mid_0[1] = {1'b0,layer_2_0[1119:1112]} - {1'b0, layer_1_0[1119:1112]};
      mid_0[2] = {1'b0,layer_2_0[1127:1120]} - {1'b0, layer_1_0[1127:1120]};
      mid_1[0] = {1'b0,layer_2_1[1111:1104]} - {1'b0, layer_1_1[1111:1104]};
      mid_1[1] = {1'b0,layer_2_1[1119:1112]} - {1'b0, layer_1_1[1119:1112]};
      mid_1[2] = {1'b0,layer_2_1[1127:1120]} - {1'b0, layer_1_1[1127:1120]};
      mid_2[0] = {1'b0,layer_2_2[1111:1104]} - {1'b0, layer_1_2[1111:1104]};
      mid_2[1] = {1'b0,layer_2_2[1119:1112]} - {1'b0, layer_1_2[1119:1112]};
      mid_2[2] = {1'b0,layer_2_2[1127:1120]} - {1'b0, layer_1_2[1127:1120]};
      btm_0[0] = {1'b0,layer_3_0[1111:1104]} - {1'b0, layer_2_0[1111:1104]};
      btm_0[1] = {1'b0,layer_3_0[1119:1112]} - {1'b0, layer_2_0[1119:1112]};
      btm_0[2] = {1'b0,layer_3_0[1127:1120]} - {1'b0, layer_2_0[1127:1120]};
      btm_1[0] = {1'b0,layer_3_1[1111:1104]} - {1'b0, layer_2_1[1111:1104]};
      btm_1[1] = {1'b0,layer_3_1[1119:1112]} - {1'b0, layer_2_1[1119:1112]};
      btm_1[2] = {1'b0,layer_3_1[1127:1120]} - {1'b0, layer_2_1[1127:1120]};
      btm_2[0] = {1'b0,layer_3_2[1111:1104]} - {1'b0, layer_2_2[1111:1104]};
      btm_2[1] = {1'b0,layer_3_2[1119:1112]} - {1'b0, layer_2_2[1119:1112]};
      btm_2[2] = {1'b0,layer_3_2[1127:1120]} - {1'b0, layer_2_2[1127:1120]};
    end
    'd140: begin
      top_0[0] = {1'b0,layer_1_0[1119:1112]} - {1'b0, layer_0_0[1119:1112]};
      top_0[1] = {1'b0,layer_1_0[1127:1120]} - {1'b0, layer_0_0[1127:1120]};
      top_0[2] = {1'b0,layer_1_0[1135:1128]} - {1'b0, layer_0_0[1135:1128]};
      top_1[0] = {1'b0,layer_1_1[1119:1112]} - {1'b0, layer_0_1[1119:1112]};
      top_1[1] = {1'b0,layer_1_1[1127:1120]} - {1'b0, layer_0_1[1127:1120]};
      top_1[2] = {1'b0,layer_1_1[1135:1128]} - {1'b0, layer_0_1[1135:1128]};
      top_2[0] = {1'b0,layer_1_2[1119:1112]} - {1'b0, layer_0_2[1119:1112]};
      top_2[1] = {1'b0,layer_1_2[1127:1120]} - {1'b0, layer_0_2[1127:1120]};
      top_2[2] = {1'b0,layer_1_2[1135:1128]} - {1'b0, layer_0_2[1135:1128]};
      mid_0[0] = {1'b0,layer_2_0[1119:1112]} - {1'b0, layer_1_0[1119:1112]};
      mid_0[1] = {1'b0,layer_2_0[1127:1120]} - {1'b0, layer_1_0[1127:1120]};
      mid_0[2] = {1'b0,layer_2_0[1135:1128]} - {1'b0, layer_1_0[1135:1128]};
      mid_1[0] = {1'b0,layer_2_1[1119:1112]} - {1'b0, layer_1_1[1119:1112]};
      mid_1[1] = {1'b0,layer_2_1[1127:1120]} - {1'b0, layer_1_1[1127:1120]};
      mid_1[2] = {1'b0,layer_2_1[1135:1128]} - {1'b0, layer_1_1[1135:1128]};
      mid_2[0] = {1'b0,layer_2_2[1119:1112]} - {1'b0, layer_1_2[1119:1112]};
      mid_2[1] = {1'b0,layer_2_2[1127:1120]} - {1'b0, layer_1_2[1127:1120]};
      mid_2[2] = {1'b0,layer_2_2[1135:1128]} - {1'b0, layer_1_2[1135:1128]};
      btm_0[0] = {1'b0,layer_3_0[1119:1112]} - {1'b0, layer_2_0[1119:1112]};
      btm_0[1] = {1'b0,layer_3_0[1127:1120]} - {1'b0, layer_2_0[1127:1120]};
      btm_0[2] = {1'b0,layer_3_0[1135:1128]} - {1'b0, layer_2_0[1135:1128]};
      btm_1[0] = {1'b0,layer_3_1[1119:1112]} - {1'b0, layer_2_1[1119:1112]};
      btm_1[1] = {1'b0,layer_3_1[1127:1120]} - {1'b0, layer_2_1[1127:1120]};
      btm_1[2] = {1'b0,layer_3_1[1135:1128]} - {1'b0, layer_2_1[1135:1128]};
      btm_2[0] = {1'b0,layer_3_2[1119:1112]} - {1'b0, layer_2_2[1119:1112]};
      btm_2[1] = {1'b0,layer_3_2[1127:1120]} - {1'b0, layer_2_2[1127:1120]};
      btm_2[2] = {1'b0,layer_3_2[1135:1128]} - {1'b0, layer_2_2[1135:1128]};
    end
    'd141: begin
      top_0[0] = {1'b0,layer_1_0[1127:1120]} - {1'b0, layer_0_0[1127:1120]};
      top_0[1] = {1'b0,layer_1_0[1135:1128]} - {1'b0, layer_0_0[1135:1128]};
      top_0[2] = {1'b0,layer_1_0[1143:1136]} - {1'b0, layer_0_0[1143:1136]};
      top_1[0] = {1'b0,layer_1_1[1127:1120]} - {1'b0, layer_0_1[1127:1120]};
      top_1[1] = {1'b0,layer_1_1[1135:1128]} - {1'b0, layer_0_1[1135:1128]};
      top_1[2] = {1'b0,layer_1_1[1143:1136]} - {1'b0, layer_0_1[1143:1136]};
      top_2[0] = {1'b0,layer_1_2[1127:1120]} - {1'b0, layer_0_2[1127:1120]};
      top_2[1] = {1'b0,layer_1_2[1135:1128]} - {1'b0, layer_0_2[1135:1128]};
      top_2[2] = {1'b0,layer_1_2[1143:1136]} - {1'b0, layer_0_2[1143:1136]};
      mid_0[0] = {1'b0,layer_2_0[1127:1120]} - {1'b0, layer_1_0[1127:1120]};
      mid_0[1] = {1'b0,layer_2_0[1135:1128]} - {1'b0, layer_1_0[1135:1128]};
      mid_0[2] = {1'b0,layer_2_0[1143:1136]} - {1'b0, layer_1_0[1143:1136]};
      mid_1[0] = {1'b0,layer_2_1[1127:1120]} - {1'b0, layer_1_1[1127:1120]};
      mid_1[1] = {1'b0,layer_2_1[1135:1128]} - {1'b0, layer_1_1[1135:1128]};
      mid_1[2] = {1'b0,layer_2_1[1143:1136]} - {1'b0, layer_1_1[1143:1136]};
      mid_2[0] = {1'b0,layer_2_2[1127:1120]} - {1'b0, layer_1_2[1127:1120]};
      mid_2[1] = {1'b0,layer_2_2[1135:1128]} - {1'b0, layer_1_2[1135:1128]};
      mid_2[2] = {1'b0,layer_2_2[1143:1136]} - {1'b0, layer_1_2[1143:1136]};
      btm_0[0] = {1'b0,layer_3_0[1127:1120]} - {1'b0, layer_2_0[1127:1120]};
      btm_0[1] = {1'b0,layer_3_0[1135:1128]} - {1'b0, layer_2_0[1135:1128]};
      btm_0[2] = {1'b0,layer_3_0[1143:1136]} - {1'b0, layer_2_0[1143:1136]};
      btm_1[0] = {1'b0,layer_3_1[1127:1120]} - {1'b0, layer_2_1[1127:1120]};
      btm_1[1] = {1'b0,layer_3_1[1135:1128]} - {1'b0, layer_2_1[1135:1128]};
      btm_1[2] = {1'b0,layer_3_1[1143:1136]} - {1'b0, layer_2_1[1143:1136]};
      btm_2[0] = {1'b0,layer_3_2[1127:1120]} - {1'b0, layer_2_2[1127:1120]};
      btm_2[1] = {1'b0,layer_3_2[1135:1128]} - {1'b0, layer_2_2[1135:1128]};
      btm_2[2] = {1'b0,layer_3_2[1143:1136]} - {1'b0, layer_2_2[1143:1136]};
    end
    'd142: begin
      top_0[0] = {1'b0,layer_1_0[1135:1128]} - {1'b0, layer_0_0[1135:1128]};
      top_0[1] = {1'b0,layer_1_0[1143:1136]} - {1'b0, layer_0_0[1143:1136]};
      top_0[2] = {1'b0,layer_1_0[1151:1144]} - {1'b0, layer_0_0[1151:1144]};
      top_1[0] = {1'b0,layer_1_1[1135:1128]} - {1'b0, layer_0_1[1135:1128]};
      top_1[1] = {1'b0,layer_1_1[1143:1136]} - {1'b0, layer_0_1[1143:1136]};
      top_1[2] = {1'b0,layer_1_1[1151:1144]} - {1'b0, layer_0_1[1151:1144]};
      top_2[0] = {1'b0,layer_1_2[1135:1128]} - {1'b0, layer_0_2[1135:1128]};
      top_2[1] = {1'b0,layer_1_2[1143:1136]} - {1'b0, layer_0_2[1143:1136]};
      top_2[2] = {1'b0,layer_1_2[1151:1144]} - {1'b0, layer_0_2[1151:1144]};
      mid_0[0] = {1'b0,layer_2_0[1135:1128]} - {1'b0, layer_1_0[1135:1128]};
      mid_0[1] = {1'b0,layer_2_0[1143:1136]} - {1'b0, layer_1_0[1143:1136]};
      mid_0[2] = {1'b0,layer_2_0[1151:1144]} - {1'b0, layer_1_0[1151:1144]};
      mid_1[0] = {1'b0,layer_2_1[1135:1128]} - {1'b0, layer_1_1[1135:1128]};
      mid_1[1] = {1'b0,layer_2_1[1143:1136]} - {1'b0, layer_1_1[1143:1136]};
      mid_1[2] = {1'b0,layer_2_1[1151:1144]} - {1'b0, layer_1_1[1151:1144]};
      mid_2[0] = {1'b0,layer_2_2[1135:1128]} - {1'b0, layer_1_2[1135:1128]};
      mid_2[1] = {1'b0,layer_2_2[1143:1136]} - {1'b0, layer_1_2[1143:1136]};
      mid_2[2] = {1'b0,layer_2_2[1151:1144]} - {1'b0, layer_1_2[1151:1144]};
      btm_0[0] = {1'b0,layer_3_0[1135:1128]} - {1'b0, layer_2_0[1135:1128]};
      btm_0[1] = {1'b0,layer_3_0[1143:1136]} - {1'b0, layer_2_0[1143:1136]};
      btm_0[2] = {1'b0,layer_3_0[1151:1144]} - {1'b0, layer_2_0[1151:1144]};
      btm_1[0] = {1'b0,layer_3_1[1135:1128]} - {1'b0, layer_2_1[1135:1128]};
      btm_1[1] = {1'b0,layer_3_1[1143:1136]} - {1'b0, layer_2_1[1143:1136]};
      btm_1[2] = {1'b0,layer_3_1[1151:1144]} - {1'b0, layer_2_1[1151:1144]};
      btm_2[0] = {1'b0,layer_3_2[1135:1128]} - {1'b0, layer_2_2[1135:1128]};
      btm_2[1] = {1'b0,layer_3_2[1143:1136]} - {1'b0, layer_2_2[1143:1136]};
      btm_2[2] = {1'b0,layer_3_2[1151:1144]} - {1'b0, layer_2_2[1151:1144]};
    end
    'd143: begin
      top_0[0] = {1'b0,layer_1_0[1143:1136]} - {1'b0, layer_0_0[1143:1136]};
      top_0[1] = {1'b0,layer_1_0[1151:1144]} - {1'b0, layer_0_0[1151:1144]};
      top_0[2] = {1'b0,layer_1_0[1159:1152]} - {1'b0, layer_0_0[1159:1152]};
      top_1[0] = {1'b0,layer_1_1[1143:1136]} - {1'b0, layer_0_1[1143:1136]};
      top_1[1] = {1'b0,layer_1_1[1151:1144]} - {1'b0, layer_0_1[1151:1144]};
      top_1[2] = {1'b0,layer_1_1[1159:1152]} - {1'b0, layer_0_1[1159:1152]};
      top_2[0] = {1'b0,layer_1_2[1143:1136]} - {1'b0, layer_0_2[1143:1136]};
      top_2[1] = {1'b0,layer_1_2[1151:1144]} - {1'b0, layer_0_2[1151:1144]};
      top_2[2] = {1'b0,layer_1_2[1159:1152]} - {1'b0, layer_0_2[1159:1152]};
      mid_0[0] = {1'b0,layer_2_0[1143:1136]} - {1'b0, layer_1_0[1143:1136]};
      mid_0[1] = {1'b0,layer_2_0[1151:1144]} - {1'b0, layer_1_0[1151:1144]};
      mid_0[2] = {1'b0,layer_2_0[1159:1152]} - {1'b0, layer_1_0[1159:1152]};
      mid_1[0] = {1'b0,layer_2_1[1143:1136]} - {1'b0, layer_1_1[1143:1136]};
      mid_1[1] = {1'b0,layer_2_1[1151:1144]} - {1'b0, layer_1_1[1151:1144]};
      mid_1[2] = {1'b0,layer_2_1[1159:1152]} - {1'b0, layer_1_1[1159:1152]};
      mid_2[0] = {1'b0,layer_2_2[1143:1136]} - {1'b0, layer_1_2[1143:1136]};
      mid_2[1] = {1'b0,layer_2_2[1151:1144]} - {1'b0, layer_1_2[1151:1144]};
      mid_2[2] = {1'b0,layer_2_2[1159:1152]} - {1'b0, layer_1_2[1159:1152]};
      btm_0[0] = {1'b0,layer_3_0[1143:1136]} - {1'b0, layer_2_0[1143:1136]};
      btm_0[1] = {1'b0,layer_3_0[1151:1144]} - {1'b0, layer_2_0[1151:1144]};
      btm_0[2] = {1'b0,layer_3_0[1159:1152]} - {1'b0, layer_2_0[1159:1152]};
      btm_1[0] = {1'b0,layer_3_1[1143:1136]} - {1'b0, layer_2_1[1143:1136]};
      btm_1[1] = {1'b0,layer_3_1[1151:1144]} - {1'b0, layer_2_1[1151:1144]};
      btm_1[2] = {1'b0,layer_3_1[1159:1152]} - {1'b0, layer_2_1[1159:1152]};
      btm_2[0] = {1'b0,layer_3_2[1143:1136]} - {1'b0, layer_2_2[1143:1136]};
      btm_2[1] = {1'b0,layer_3_2[1151:1144]} - {1'b0, layer_2_2[1151:1144]};
      btm_2[2] = {1'b0,layer_3_2[1159:1152]} - {1'b0, layer_2_2[1159:1152]};
    end
    'd144: begin
      top_0[0] = {1'b0,layer_1_0[1151:1144]} - {1'b0, layer_0_0[1151:1144]};
      top_0[1] = {1'b0,layer_1_0[1159:1152]} - {1'b0, layer_0_0[1159:1152]};
      top_0[2] = {1'b0,layer_1_0[1167:1160]} - {1'b0, layer_0_0[1167:1160]};
      top_1[0] = {1'b0,layer_1_1[1151:1144]} - {1'b0, layer_0_1[1151:1144]};
      top_1[1] = {1'b0,layer_1_1[1159:1152]} - {1'b0, layer_0_1[1159:1152]};
      top_1[2] = {1'b0,layer_1_1[1167:1160]} - {1'b0, layer_0_1[1167:1160]};
      top_2[0] = {1'b0,layer_1_2[1151:1144]} - {1'b0, layer_0_2[1151:1144]};
      top_2[1] = {1'b0,layer_1_2[1159:1152]} - {1'b0, layer_0_2[1159:1152]};
      top_2[2] = {1'b0,layer_1_2[1167:1160]} - {1'b0, layer_0_2[1167:1160]};
      mid_0[0] = {1'b0,layer_2_0[1151:1144]} - {1'b0, layer_1_0[1151:1144]};
      mid_0[1] = {1'b0,layer_2_0[1159:1152]} - {1'b0, layer_1_0[1159:1152]};
      mid_0[2] = {1'b0,layer_2_0[1167:1160]} - {1'b0, layer_1_0[1167:1160]};
      mid_1[0] = {1'b0,layer_2_1[1151:1144]} - {1'b0, layer_1_1[1151:1144]};
      mid_1[1] = {1'b0,layer_2_1[1159:1152]} - {1'b0, layer_1_1[1159:1152]};
      mid_1[2] = {1'b0,layer_2_1[1167:1160]} - {1'b0, layer_1_1[1167:1160]};
      mid_2[0] = {1'b0,layer_2_2[1151:1144]} - {1'b0, layer_1_2[1151:1144]};
      mid_2[1] = {1'b0,layer_2_2[1159:1152]} - {1'b0, layer_1_2[1159:1152]};
      mid_2[2] = {1'b0,layer_2_2[1167:1160]} - {1'b0, layer_1_2[1167:1160]};
      btm_0[0] = {1'b0,layer_3_0[1151:1144]} - {1'b0, layer_2_0[1151:1144]};
      btm_0[1] = {1'b0,layer_3_0[1159:1152]} - {1'b0, layer_2_0[1159:1152]};
      btm_0[2] = {1'b0,layer_3_0[1167:1160]} - {1'b0, layer_2_0[1167:1160]};
      btm_1[0] = {1'b0,layer_3_1[1151:1144]} - {1'b0, layer_2_1[1151:1144]};
      btm_1[1] = {1'b0,layer_3_1[1159:1152]} - {1'b0, layer_2_1[1159:1152]};
      btm_1[2] = {1'b0,layer_3_1[1167:1160]} - {1'b0, layer_2_1[1167:1160]};
      btm_2[0] = {1'b0,layer_3_2[1151:1144]} - {1'b0, layer_2_2[1151:1144]};
      btm_2[1] = {1'b0,layer_3_2[1159:1152]} - {1'b0, layer_2_2[1159:1152]};
      btm_2[2] = {1'b0,layer_3_2[1167:1160]} - {1'b0, layer_2_2[1167:1160]};
    end
    'd145: begin
      top_0[0] = {1'b0,layer_1_0[1159:1152]} - {1'b0, layer_0_0[1159:1152]};
      top_0[1] = {1'b0,layer_1_0[1167:1160]} - {1'b0, layer_0_0[1167:1160]};
      top_0[2] = {1'b0,layer_1_0[1175:1168]} - {1'b0, layer_0_0[1175:1168]};
      top_1[0] = {1'b0,layer_1_1[1159:1152]} - {1'b0, layer_0_1[1159:1152]};
      top_1[1] = {1'b0,layer_1_1[1167:1160]} - {1'b0, layer_0_1[1167:1160]};
      top_1[2] = {1'b0,layer_1_1[1175:1168]} - {1'b0, layer_0_1[1175:1168]};
      top_2[0] = {1'b0,layer_1_2[1159:1152]} - {1'b0, layer_0_2[1159:1152]};
      top_2[1] = {1'b0,layer_1_2[1167:1160]} - {1'b0, layer_0_2[1167:1160]};
      top_2[2] = {1'b0,layer_1_2[1175:1168]} - {1'b0, layer_0_2[1175:1168]};
      mid_0[0] = {1'b0,layer_2_0[1159:1152]} - {1'b0, layer_1_0[1159:1152]};
      mid_0[1] = {1'b0,layer_2_0[1167:1160]} - {1'b0, layer_1_0[1167:1160]};
      mid_0[2] = {1'b0,layer_2_0[1175:1168]} - {1'b0, layer_1_0[1175:1168]};
      mid_1[0] = {1'b0,layer_2_1[1159:1152]} - {1'b0, layer_1_1[1159:1152]};
      mid_1[1] = {1'b0,layer_2_1[1167:1160]} - {1'b0, layer_1_1[1167:1160]};
      mid_1[2] = {1'b0,layer_2_1[1175:1168]} - {1'b0, layer_1_1[1175:1168]};
      mid_2[0] = {1'b0,layer_2_2[1159:1152]} - {1'b0, layer_1_2[1159:1152]};
      mid_2[1] = {1'b0,layer_2_2[1167:1160]} - {1'b0, layer_1_2[1167:1160]};
      mid_2[2] = {1'b0,layer_2_2[1175:1168]} - {1'b0, layer_1_2[1175:1168]};
      btm_0[0] = {1'b0,layer_3_0[1159:1152]} - {1'b0, layer_2_0[1159:1152]};
      btm_0[1] = {1'b0,layer_3_0[1167:1160]} - {1'b0, layer_2_0[1167:1160]};
      btm_0[2] = {1'b0,layer_3_0[1175:1168]} - {1'b0, layer_2_0[1175:1168]};
      btm_1[0] = {1'b0,layer_3_1[1159:1152]} - {1'b0, layer_2_1[1159:1152]};
      btm_1[1] = {1'b0,layer_3_1[1167:1160]} - {1'b0, layer_2_1[1167:1160]};
      btm_1[2] = {1'b0,layer_3_1[1175:1168]} - {1'b0, layer_2_1[1175:1168]};
      btm_2[0] = {1'b0,layer_3_2[1159:1152]} - {1'b0, layer_2_2[1159:1152]};
      btm_2[1] = {1'b0,layer_3_2[1167:1160]} - {1'b0, layer_2_2[1167:1160]};
      btm_2[2] = {1'b0,layer_3_2[1175:1168]} - {1'b0, layer_2_2[1175:1168]};
    end
    'd146: begin
      top_0[0] = {1'b0,layer_1_0[1167:1160]} - {1'b0, layer_0_0[1167:1160]};
      top_0[1] = {1'b0,layer_1_0[1175:1168]} - {1'b0, layer_0_0[1175:1168]};
      top_0[2] = {1'b0,layer_1_0[1183:1176]} - {1'b0, layer_0_0[1183:1176]};
      top_1[0] = {1'b0,layer_1_1[1167:1160]} - {1'b0, layer_0_1[1167:1160]};
      top_1[1] = {1'b0,layer_1_1[1175:1168]} - {1'b0, layer_0_1[1175:1168]};
      top_1[2] = {1'b0,layer_1_1[1183:1176]} - {1'b0, layer_0_1[1183:1176]};
      top_2[0] = {1'b0,layer_1_2[1167:1160]} - {1'b0, layer_0_2[1167:1160]};
      top_2[1] = {1'b0,layer_1_2[1175:1168]} - {1'b0, layer_0_2[1175:1168]};
      top_2[2] = {1'b0,layer_1_2[1183:1176]} - {1'b0, layer_0_2[1183:1176]};
      mid_0[0] = {1'b0,layer_2_0[1167:1160]} - {1'b0, layer_1_0[1167:1160]};
      mid_0[1] = {1'b0,layer_2_0[1175:1168]} - {1'b0, layer_1_0[1175:1168]};
      mid_0[2] = {1'b0,layer_2_0[1183:1176]} - {1'b0, layer_1_0[1183:1176]};
      mid_1[0] = {1'b0,layer_2_1[1167:1160]} - {1'b0, layer_1_1[1167:1160]};
      mid_1[1] = {1'b0,layer_2_1[1175:1168]} - {1'b0, layer_1_1[1175:1168]};
      mid_1[2] = {1'b0,layer_2_1[1183:1176]} - {1'b0, layer_1_1[1183:1176]};
      mid_2[0] = {1'b0,layer_2_2[1167:1160]} - {1'b0, layer_1_2[1167:1160]};
      mid_2[1] = {1'b0,layer_2_2[1175:1168]} - {1'b0, layer_1_2[1175:1168]};
      mid_2[2] = {1'b0,layer_2_2[1183:1176]} - {1'b0, layer_1_2[1183:1176]};
      btm_0[0] = {1'b0,layer_3_0[1167:1160]} - {1'b0, layer_2_0[1167:1160]};
      btm_0[1] = {1'b0,layer_3_0[1175:1168]} - {1'b0, layer_2_0[1175:1168]};
      btm_0[2] = {1'b0,layer_3_0[1183:1176]} - {1'b0, layer_2_0[1183:1176]};
      btm_1[0] = {1'b0,layer_3_1[1167:1160]} - {1'b0, layer_2_1[1167:1160]};
      btm_1[1] = {1'b0,layer_3_1[1175:1168]} - {1'b0, layer_2_1[1175:1168]};
      btm_1[2] = {1'b0,layer_3_1[1183:1176]} - {1'b0, layer_2_1[1183:1176]};
      btm_2[0] = {1'b0,layer_3_2[1167:1160]} - {1'b0, layer_2_2[1167:1160]};
      btm_2[1] = {1'b0,layer_3_2[1175:1168]} - {1'b0, layer_2_2[1175:1168]};
      btm_2[2] = {1'b0,layer_3_2[1183:1176]} - {1'b0, layer_2_2[1183:1176]};
    end
    'd147: begin
      top_0[0] = {1'b0,layer_1_0[1175:1168]} - {1'b0, layer_0_0[1175:1168]};
      top_0[1] = {1'b0,layer_1_0[1183:1176]} - {1'b0, layer_0_0[1183:1176]};
      top_0[2] = {1'b0,layer_1_0[1191:1184]} - {1'b0, layer_0_0[1191:1184]};
      top_1[0] = {1'b0,layer_1_1[1175:1168]} - {1'b0, layer_0_1[1175:1168]};
      top_1[1] = {1'b0,layer_1_1[1183:1176]} - {1'b0, layer_0_1[1183:1176]};
      top_1[2] = {1'b0,layer_1_1[1191:1184]} - {1'b0, layer_0_1[1191:1184]};
      top_2[0] = {1'b0,layer_1_2[1175:1168]} - {1'b0, layer_0_2[1175:1168]};
      top_2[1] = {1'b0,layer_1_2[1183:1176]} - {1'b0, layer_0_2[1183:1176]};
      top_2[2] = {1'b0,layer_1_2[1191:1184]} - {1'b0, layer_0_2[1191:1184]};
      mid_0[0] = {1'b0,layer_2_0[1175:1168]} - {1'b0, layer_1_0[1175:1168]};
      mid_0[1] = {1'b0,layer_2_0[1183:1176]} - {1'b0, layer_1_0[1183:1176]};
      mid_0[2] = {1'b0,layer_2_0[1191:1184]} - {1'b0, layer_1_0[1191:1184]};
      mid_1[0] = {1'b0,layer_2_1[1175:1168]} - {1'b0, layer_1_1[1175:1168]};
      mid_1[1] = {1'b0,layer_2_1[1183:1176]} - {1'b0, layer_1_1[1183:1176]};
      mid_1[2] = {1'b0,layer_2_1[1191:1184]} - {1'b0, layer_1_1[1191:1184]};
      mid_2[0] = {1'b0,layer_2_2[1175:1168]} - {1'b0, layer_1_2[1175:1168]};
      mid_2[1] = {1'b0,layer_2_2[1183:1176]} - {1'b0, layer_1_2[1183:1176]};
      mid_2[2] = {1'b0,layer_2_2[1191:1184]} - {1'b0, layer_1_2[1191:1184]};
      btm_0[0] = {1'b0,layer_3_0[1175:1168]} - {1'b0, layer_2_0[1175:1168]};
      btm_0[1] = {1'b0,layer_3_0[1183:1176]} - {1'b0, layer_2_0[1183:1176]};
      btm_0[2] = {1'b0,layer_3_0[1191:1184]} - {1'b0, layer_2_0[1191:1184]};
      btm_1[0] = {1'b0,layer_3_1[1175:1168]} - {1'b0, layer_2_1[1175:1168]};
      btm_1[1] = {1'b0,layer_3_1[1183:1176]} - {1'b0, layer_2_1[1183:1176]};
      btm_1[2] = {1'b0,layer_3_1[1191:1184]} - {1'b0, layer_2_1[1191:1184]};
      btm_2[0] = {1'b0,layer_3_2[1175:1168]} - {1'b0, layer_2_2[1175:1168]};
      btm_2[1] = {1'b0,layer_3_2[1183:1176]} - {1'b0, layer_2_2[1183:1176]};
      btm_2[2] = {1'b0,layer_3_2[1191:1184]} - {1'b0, layer_2_2[1191:1184]};
    end
    'd148: begin
      top_0[0] = {1'b0,layer_1_0[1183:1176]} - {1'b0, layer_0_0[1183:1176]};
      top_0[1] = {1'b0,layer_1_0[1191:1184]} - {1'b0, layer_0_0[1191:1184]};
      top_0[2] = {1'b0,layer_1_0[1199:1192]} - {1'b0, layer_0_0[1199:1192]};
      top_1[0] = {1'b0,layer_1_1[1183:1176]} - {1'b0, layer_0_1[1183:1176]};
      top_1[1] = {1'b0,layer_1_1[1191:1184]} - {1'b0, layer_0_1[1191:1184]};
      top_1[2] = {1'b0,layer_1_1[1199:1192]} - {1'b0, layer_0_1[1199:1192]};
      top_2[0] = {1'b0,layer_1_2[1183:1176]} - {1'b0, layer_0_2[1183:1176]};
      top_2[1] = {1'b0,layer_1_2[1191:1184]} - {1'b0, layer_0_2[1191:1184]};
      top_2[2] = {1'b0,layer_1_2[1199:1192]} - {1'b0, layer_0_2[1199:1192]};
      mid_0[0] = {1'b0,layer_2_0[1183:1176]} - {1'b0, layer_1_0[1183:1176]};
      mid_0[1] = {1'b0,layer_2_0[1191:1184]} - {1'b0, layer_1_0[1191:1184]};
      mid_0[2] = {1'b0,layer_2_0[1199:1192]} - {1'b0, layer_1_0[1199:1192]};
      mid_1[0] = {1'b0,layer_2_1[1183:1176]} - {1'b0, layer_1_1[1183:1176]};
      mid_1[1] = {1'b0,layer_2_1[1191:1184]} - {1'b0, layer_1_1[1191:1184]};
      mid_1[2] = {1'b0,layer_2_1[1199:1192]} - {1'b0, layer_1_1[1199:1192]};
      mid_2[0] = {1'b0,layer_2_2[1183:1176]} - {1'b0, layer_1_2[1183:1176]};
      mid_2[1] = {1'b0,layer_2_2[1191:1184]} - {1'b0, layer_1_2[1191:1184]};
      mid_2[2] = {1'b0,layer_2_2[1199:1192]} - {1'b0, layer_1_2[1199:1192]};
      btm_0[0] = {1'b0,layer_3_0[1183:1176]} - {1'b0, layer_2_0[1183:1176]};
      btm_0[1] = {1'b0,layer_3_0[1191:1184]} - {1'b0, layer_2_0[1191:1184]};
      btm_0[2] = {1'b0,layer_3_0[1199:1192]} - {1'b0, layer_2_0[1199:1192]};
      btm_1[0] = {1'b0,layer_3_1[1183:1176]} - {1'b0, layer_2_1[1183:1176]};
      btm_1[1] = {1'b0,layer_3_1[1191:1184]} - {1'b0, layer_2_1[1191:1184]};
      btm_1[2] = {1'b0,layer_3_1[1199:1192]} - {1'b0, layer_2_1[1199:1192]};
      btm_2[0] = {1'b0,layer_3_2[1183:1176]} - {1'b0, layer_2_2[1183:1176]};
      btm_2[1] = {1'b0,layer_3_2[1191:1184]} - {1'b0, layer_2_2[1191:1184]};
      btm_2[2] = {1'b0,layer_3_2[1199:1192]} - {1'b0, layer_2_2[1199:1192]};
    end
    'd149: begin
      top_0[0] = {1'b0,layer_1_0[1191:1184]} - {1'b0, layer_0_0[1191:1184]};
      top_0[1] = {1'b0,layer_1_0[1199:1192]} - {1'b0, layer_0_0[1199:1192]};
      top_0[2] = {1'b0,layer_1_0[1207:1200]} - {1'b0, layer_0_0[1207:1200]};
      top_1[0] = {1'b0,layer_1_1[1191:1184]} - {1'b0, layer_0_1[1191:1184]};
      top_1[1] = {1'b0,layer_1_1[1199:1192]} - {1'b0, layer_0_1[1199:1192]};
      top_1[2] = {1'b0,layer_1_1[1207:1200]} - {1'b0, layer_0_1[1207:1200]};
      top_2[0] = {1'b0,layer_1_2[1191:1184]} - {1'b0, layer_0_2[1191:1184]};
      top_2[1] = {1'b0,layer_1_2[1199:1192]} - {1'b0, layer_0_2[1199:1192]};
      top_2[2] = {1'b0,layer_1_2[1207:1200]} - {1'b0, layer_0_2[1207:1200]};
      mid_0[0] = {1'b0,layer_2_0[1191:1184]} - {1'b0, layer_1_0[1191:1184]};
      mid_0[1] = {1'b0,layer_2_0[1199:1192]} - {1'b0, layer_1_0[1199:1192]};
      mid_0[2] = {1'b0,layer_2_0[1207:1200]} - {1'b0, layer_1_0[1207:1200]};
      mid_1[0] = {1'b0,layer_2_1[1191:1184]} - {1'b0, layer_1_1[1191:1184]};
      mid_1[1] = {1'b0,layer_2_1[1199:1192]} - {1'b0, layer_1_1[1199:1192]};
      mid_1[2] = {1'b0,layer_2_1[1207:1200]} - {1'b0, layer_1_1[1207:1200]};
      mid_2[0] = {1'b0,layer_2_2[1191:1184]} - {1'b0, layer_1_2[1191:1184]};
      mid_2[1] = {1'b0,layer_2_2[1199:1192]} - {1'b0, layer_1_2[1199:1192]};
      mid_2[2] = {1'b0,layer_2_2[1207:1200]} - {1'b0, layer_1_2[1207:1200]};
      btm_0[0] = {1'b0,layer_3_0[1191:1184]} - {1'b0, layer_2_0[1191:1184]};
      btm_0[1] = {1'b0,layer_3_0[1199:1192]} - {1'b0, layer_2_0[1199:1192]};
      btm_0[2] = {1'b0,layer_3_0[1207:1200]} - {1'b0, layer_2_0[1207:1200]};
      btm_1[0] = {1'b0,layer_3_1[1191:1184]} - {1'b0, layer_2_1[1191:1184]};
      btm_1[1] = {1'b0,layer_3_1[1199:1192]} - {1'b0, layer_2_1[1199:1192]};
      btm_1[2] = {1'b0,layer_3_1[1207:1200]} - {1'b0, layer_2_1[1207:1200]};
      btm_2[0] = {1'b0,layer_3_2[1191:1184]} - {1'b0, layer_2_2[1191:1184]};
      btm_2[1] = {1'b0,layer_3_2[1199:1192]} - {1'b0, layer_2_2[1199:1192]};
      btm_2[2] = {1'b0,layer_3_2[1207:1200]} - {1'b0, layer_2_2[1207:1200]};
    end
    'd150: begin
      top_0[0] = {1'b0,layer_1_0[1199:1192]} - {1'b0, layer_0_0[1199:1192]};
      top_0[1] = {1'b0,layer_1_0[1207:1200]} - {1'b0, layer_0_0[1207:1200]};
      top_0[2] = {1'b0,layer_1_0[1215:1208]} - {1'b0, layer_0_0[1215:1208]};
      top_1[0] = {1'b0,layer_1_1[1199:1192]} - {1'b0, layer_0_1[1199:1192]};
      top_1[1] = {1'b0,layer_1_1[1207:1200]} - {1'b0, layer_0_1[1207:1200]};
      top_1[2] = {1'b0,layer_1_1[1215:1208]} - {1'b0, layer_0_1[1215:1208]};
      top_2[0] = {1'b0,layer_1_2[1199:1192]} - {1'b0, layer_0_2[1199:1192]};
      top_2[1] = {1'b0,layer_1_2[1207:1200]} - {1'b0, layer_0_2[1207:1200]};
      top_2[2] = {1'b0,layer_1_2[1215:1208]} - {1'b0, layer_0_2[1215:1208]};
      mid_0[0] = {1'b0,layer_2_0[1199:1192]} - {1'b0, layer_1_0[1199:1192]};
      mid_0[1] = {1'b0,layer_2_0[1207:1200]} - {1'b0, layer_1_0[1207:1200]};
      mid_0[2] = {1'b0,layer_2_0[1215:1208]} - {1'b0, layer_1_0[1215:1208]};
      mid_1[0] = {1'b0,layer_2_1[1199:1192]} - {1'b0, layer_1_1[1199:1192]};
      mid_1[1] = {1'b0,layer_2_1[1207:1200]} - {1'b0, layer_1_1[1207:1200]};
      mid_1[2] = {1'b0,layer_2_1[1215:1208]} - {1'b0, layer_1_1[1215:1208]};
      mid_2[0] = {1'b0,layer_2_2[1199:1192]} - {1'b0, layer_1_2[1199:1192]};
      mid_2[1] = {1'b0,layer_2_2[1207:1200]} - {1'b0, layer_1_2[1207:1200]};
      mid_2[2] = {1'b0,layer_2_2[1215:1208]} - {1'b0, layer_1_2[1215:1208]};
      btm_0[0] = {1'b0,layer_3_0[1199:1192]} - {1'b0, layer_2_0[1199:1192]};
      btm_0[1] = {1'b0,layer_3_0[1207:1200]} - {1'b0, layer_2_0[1207:1200]};
      btm_0[2] = {1'b0,layer_3_0[1215:1208]} - {1'b0, layer_2_0[1215:1208]};
      btm_1[0] = {1'b0,layer_3_1[1199:1192]} - {1'b0, layer_2_1[1199:1192]};
      btm_1[1] = {1'b0,layer_3_1[1207:1200]} - {1'b0, layer_2_1[1207:1200]};
      btm_1[2] = {1'b0,layer_3_1[1215:1208]} - {1'b0, layer_2_1[1215:1208]};
      btm_2[0] = {1'b0,layer_3_2[1199:1192]} - {1'b0, layer_2_2[1199:1192]};
      btm_2[1] = {1'b0,layer_3_2[1207:1200]} - {1'b0, layer_2_2[1207:1200]};
      btm_2[2] = {1'b0,layer_3_2[1215:1208]} - {1'b0, layer_2_2[1215:1208]};
    end
    'd151: begin
      top_0[0] = {1'b0,layer_1_0[1207:1200]} - {1'b0, layer_0_0[1207:1200]};
      top_0[1] = {1'b0,layer_1_0[1215:1208]} - {1'b0, layer_0_0[1215:1208]};
      top_0[2] = {1'b0,layer_1_0[1223:1216]} - {1'b0, layer_0_0[1223:1216]};
      top_1[0] = {1'b0,layer_1_1[1207:1200]} - {1'b0, layer_0_1[1207:1200]};
      top_1[1] = {1'b0,layer_1_1[1215:1208]} - {1'b0, layer_0_1[1215:1208]};
      top_1[2] = {1'b0,layer_1_1[1223:1216]} - {1'b0, layer_0_1[1223:1216]};
      top_2[0] = {1'b0,layer_1_2[1207:1200]} - {1'b0, layer_0_2[1207:1200]};
      top_2[1] = {1'b0,layer_1_2[1215:1208]} - {1'b0, layer_0_2[1215:1208]};
      top_2[2] = {1'b0,layer_1_2[1223:1216]} - {1'b0, layer_0_2[1223:1216]};
      mid_0[0] = {1'b0,layer_2_0[1207:1200]} - {1'b0, layer_1_0[1207:1200]};
      mid_0[1] = {1'b0,layer_2_0[1215:1208]} - {1'b0, layer_1_0[1215:1208]};
      mid_0[2] = {1'b0,layer_2_0[1223:1216]} - {1'b0, layer_1_0[1223:1216]};
      mid_1[0] = {1'b0,layer_2_1[1207:1200]} - {1'b0, layer_1_1[1207:1200]};
      mid_1[1] = {1'b0,layer_2_1[1215:1208]} - {1'b0, layer_1_1[1215:1208]};
      mid_1[2] = {1'b0,layer_2_1[1223:1216]} - {1'b0, layer_1_1[1223:1216]};
      mid_2[0] = {1'b0,layer_2_2[1207:1200]} - {1'b0, layer_1_2[1207:1200]};
      mid_2[1] = {1'b0,layer_2_2[1215:1208]} - {1'b0, layer_1_2[1215:1208]};
      mid_2[2] = {1'b0,layer_2_2[1223:1216]} - {1'b0, layer_1_2[1223:1216]};
      btm_0[0] = {1'b0,layer_3_0[1207:1200]} - {1'b0, layer_2_0[1207:1200]};
      btm_0[1] = {1'b0,layer_3_0[1215:1208]} - {1'b0, layer_2_0[1215:1208]};
      btm_0[2] = {1'b0,layer_3_0[1223:1216]} - {1'b0, layer_2_0[1223:1216]};
      btm_1[0] = {1'b0,layer_3_1[1207:1200]} - {1'b0, layer_2_1[1207:1200]};
      btm_1[1] = {1'b0,layer_3_1[1215:1208]} - {1'b0, layer_2_1[1215:1208]};
      btm_1[2] = {1'b0,layer_3_1[1223:1216]} - {1'b0, layer_2_1[1223:1216]};
      btm_2[0] = {1'b0,layer_3_2[1207:1200]} - {1'b0, layer_2_2[1207:1200]};
      btm_2[1] = {1'b0,layer_3_2[1215:1208]} - {1'b0, layer_2_2[1215:1208]};
      btm_2[2] = {1'b0,layer_3_2[1223:1216]} - {1'b0, layer_2_2[1223:1216]};
    end
    'd152: begin
      top_0[0] = {1'b0,layer_1_0[1215:1208]} - {1'b0, layer_0_0[1215:1208]};
      top_0[1] = {1'b0,layer_1_0[1223:1216]} - {1'b0, layer_0_0[1223:1216]};
      top_0[2] = {1'b0,layer_1_0[1231:1224]} - {1'b0, layer_0_0[1231:1224]};
      top_1[0] = {1'b0,layer_1_1[1215:1208]} - {1'b0, layer_0_1[1215:1208]};
      top_1[1] = {1'b0,layer_1_1[1223:1216]} - {1'b0, layer_0_1[1223:1216]};
      top_1[2] = {1'b0,layer_1_1[1231:1224]} - {1'b0, layer_0_1[1231:1224]};
      top_2[0] = {1'b0,layer_1_2[1215:1208]} - {1'b0, layer_0_2[1215:1208]};
      top_2[1] = {1'b0,layer_1_2[1223:1216]} - {1'b0, layer_0_2[1223:1216]};
      top_2[2] = {1'b0,layer_1_2[1231:1224]} - {1'b0, layer_0_2[1231:1224]};
      mid_0[0] = {1'b0,layer_2_0[1215:1208]} - {1'b0, layer_1_0[1215:1208]};
      mid_0[1] = {1'b0,layer_2_0[1223:1216]} - {1'b0, layer_1_0[1223:1216]};
      mid_0[2] = {1'b0,layer_2_0[1231:1224]} - {1'b0, layer_1_0[1231:1224]};
      mid_1[0] = {1'b0,layer_2_1[1215:1208]} - {1'b0, layer_1_1[1215:1208]};
      mid_1[1] = {1'b0,layer_2_1[1223:1216]} - {1'b0, layer_1_1[1223:1216]};
      mid_1[2] = {1'b0,layer_2_1[1231:1224]} - {1'b0, layer_1_1[1231:1224]};
      mid_2[0] = {1'b0,layer_2_2[1215:1208]} - {1'b0, layer_1_2[1215:1208]};
      mid_2[1] = {1'b0,layer_2_2[1223:1216]} - {1'b0, layer_1_2[1223:1216]};
      mid_2[2] = {1'b0,layer_2_2[1231:1224]} - {1'b0, layer_1_2[1231:1224]};
      btm_0[0] = {1'b0,layer_3_0[1215:1208]} - {1'b0, layer_2_0[1215:1208]};
      btm_0[1] = {1'b0,layer_3_0[1223:1216]} - {1'b0, layer_2_0[1223:1216]};
      btm_0[2] = {1'b0,layer_3_0[1231:1224]} - {1'b0, layer_2_0[1231:1224]};
      btm_1[0] = {1'b0,layer_3_1[1215:1208]} - {1'b0, layer_2_1[1215:1208]};
      btm_1[1] = {1'b0,layer_3_1[1223:1216]} - {1'b0, layer_2_1[1223:1216]};
      btm_1[2] = {1'b0,layer_3_1[1231:1224]} - {1'b0, layer_2_1[1231:1224]};
      btm_2[0] = {1'b0,layer_3_2[1215:1208]} - {1'b0, layer_2_2[1215:1208]};
      btm_2[1] = {1'b0,layer_3_2[1223:1216]} - {1'b0, layer_2_2[1223:1216]};
      btm_2[2] = {1'b0,layer_3_2[1231:1224]} - {1'b0, layer_2_2[1231:1224]};
    end
    'd153: begin
      top_0[0] = {1'b0,layer_1_0[1223:1216]} - {1'b0, layer_0_0[1223:1216]};
      top_0[1] = {1'b0,layer_1_0[1231:1224]} - {1'b0, layer_0_0[1231:1224]};
      top_0[2] = {1'b0,layer_1_0[1239:1232]} - {1'b0, layer_0_0[1239:1232]};
      top_1[0] = {1'b0,layer_1_1[1223:1216]} - {1'b0, layer_0_1[1223:1216]};
      top_1[1] = {1'b0,layer_1_1[1231:1224]} - {1'b0, layer_0_1[1231:1224]};
      top_1[2] = {1'b0,layer_1_1[1239:1232]} - {1'b0, layer_0_1[1239:1232]};
      top_2[0] = {1'b0,layer_1_2[1223:1216]} - {1'b0, layer_0_2[1223:1216]};
      top_2[1] = {1'b0,layer_1_2[1231:1224]} - {1'b0, layer_0_2[1231:1224]};
      top_2[2] = {1'b0,layer_1_2[1239:1232]} - {1'b0, layer_0_2[1239:1232]};
      mid_0[0] = {1'b0,layer_2_0[1223:1216]} - {1'b0, layer_1_0[1223:1216]};
      mid_0[1] = {1'b0,layer_2_0[1231:1224]} - {1'b0, layer_1_0[1231:1224]};
      mid_0[2] = {1'b0,layer_2_0[1239:1232]} - {1'b0, layer_1_0[1239:1232]};
      mid_1[0] = {1'b0,layer_2_1[1223:1216]} - {1'b0, layer_1_1[1223:1216]};
      mid_1[1] = {1'b0,layer_2_1[1231:1224]} - {1'b0, layer_1_1[1231:1224]};
      mid_1[2] = {1'b0,layer_2_1[1239:1232]} - {1'b0, layer_1_1[1239:1232]};
      mid_2[0] = {1'b0,layer_2_2[1223:1216]} - {1'b0, layer_1_2[1223:1216]};
      mid_2[1] = {1'b0,layer_2_2[1231:1224]} - {1'b0, layer_1_2[1231:1224]};
      mid_2[2] = {1'b0,layer_2_2[1239:1232]} - {1'b0, layer_1_2[1239:1232]};
      btm_0[0] = {1'b0,layer_3_0[1223:1216]} - {1'b0, layer_2_0[1223:1216]};
      btm_0[1] = {1'b0,layer_3_0[1231:1224]} - {1'b0, layer_2_0[1231:1224]};
      btm_0[2] = {1'b0,layer_3_0[1239:1232]} - {1'b0, layer_2_0[1239:1232]};
      btm_1[0] = {1'b0,layer_3_1[1223:1216]} - {1'b0, layer_2_1[1223:1216]};
      btm_1[1] = {1'b0,layer_3_1[1231:1224]} - {1'b0, layer_2_1[1231:1224]};
      btm_1[2] = {1'b0,layer_3_1[1239:1232]} - {1'b0, layer_2_1[1239:1232]};
      btm_2[0] = {1'b0,layer_3_2[1223:1216]} - {1'b0, layer_2_2[1223:1216]};
      btm_2[1] = {1'b0,layer_3_2[1231:1224]} - {1'b0, layer_2_2[1231:1224]};
      btm_2[2] = {1'b0,layer_3_2[1239:1232]} - {1'b0, layer_2_2[1239:1232]};
    end
    'd154: begin
      top_0[0] = {1'b0,layer_1_0[1231:1224]} - {1'b0, layer_0_0[1231:1224]};
      top_0[1] = {1'b0,layer_1_0[1239:1232]} - {1'b0, layer_0_0[1239:1232]};
      top_0[2] = {1'b0,layer_1_0[1247:1240]} - {1'b0, layer_0_0[1247:1240]};
      top_1[0] = {1'b0,layer_1_1[1231:1224]} - {1'b0, layer_0_1[1231:1224]};
      top_1[1] = {1'b0,layer_1_1[1239:1232]} - {1'b0, layer_0_1[1239:1232]};
      top_1[2] = {1'b0,layer_1_1[1247:1240]} - {1'b0, layer_0_1[1247:1240]};
      top_2[0] = {1'b0,layer_1_2[1231:1224]} - {1'b0, layer_0_2[1231:1224]};
      top_2[1] = {1'b0,layer_1_2[1239:1232]} - {1'b0, layer_0_2[1239:1232]};
      top_2[2] = {1'b0,layer_1_2[1247:1240]} - {1'b0, layer_0_2[1247:1240]};
      mid_0[0] = {1'b0,layer_2_0[1231:1224]} - {1'b0, layer_1_0[1231:1224]};
      mid_0[1] = {1'b0,layer_2_0[1239:1232]} - {1'b0, layer_1_0[1239:1232]};
      mid_0[2] = {1'b0,layer_2_0[1247:1240]} - {1'b0, layer_1_0[1247:1240]};
      mid_1[0] = {1'b0,layer_2_1[1231:1224]} - {1'b0, layer_1_1[1231:1224]};
      mid_1[1] = {1'b0,layer_2_1[1239:1232]} - {1'b0, layer_1_1[1239:1232]};
      mid_1[2] = {1'b0,layer_2_1[1247:1240]} - {1'b0, layer_1_1[1247:1240]};
      mid_2[0] = {1'b0,layer_2_2[1231:1224]} - {1'b0, layer_1_2[1231:1224]};
      mid_2[1] = {1'b0,layer_2_2[1239:1232]} - {1'b0, layer_1_2[1239:1232]};
      mid_2[2] = {1'b0,layer_2_2[1247:1240]} - {1'b0, layer_1_2[1247:1240]};
      btm_0[0] = {1'b0,layer_3_0[1231:1224]} - {1'b0, layer_2_0[1231:1224]};
      btm_0[1] = {1'b0,layer_3_0[1239:1232]} - {1'b0, layer_2_0[1239:1232]};
      btm_0[2] = {1'b0,layer_3_0[1247:1240]} - {1'b0, layer_2_0[1247:1240]};
      btm_1[0] = {1'b0,layer_3_1[1231:1224]} - {1'b0, layer_2_1[1231:1224]};
      btm_1[1] = {1'b0,layer_3_1[1239:1232]} - {1'b0, layer_2_1[1239:1232]};
      btm_1[2] = {1'b0,layer_3_1[1247:1240]} - {1'b0, layer_2_1[1247:1240]};
      btm_2[0] = {1'b0,layer_3_2[1231:1224]} - {1'b0, layer_2_2[1231:1224]};
      btm_2[1] = {1'b0,layer_3_2[1239:1232]} - {1'b0, layer_2_2[1239:1232]};
      btm_2[2] = {1'b0,layer_3_2[1247:1240]} - {1'b0, layer_2_2[1247:1240]};
    end
    'd155: begin
      top_0[0] = {1'b0,layer_1_0[1239:1232]} - {1'b0, layer_0_0[1239:1232]};
      top_0[1] = {1'b0,layer_1_0[1247:1240]} - {1'b0, layer_0_0[1247:1240]};
      top_0[2] = {1'b0,layer_1_0[1255:1248]} - {1'b0, layer_0_0[1255:1248]};
      top_1[0] = {1'b0,layer_1_1[1239:1232]} - {1'b0, layer_0_1[1239:1232]};
      top_1[1] = {1'b0,layer_1_1[1247:1240]} - {1'b0, layer_0_1[1247:1240]};
      top_1[2] = {1'b0,layer_1_1[1255:1248]} - {1'b0, layer_0_1[1255:1248]};
      top_2[0] = {1'b0,layer_1_2[1239:1232]} - {1'b0, layer_0_2[1239:1232]};
      top_2[1] = {1'b0,layer_1_2[1247:1240]} - {1'b0, layer_0_2[1247:1240]};
      top_2[2] = {1'b0,layer_1_2[1255:1248]} - {1'b0, layer_0_2[1255:1248]};
      mid_0[0] = {1'b0,layer_2_0[1239:1232]} - {1'b0, layer_1_0[1239:1232]};
      mid_0[1] = {1'b0,layer_2_0[1247:1240]} - {1'b0, layer_1_0[1247:1240]};
      mid_0[2] = {1'b0,layer_2_0[1255:1248]} - {1'b0, layer_1_0[1255:1248]};
      mid_1[0] = {1'b0,layer_2_1[1239:1232]} - {1'b0, layer_1_1[1239:1232]};
      mid_1[1] = {1'b0,layer_2_1[1247:1240]} - {1'b0, layer_1_1[1247:1240]};
      mid_1[2] = {1'b0,layer_2_1[1255:1248]} - {1'b0, layer_1_1[1255:1248]};
      mid_2[0] = {1'b0,layer_2_2[1239:1232]} - {1'b0, layer_1_2[1239:1232]};
      mid_2[1] = {1'b0,layer_2_2[1247:1240]} - {1'b0, layer_1_2[1247:1240]};
      mid_2[2] = {1'b0,layer_2_2[1255:1248]} - {1'b0, layer_1_2[1255:1248]};
      btm_0[0] = {1'b0,layer_3_0[1239:1232]} - {1'b0, layer_2_0[1239:1232]};
      btm_0[1] = {1'b0,layer_3_0[1247:1240]} - {1'b0, layer_2_0[1247:1240]};
      btm_0[2] = {1'b0,layer_3_0[1255:1248]} - {1'b0, layer_2_0[1255:1248]};
      btm_1[0] = {1'b0,layer_3_1[1239:1232]} - {1'b0, layer_2_1[1239:1232]};
      btm_1[1] = {1'b0,layer_3_1[1247:1240]} - {1'b0, layer_2_1[1247:1240]};
      btm_1[2] = {1'b0,layer_3_1[1255:1248]} - {1'b0, layer_2_1[1255:1248]};
      btm_2[0] = {1'b0,layer_3_2[1239:1232]} - {1'b0, layer_2_2[1239:1232]};
      btm_2[1] = {1'b0,layer_3_2[1247:1240]} - {1'b0, layer_2_2[1247:1240]};
      btm_2[2] = {1'b0,layer_3_2[1255:1248]} - {1'b0, layer_2_2[1255:1248]};
    end
    'd156: begin
      top_0[0] = {1'b0,layer_1_0[1247:1240]} - {1'b0, layer_0_0[1247:1240]};
      top_0[1] = {1'b0,layer_1_0[1255:1248]} - {1'b0, layer_0_0[1255:1248]};
      top_0[2] = {1'b0,layer_1_0[1263:1256]} - {1'b0, layer_0_0[1263:1256]};
      top_1[0] = {1'b0,layer_1_1[1247:1240]} - {1'b0, layer_0_1[1247:1240]};
      top_1[1] = {1'b0,layer_1_1[1255:1248]} - {1'b0, layer_0_1[1255:1248]};
      top_1[2] = {1'b0,layer_1_1[1263:1256]} - {1'b0, layer_0_1[1263:1256]};
      top_2[0] = {1'b0,layer_1_2[1247:1240]} - {1'b0, layer_0_2[1247:1240]};
      top_2[1] = {1'b0,layer_1_2[1255:1248]} - {1'b0, layer_0_2[1255:1248]};
      top_2[2] = {1'b0,layer_1_2[1263:1256]} - {1'b0, layer_0_2[1263:1256]};
      mid_0[0] = {1'b0,layer_2_0[1247:1240]} - {1'b0, layer_1_0[1247:1240]};
      mid_0[1] = {1'b0,layer_2_0[1255:1248]} - {1'b0, layer_1_0[1255:1248]};
      mid_0[2] = {1'b0,layer_2_0[1263:1256]} - {1'b0, layer_1_0[1263:1256]};
      mid_1[0] = {1'b0,layer_2_1[1247:1240]} - {1'b0, layer_1_1[1247:1240]};
      mid_1[1] = {1'b0,layer_2_1[1255:1248]} - {1'b0, layer_1_1[1255:1248]};
      mid_1[2] = {1'b0,layer_2_1[1263:1256]} - {1'b0, layer_1_1[1263:1256]};
      mid_2[0] = {1'b0,layer_2_2[1247:1240]} - {1'b0, layer_1_2[1247:1240]};
      mid_2[1] = {1'b0,layer_2_2[1255:1248]} - {1'b0, layer_1_2[1255:1248]};
      mid_2[2] = {1'b0,layer_2_2[1263:1256]} - {1'b0, layer_1_2[1263:1256]};
      btm_0[0] = {1'b0,layer_3_0[1247:1240]} - {1'b0, layer_2_0[1247:1240]};
      btm_0[1] = {1'b0,layer_3_0[1255:1248]} - {1'b0, layer_2_0[1255:1248]};
      btm_0[2] = {1'b0,layer_3_0[1263:1256]} - {1'b0, layer_2_0[1263:1256]};
      btm_1[0] = {1'b0,layer_3_1[1247:1240]} - {1'b0, layer_2_1[1247:1240]};
      btm_1[1] = {1'b0,layer_3_1[1255:1248]} - {1'b0, layer_2_1[1255:1248]};
      btm_1[2] = {1'b0,layer_3_1[1263:1256]} - {1'b0, layer_2_1[1263:1256]};
      btm_2[0] = {1'b0,layer_3_2[1247:1240]} - {1'b0, layer_2_2[1247:1240]};
      btm_2[1] = {1'b0,layer_3_2[1255:1248]} - {1'b0, layer_2_2[1255:1248]};
      btm_2[2] = {1'b0,layer_3_2[1263:1256]} - {1'b0, layer_2_2[1263:1256]};
    end
    'd157: begin
      top_0[0] = {1'b0,layer_1_0[1255:1248]} - {1'b0, layer_0_0[1255:1248]};
      top_0[1] = {1'b0,layer_1_0[1263:1256]} - {1'b0, layer_0_0[1263:1256]};
      top_0[2] = {1'b0,layer_1_0[1271:1264]} - {1'b0, layer_0_0[1271:1264]};
      top_1[0] = {1'b0,layer_1_1[1255:1248]} - {1'b0, layer_0_1[1255:1248]};
      top_1[1] = {1'b0,layer_1_1[1263:1256]} - {1'b0, layer_0_1[1263:1256]};
      top_1[2] = {1'b0,layer_1_1[1271:1264]} - {1'b0, layer_0_1[1271:1264]};
      top_2[0] = {1'b0,layer_1_2[1255:1248]} - {1'b0, layer_0_2[1255:1248]};
      top_2[1] = {1'b0,layer_1_2[1263:1256]} - {1'b0, layer_0_2[1263:1256]};
      top_2[2] = {1'b0,layer_1_2[1271:1264]} - {1'b0, layer_0_2[1271:1264]};
      mid_0[0] = {1'b0,layer_2_0[1255:1248]} - {1'b0, layer_1_0[1255:1248]};
      mid_0[1] = {1'b0,layer_2_0[1263:1256]} - {1'b0, layer_1_0[1263:1256]};
      mid_0[2] = {1'b0,layer_2_0[1271:1264]} - {1'b0, layer_1_0[1271:1264]};
      mid_1[0] = {1'b0,layer_2_1[1255:1248]} - {1'b0, layer_1_1[1255:1248]};
      mid_1[1] = {1'b0,layer_2_1[1263:1256]} - {1'b0, layer_1_1[1263:1256]};
      mid_1[2] = {1'b0,layer_2_1[1271:1264]} - {1'b0, layer_1_1[1271:1264]};
      mid_2[0] = {1'b0,layer_2_2[1255:1248]} - {1'b0, layer_1_2[1255:1248]};
      mid_2[1] = {1'b0,layer_2_2[1263:1256]} - {1'b0, layer_1_2[1263:1256]};
      mid_2[2] = {1'b0,layer_2_2[1271:1264]} - {1'b0, layer_1_2[1271:1264]};
      btm_0[0] = {1'b0,layer_3_0[1255:1248]} - {1'b0, layer_2_0[1255:1248]};
      btm_0[1] = {1'b0,layer_3_0[1263:1256]} - {1'b0, layer_2_0[1263:1256]};
      btm_0[2] = {1'b0,layer_3_0[1271:1264]} - {1'b0, layer_2_0[1271:1264]};
      btm_1[0] = {1'b0,layer_3_1[1255:1248]} - {1'b0, layer_2_1[1255:1248]};
      btm_1[1] = {1'b0,layer_3_1[1263:1256]} - {1'b0, layer_2_1[1263:1256]};
      btm_1[2] = {1'b0,layer_3_1[1271:1264]} - {1'b0, layer_2_1[1271:1264]};
      btm_2[0] = {1'b0,layer_3_2[1255:1248]} - {1'b0, layer_2_2[1255:1248]};
      btm_2[1] = {1'b0,layer_3_2[1263:1256]} - {1'b0, layer_2_2[1263:1256]};
      btm_2[2] = {1'b0,layer_3_2[1271:1264]} - {1'b0, layer_2_2[1271:1264]};
    end
    'd158: begin
      top_0[0] = {1'b0,layer_1_0[1263:1256]} - {1'b0, layer_0_0[1263:1256]};
      top_0[1] = {1'b0,layer_1_0[1271:1264]} - {1'b0, layer_0_0[1271:1264]};
      top_0[2] = {1'b0,layer_1_0[1279:1272]} - {1'b0, layer_0_0[1279:1272]};
      top_1[0] = {1'b0,layer_1_1[1263:1256]} - {1'b0, layer_0_1[1263:1256]};
      top_1[1] = {1'b0,layer_1_1[1271:1264]} - {1'b0, layer_0_1[1271:1264]};
      top_1[2] = {1'b0,layer_1_1[1279:1272]} - {1'b0, layer_0_1[1279:1272]};
      top_2[0] = {1'b0,layer_1_2[1263:1256]} - {1'b0, layer_0_2[1263:1256]};
      top_2[1] = {1'b0,layer_1_2[1271:1264]} - {1'b0, layer_0_2[1271:1264]};
      top_2[2] = {1'b0,layer_1_2[1279:1272]} - {1'b0, layer_0_2[1279:1272]};
      mid_0[0] = {1'b0,layer_2_0[1263:1256]} - {1'b0, layer_1_0[1263:1256]};
      mid_0[1] = {1'b0,layer_2_0[1271:1264]} - {1'b0, layer_1_0[1271:1264]};
      mid_0[2] = {1'b0,layer_2_0[1279:1272]} - {1'b0, layer_1_0[1279:1272]};
      mid_1[0] = {1'b0,layer_2_1[1263:1256]} - {1'b0, layer_1_1[1263:1256]};
      mid_1[1] = {1'b0,layer_2_1[1271:1264]} - {1'b0, layer_1_1[1271:1264]};
      mid_1[2] = {1'b0,layer_2_1[1279:1272]} - {1'b0, layer_1_1[1279:1272]};
      mid_2[0] = {1'b0,layer_2_2[1263:1256]} - {1'b0, layer_1_2[1263:1256]};
      mid_2[1] = {1'b0,layer_2_2[1271:1264]} - {1'b0, layer_1_2[1271:1264]};
      mid_2[2] = {1'b0,layer_2_2[1279:1272]} - {1'b0, layer_1_2[1279:1272]};
      btm_0[0] = {1'b0,layer_3_0[1263:1256]} - {1'b0, layer_2_0[1263:1256]};
      btm_0[1] = {1'b0,layer_3_0[1271:1264]} - {1'b0, layer_2_0[1271:1264]};
      btm_0[2] = {1'b0,layer_3_0[1279:1272]} - {1'b0, layer_2_0[1279:1272]};
      btm_1[0] = {1'b0,layer_3_1[1263:1256]} - {1'b0, layer_2_1[1263:1256]};
      btm_1[1] = {1'b0,layer_3_1[1271:1264]} - {1'b0, layer_2_1[1271:1264]};
      btm_1[2] = {1'b0,layer_3_1[1279:1272]} - {1'b0, layer_2_1[1279:1272]};
      btm_2[0] = {1'b0,layer_3_2[1263:1256]} - {1'b0, layer_2_2[1263:1256]};
      btm_2[1] = {1'b0,layer_3_2[1271:1264]} - {1'b0, layer_2_2[1271:1264]};
      btm_2[2] = {1'b0,layer_3_2[1279:1272]} - {1'b0, layer_2_2[1279:1272]};
    end
    'd159: begin
      top_0[0] = {1'b0,layer_1_0[1271:1264]} - {1'b0, layer_0_0[1271:1264]};
      top_0[1] = {1'b0,layer_1_0[1279:1272]} - {1'b0, layer_0_0[1279:1272]};
      top_0[2] = {1'b0,layer_1_0[1287:1280]} - {1'b0, layer_0_0[1287:1280]};
      top_1[0] = {1'b0,layer_1_1[1271:1264]} - {1'b0, layer_0_1[1271:1264]};
      top_1[1] = {1'b0,layer_1_1[1279:1272]} - {1'b0, layer_0_1[1279:1272]};
      top_1[2] = {1'b0,layer_1_1[1287:1280]} - {1'b0, layer_0_1[1287:1280]};
      top_2[0] = {1'b0,layer_1_2[1271:1264]} - {1'b0, layer_0_2[1271:1264]};
      top_2[1] = {1'b0,layer_1_2[1279:1272]} - {1'b0, layer_0_2[1279:1272]};
      top_2[2] = {1'b0,layer_1_2[1287:1280]} - {1'b0, layer_0_2[1287:1280]};
      mid_0[0] = {1'b0,layer_2_0[1271:1264]} - {1'b0, layer_1_0[1271:1264]};
      mid_0[1] = {1'b0,layer_2_0[1279:1272]} - {1'b0, layer_1_0[1279:1272]};
      mid_0[2] = {1'b0,layer_2_0[1287:1280]} - {1'b0, layer_1_0[1287:1280]};
      mid_1[0] = {1'b0,layer_2_1[1271:1264]} - {1'b0, layer_1_1[1271:1264]};
      mid_1[1] = {1'b0,layer_2_1[1279:1272]} - {1'b0, layer_1_1[1279:1272]};
      mid_1[2] = {1'b0,layer_2_1[1287:1280]} - {1'b0, layer_1_1[1287:1280]};
      mid_2[0] = {1'b0,layer_2_2[1271:1264]} - {1'b0, layer_1_2[1271:1264]};
      mid_2[1] = {1'b0,layer_2_2[1279:1272]} - {1'b0, layer_1_2[1279:1272]};
      mid_2[2] = {1'b0,layer_2_2[1287:1280]} - {1'b0, layer_1_2[1287:1280]};
      btm_0[0] = {1'b0,layer_3_0[1271:1264]} - {1'b0, layer_2_0[1271:1264]};
      btm_0[1] = {1'b0,layer_3_0[1279:1272]} - {1'b0, layer_2_0[1279:1272]};
      btm_0[2] = {1'b0,layer_3_0[1287:1280]} - {1'b0, layer_2_0[1287:1280]};
      btm_1[0] = {1'b0,layer_3_1[1271:1264]} - {1'b0, layer_2_1[1271:1264]};
      btm_1[1] = {1'b0,layer_3_1[1279:1272]} - {1'b0, layer_2_1[1279:1272]};
      btm_1[2] = {1'b0,layer_3_1[1287:1280]} - {1'b0, layer_2_1[1287:1280]};
      btm_2[0] = {1'b0,layer_3_2[1271:1264]} - {1'b0, layer_2_2[1271:1264]};
      btm_2[1] = {1'b0,layer_3_2[1279:1272]} - {1'b0, layer_2_2[1279:1272]};
      btm_2[2] = {1'b0,layer_3_2[1287:1280]} - {1'b0, layer_2_2[1287:1280]};
    end
    'd160: begin
      top_0[0] = {1'b0,layer_1_0[1279:1272]} - {1'b0, layer_0_0[1279:1272]};
      top_0[1] = {1'b0,layer_1_0[1287:1280]} - {1'b0, layer_0_0[1287:1280]};
      top_0[2] = {1'b0,layer_1_0[1295:1288]} - {1'b0, layer_0_0[1295:1288]};
      top_1[0] = {1'b0,layer_1_1[1279:1272]} - {1'b0, layer_0_1[1279:1272]};
      top_1[1] = {1'b0,layer_1_1[1287:1280]} - {1'b0, layer_0_1[1287:1280]};
      top_1[2] = {1'b0,layer_1_1[1295:1288]} - {1'b0, layer_0_1[1295:1288]};
      top_2[0] = {1'b0,layer_1_2[1279:1272]} - {1'b0, layer_0_2[1279:1272]};
      top_2[1] = {1'b0,layer_1_2[1287:1280]} - {1'b0, layer_0_2[1287:1280]};
      top_2[2] = {1'b0,layer_1_2[1295:1288]} - {1'b0, layer_0_2[1295:1288]};
      mid_0[0] = {1'b0,layer_2_0[1279:1272]} - {1'b0, layer_1_0[1279:1272]};
      mid_0[1] = {1'b0,layer_2_0[1287:1280]} - {1'b0, layer_1_0[1287:1280]};
      mid_0[2] = {1'b0,layer_2_0[1295:1288]} - {1'b0, layer_1_0[1295:1288]};
      mid_1[0] = {1'b0,layer_2_1[1279:1272]} - {1'b0, layer_1_1[1279:1272]};
      mid_1[1] = {1'b0,layer_2_1[1287:1280]} - {1'b0, layer_1_1[1287:1280]};
      mid_1[2] = {1'b0,layer_2_1[1295:1288]} - {1'b0, layer_1_1[1295:1288]};
      mid_2[0] = {1'b0,layer_2_2[1279:1272]} - {1'b0, layer_1_2[1279:1272]};
      mid_2[1] = {1'b0,layer_2_2[1287:1280]} - {1'b0, layer_1_2[1287:1280]};
      mid_2[2] = {1'b0,layer_2_2[1295:1288]} - {1'b0, layer_1_2[1295:1288]};
      btm_0[0] = {1'b0,layer_3_0[1279:1272]} - {1'b0, layer_2_0[1279:1272]};
      btm_0[1] = {1'b0,layer_3_0[1287:1280]} - {1'b0, layer_2_0[1287:1280]};
      btm_0[2] = {1'b0,layer_3_0[1295:1288]} - {1'b0, layer_2_0[1295:1288]};
      btm_1[0] = {1'b0,layer_3_1[1279:1272]} - {1'b0, layer_2_1[1279:1272]};
      btm_1[1] = {1'b0,layer_3_1[1287:1280]} - {1'b0, layer_2_1[1287:1280]};
      btm_1[2] = {1'b0,layer_3_1[1295:1288]} - {1'b0, layer_2_1[1295:1288]};
      btm_2[0] = {1'b0,layer_3_2[1279:1272]} - {1'b0, layer_2_2[1279:1272]};
      btm_2[1] = {1'b0,layer_3_2[1287:1280]} - {1'b0, layer_2_2[1287:1280]};
      btm_2[2] = {1'b0,layer_3_2[1295:1288]} - {1'b0, layer_2_2[1295:1288]};
    end
    'd161: begin
      top_0[0] = {1'b0,layer_1_0[1287:1280]} - {1'b0, layer_0_0[1287:1280]};
      top_0[1] = {1'b0,layer_1_0[1295:1288]} - {1'b0, layer_0_0[1295:1288]};
      top_0[2] = {1'b0,layer_1_0[1303:1296]} - {1'b0, layer_0_0[1303:1296]};
      top_1[0] = {1'b0,layer_1_1[1287:1280]} - {1'b0, layer_0_1[1287:1280]};
      top_1[1] = {1'b0,layer_1_1[1295:1288]} - {1'b0, layer_0_1[1295:1288]};
      top_1[2] = {1'b0,layer_1_1[1303:1296]} - {1'b0, layer_0_1[1303:1296]};
      top_2[0] = {1'b0,layer_1_2[1287:1280]} - {1'b0, layer_0_2[1287:1280]};
      top_2[1] = {1'b0,layer_1_2[1295:1288]} - {1'b0, layer_0_2[1295:1288]};
      top_2[2] = {1'b0,layer_1_2[1303:1296]} - {1'b0, layer_0_2[1303:1296]};
      mid_0[0] = {1'b0,layer_2_0[1287:1280]} - {1'b0, layer_1_0[1287:1280]};
      mid_0[1] = {1'b0,layer_2_0[1295:1288]} - {1'b0, layer_1_0[1295:1288]};
      mid_0[2] = {1'b0,layer_2_0[1303:1296]} - {1'b0, layer_1_0[1303:1296]};
      mid_1[0] = {1'b0,layer_2_1[1287:1280]} - {1'b0, layer_1_1[1287:1280]};
      mid_1[1] = {1'b0,layer_2_1[1295:1288]} - {1'b0, layer_1_1[1295:1288]};
      mid_1[2] = {1'b0,layer_2_1[1303:1296]} - {1'b0, layer_1_1[1303:1296]};
      mid_2[0] = {1'b0,layer_2_2[1287:1280]} - {1'b0, layer_1_2[1287:1280]};
      mid_2[1] = {1'b0,layer_2_2[1295:1288]} - {1'b0, layer_1_2[1295:1288]};
      mid_2[2] = {1'b0,layer_2_2[1303:1296]} - {1'b0, layer_1_2[1303:1296]};
      btm_0[0] = {1'b0,layer_3_0[1287:1280]} - {1'b0, layer_2_0[1287:1280]};
      btm_0[1] = {1'b0,layer_3_0[1295:1288]} - {1'b0, layer_2_0[1295:1288]};
      btm_0[2] = {1'b0,layer_3_0[1303:1296]} - {1'b0, layer_2_0[1303:1296]};
      btm_1[0] = {1'b0,layer_3_1[1287:1280]} - {1'b0, layer_2_1[1287:1280]};
      btm_1[1] = {1'b0,layer_3_1[1295:1288]} - {1'b0, layer_2_1[1295:1288]};
      btm_1[2] = {1'b0,layer_3_1[1303:1296]} - {1'b0, layer_2_1[1303:1296]};
      btm_2[0] = {1'b0,layer_3_2[1287:1280]} - {1'b0, layer_2_2[1287:1280]};
      btm_2[1] = {1'b0,layer_3_2[1295:1288]} - {1'b0, layer_2_2[1295:1288]};
      btm_2[2] = {1'b0,layer_3_2[1303:1296]} - {1'b0, layer_2_2[1303:1296]};
    end
    'd162: begin
      top_0[0] = {1'b0,layer_1_0[1295:1288]} - {1'b0, layer_0_0[1295:1288]};
      top_0[1] = {1'b0,layer_1_0[1303:1296]} - {1'b0, layer_0_0[1303:1296]};
      top_0[2] = {1'b0,layer_1_0[1311:1304]} - {1'b0, layer_0_0[1311:1304]};
      top_1[0] = {1'b0,layer_1_1[1295:1288]} - {1'b0, layer_0_1[1295:1288]};
      top_1[1] = {1'b0,layer_1_1[1303:1296]} - {1'b0, layer_0_1[1303:1296]};
      top_1[2] = {1'b0,layer_1_1[1311:1304]} - {1'b0, layer_0_1[1311:1304]};
      top_2[0] = {1'b0,layer_1_2[1295:1288]} - {1'b0, layer_0_2[1295:1288]};
      top_2[1] = {1'b0,layer_1_2[1303:1296]} - {1'b0, layer_0_2[1303:1296]};
      top_2[2] = {1'b0,layer_1_2[1311:1304]} - {1'b0, layer_0_2[1311:1304]};
      mid_0[0] = {1'b0,layer_2_0[1295:1288]} - {1'b0, layer_1_0[1295:1288]};
      mid_0[1] = {1'b0,layer_2_0[1303:1296]} - {1'b0, layer_1_0[1303:1296]};
      mid_0[2] = {1'b0,layer_2_0[1311:1304]} - {1'b0, layer_1_0[1311:1304]};
      mid_1[0] = {1'b0,layer_2_1[1295:1288]} - {1'b0, layer_1_1[1295:1288]};
      mid_1[1] = {1'b0,layer_2_1[1303:1296]} - {1'b0, layer_1_1[1303:1296]};
      mid_1[2] = {1'b0,layer_2_1[1311:1304]} - {1'b0, layer_1_1[1311:1304]};
      mid_2[0] = {1'b0,layer_2_2[1295:1288]} - {1'b0, layer_1_2[1295:1288]};
      mid_2[1] = {1'b0,layer_2_2[1303:1296]} - {1'b0, layer_1_2[1303:1296]};
      mid_2[2] = {1'b0,layer_2_2[1311:1304]} - {1'b0, layer_1_2[1311:1304]};
      btm_0[0] = {1'b0,layer_3_0[1295:1288]} - {1'b0, layer_2_0[1295:1288]};
      btm_0[1] = {1'b0,layer_3_0[1303:1296]} - {1'b0, layer_2_0[1303:1296]};
      btm_0[2] = {1'b0,layer_3_0[1311:1304]} - {1'b0, layer_2_0[1311:1304]};
      btm_1[0] = {1'b0,layer_3_1[1295:1288]} - {1'b0, layer_2_1[1295:1288]};
      btm_1[1] = {1'b0,layer_3_1[1303:1296]} - {1'b0, layer_2_1[1303:1296]};
      btm_1[2] = {1'b0,layer_3_1[1311:1304]} - {1'b0, layer_2_1[1311:1304]};
      btm_2[0] = {1'b0,layer_3_2[1295:1288]} - {1'b0, layer_2_2[1295:1288]};
      btm_2[1] = {1'b0,layer_3_2[1303:1296]} - {1'b0, layer_2_2[1303:1296]};
      btm_2[2] = {1'b0,layer_3_2[1311:1304]} - {1'b0, layer_2_2[1311:1304]};
    end
    'd163: begin
      top_0[0] = {1'b0,layer_1_0[1303:1296]} - {1'b0, layer_0_0[1303:1296]};
      top_0[1] = {1'b0,layer_1_0[1311:1304]} - {1'b0, layer_0_0[1311:1304]};
      top_0[2] = {1'b0,layer_1_0[1319:1312]} - {1'b0, layer_0_0[1319:1312]};
      top_1[0] = {1'b0,layer_1_1[1303:1296]} - {1'b0, layer_0_1[1303:1296]};
      top_1[1] = {1'b0,layer_1_1[1311:1304]} - {1'b0, layer_0_1[1311:1304]};
      top_1[2] = {1'b0,layer_1_1[1319:1312]} - {1'b0, layer_0_1[1319:1312]};
      top_2[0] = {1'b0,layer_1_2[1303:1296]} - {1'b0, layer_0_2[1303:1296]};
      top_2[1] = {1'b0,layer_1_2[1311:1304]} - {1'b0, layer_0_2[1311:1304]};
      top_2[2] = {1'b0,layer_1_2[1319:1312]} - {1'b0, layer_0_2[1319:1312]};
      mid_0[0] = {1'b0,layer_2_0[1303:1296]} - {1'b0, layer_1_0[1303:1296]};
      mid_0[1] = {1'b0,layer_2_0[1311:1304]} - {1'b0, layer_1_0[1311:1304]};
      mid_0[2] = {1'b0,layer_2_0[1319:1312]} - {1'b0, layer_1_0[1319:1312]};
      mid_1[0] = {1'b0,layer_2_1[1303:1296]} - {1'b0, layer_1_1[1303:1296]};
      mid_1[1] = {1'b0,layer_2_1[1311:1304]} - {1'b0, layer_1_1[1311:1304]};
      mid_1[2] = {1'b0,layer_2_1[1319:1312]} - {1'b0, layer_1_1[1319:1312]};
      mid_2[0] = {1'b0,layer_2_2[1303:1296]} - {1'b0, layer_1_2[1303:1296]};
      mid_2[1] = {1'b0,layer_2_2[1311:1304]} - {1'b0, layer_1_2[1311:1304]};
      mid_2[2] = {1'b0,layer_2_2[1319:1312]} - {1'b0, layer_1_2[1319:1312]};
      btm_0[0] = {1'b0,layer_3_0[1303:1296]} - {1'b0, layer_2_0[1303:1296]};
      btm_0[1] = {1'b0,layer_3_0[1311:1304]} - {1'b0, layer_2_0[1311:1304]};
      btm_0[2] = {1'b0,layer_3_0[1319:1312]} - {1'b0, layer_2_0[1319:1312]};
      btm_1[0] = {1'b0,layer_3_1[1303:1296]} - {1'b0, layer_2_1[1303:1296]};
      btm_1[1] = {1'b0,layer_3_1[1311:1304]} - {1'b0, layer_2_1[1311:1304]};
      btm_1[2] = {1'b0,layer_3_1[1319:1312]} - {1'b0, layer_2_1[1319:1312]};
      btm_2[0] = {1'b0,layer_3_2[1303:1296]} - {1'b0, layer_2_2[1303:1296]};
      btm_2[1] = {1'b0,layer_3_2[1311:1304]} - {1'b0, layer_2_2[1311:1304]};
      btm_2[2] = {1'b0,layer_3_2[1319:1312]} - {1'b0, layer_2_2[1319:1312]};
    end
    'd164: begin
      top_0[0] = {1'b0,layer_1_0[1311:1304]} - {1'b0, layer_0_0[1311:1304]};
      top_0[1] = {1'b0,layer_1_0[1319:1312]} - {1'b0, layer_0_0[1319:1312]};
      top_0[2] = {1'b0,layer_1_0[1327:1320]} - {1'b0, layer_0_0[1327:1320]};
      top_1[0] = {1'b0,layer_1_1[1311:1304]} - {1'b0, layer_0_1[1311:1304]};
      top_1[1] = {1'b0,layer_1_1[1319:1312]} - {1'b0, layer_0_1[1319:1312]};
      top_1[2] = {1'b0,layer_1_1[1327:1320]} - {1'b0, layer_0_1[1327:1320]};
      top_2[0] = {1'b0,layer_1_2[1311:1304]} - {1'b0, layer_0_2[1311:1304]};
      top_2[1] = {1'b0,layer_1_2[1319:1312]} - {1'b0, layer_0_2[1319:1312]};
      top_2[2] = {1'b0,layer_1_2[1327:1320]} - {1'b0, layer_0_2[1327:1320]};
      mid_0[0] = {1'b0,layer_2_0[1311:1304]} - {1'b0, layer_1_0[1311:1304]};
      mid_0[1] = {1'b0,layer_2_0[1319:1312]} - {1'b0, layer_1_0[1319:1312]};
      mid_0[2] = {1'b0,layer_2_0[1327:1320]} - {1'b0, layer_1_0[1327:1320]};
      mid_1[0] = {1'b0,layer_2_1[1311:1304]} - {1'b0, layer_1_1[1311:1304]};
      mid_1[1] = {1'b0,layer_2_1[1319:1312]} - {1'b0, layer_1_1[1319:1312]};
      mid_1[2] = {1'b0,layer_2_1[1327:1320]} - {1'b0, layer_1_1[1327:1320]};
      mid_2[0] = {1'b0,layer_2_2[1311:1304]} - {1'b0, layer_1_2[1311:1304]};
      mid_2[1] = {1'b0,layer_2_2[1319:1312]} - {1'b0, layer_1_2[1319:1312]};
      mid_2[2] = {1'b0,layer_2_2[1327:1320]} - {1'b0, layer_1_2[1327:1320]};
      btm_0[0] = {1'b0,layer_3_0[1311:1304]} - {1'b0, layer_2_0[1311:1304]};
      btm_0[1] = {1'b0,layer_3_0[1319:1312]} - {1'b0, layer_2_0[1319:1312]};
      btm_0[2] = {1'b0,layer_3_0[1327:1320]} - {1'b0, layer_2_0[1327:1320]};
      btm_1[0] = {1'b0,layer_3_1[1311:1304]} - {1'b0, layer_2_1[1311:1304]};
      btm_1[1] = {1'b0,layer_3_1[1319:1312]} - {1'b0, layer_2_1[1319:1312]};
      btm_1[2] = {1'b0,layer_3_1[1327:1320]} - {1'b0, layer_2_1[1327:1320]};
      btm_2[0] = {1'b0,layer_3_2[1311:1304]} - {1'b0, layer_2_2[1311:1304]};
      btm_2[1] = {1'b0,layer_3_2[1319:1312]} - {1'b0, layer_2_2[1319:1312]};
      btm_2[2] = {1'b0,layer_3_2[1327:1320]} - {1'b0, layer_2_2[1327:1320]};
    end
    'd165: begin
      top_0[0] = {1'b0,layer_1_0[1319:1312]} - {1'b0, layer_0_0[1319:1312]};
      top_0[1] = {1'b0,layer_1_0[1327:1320]} - {1'b0, layer_0_0[1327:1320]};
      top_0[2] = {1'b0,layer_1_0[1335:1328]} - {1'b0, layer_0_0[1335:1328]};
      top_1[0] = {1'b0,layer_1_1[1319:1312]} - {1'b0, layer_0_1[1319:1312]};
      top_1[1] = {1'b0,layer_1_1[1327:1320]} - {1'b0, layer_0_1[1327:1320]};
      top_1[2] = {1'b0,layer_1_1[1335:1328]} - {1'b0, layer_0_1[1335:1328]};
      top_2[0] = {1'b0,layer_1_2[1319:1312]} - {1'b0, layer_0_2[1319:1312]};
      top_2[1] = {1'b0,layer_1_2[1327:1320]} - {1'b0, layer_0_2[1327:1320]};
      top_2[2] = {1'b0,layer_1_2[1335:1328]} - {1'b0, layer_0_2[1335:1328]};
      mid_0[0] = {1'b0,layer_2_0[1319:1312]} - {1'b0, layer_1_0[1319:1312]};
      mid_0[1] = {1'b0,layer_2_0[1327:1320]} - {1'b0, layer_1_0[1327:1320]};
      mid_0[2] = {1'b0,layer_2_0[1335:1328]} - {1'b0, layer_1_0[1335:1328]};
      mid_1[0] = {1'b0,layer_2_1[1319:1312]} - {1'b0, layer_1_1[1319:1312]};
      mid_1[1] = {1'b0,layer_2_1[1327:1320]} - {1'b0, layer_1_1[1327:1320]};
      mid_1[2] = {1'b0,layer_2_1[1335:1328]} - {1'b0, layer_1_1[1335:1328]};
      mid_2[0] = {1'b0,layer_2_2[1319:1312]} - {1'b0, layer_1_2[1319:1312]};
      mid_2[1] = {1'b0,layer_2_2[1327:1320]} - {1'b0, layer_1_2[1327:1320]};
      mid_2[2] = {1'b0,layer_2_2[1335:1328]} - {1'b0, layer_1_2[1335:1328]};
      btm_0[0] = {1'b0,layer_3_0[1319:1312]} - {1'b0, layer_2_0[1319:1312]};
      btm_0[1] = {1'b0,layer_3_0[1327:1320]} - {1'b0, layer_2_0[1327:1320]};
      btm_0[2] = {1'b0,layer_3_0[1335:1328]} - {1'b0, layer_2_0[1335:1328]};
      btm_1[0] = {1'b0,layer_3_1[1319:1312]} - {1'b0, layer_2_1[1319:1312]};
      btm_1[1] = {1'b0,layer_3_1[1327:1320]} - {1'b0, layer_2_1[1327:1320]};
      btm_1[2] = {1'b0,layer_3_1[1335:1328]} - {1'b0, layer_2_1[1335:1328]};
      btm_2[0] = {1'b0,layer_3_2[1319:1312]} - {1'b0, layer_2_2[1319:1312]};
      btm_2[1] = {1'b0,layer_3_2[1327:1320]} - {1'b0, layer_2_2[1327:1320]};
      btm_2[2] = {1'b0,layer_3_2[1335:1328]} - {1'b0, layer_2_2[1335:1328]};
    end
    'd166: begin
      top_0[0] = {1'b0,layer_1_0[1327:1320]} - {1'b0, layer_0_0[1327:1320]};
      top_0[1] = {1'b0,layer_1_0[1335:1328]} - {1'b0, layer_0_0[1335:1328]};
      top_0[2] = {1'b0,layer_1_0[1343:1336]} - {1'b0, layer_0_0[1343:1336]};
      top_1[0] = {1'b0,layer_1_1[1327:1320]} - {1'b0, layer_0_1[1327:1320]};
      top_1[1] = {1'b0,layer_1_1[1335:1328]} - {1'b0, layer_0_1[1335:1328]};
      top_1[2] = {1'b0,layer_1_1[1343:1336]} - {1'b0, layer_0_1[1343:1336]};
      top_2[0] = {1'b0,layer_1_2[1327:1320]} - {1'b0, layer_0_2[1327:1320]};
      top_2[1] = {1'b0,layer_1_2[1335:1328]} - {1'b0, layer_0_2[1335:1328]};
      top_2[2] = {1'b0,layer_1_2[1343:1336]} - {1'b0, layer_0_2[1343:1336]};
      mid_0[0] = {1'b0,layer_2_0[1327:1320]} - {1'b0, layer_1_0[1327:1320]};
      mid_0[1] = {1'b0,layer_2_0[1335:1328]} - {1'b0, layer_1_0[1335:1328]};
      mid_0[2] = {1'b0,layer_2_0[1343:1336]} - {1'b0, layer_1_0[1343:1336]};
      mid_1[0] = {1'b0,layer_2_1[1327:1320]} - {1'b0, layer_1_1[1327:1320]};
      mid_1[1] = {1'b0,layer_2_1[1335:1328]} - {1'b0, layer_1_1[1335:1328]};
      mid_1[2] = {1'b0,layer_2_1[1343:1336]} - {1'b0, layer_1_1[1343:1336]};
      mid_2[0] = {1'b0,layer_2_2[1327:1320]} - {1'b0, layer_1_2[1327:1320]};
      mid_2[1] = {1'b0,layer_2_2[1335:1328]} - {1'b0, layer_1_2[1335:1328]};
      mid_2[2] = {1'b0,layer_2_2[1343:1336]} - {1'b0, layer_1_2[1343:1336]};
      btm_0[0] = {1'b0,layer_3_0[1327:1320]} - {1'b0, layer_2_0[1327:1320]};
      btm_0[1] = {1'b0,layer_3_0[1335:1328]} - {1'b0, layer_2_0[1335:1328]};
      btm_0[2] = {1'b0,layer_3_0[1343:1336]} - {1'b0, layer_2_0[1343:1336]};
      btm_1[0] = {1'b0,layer_3_1[1327:1320]} - {1'b0, layer_2_1[1327:1320]};
      btm_1[1] = {1'b0,layer_3_1[1335:1328]} - {1'b0, layer_2_1[1335:1328]};
      btm_1[2] = {1'b0,layer_3_1[1343:1336]} - {1'b0, layer_2_1[1343:1336]};
      btm_2[0] = {1'b0,layer_3_2[1327:1320]} - {1'b0, layer_2_2[1327:1320]};
      btm_2[1] = {1'b0,layer_3_2[1335:1328]} - {1'b0, layer_2_2[1335:1328]};
      btm_2[2] = {1'b0,layer_3_2[1343:1336]} - {1'b0, layer_2_2[1343:1336]};
    end
    'd167: begin
      top_0[0] = {1'b0,layer_1_0[1335:1328]} - {1'b0, layer_0_0[1335:1328]};
      top_0[1] = {1'b0,layer_1_0[1343:1336]} - {1'b0, layer_0_0[1343:1336]};
      top_0[2] = {1'b0,layer_1_0[1351:1344]} - {1'b0, layer_0_0[1351:1344]};
      top_1[0] = {1'b0,layer_1_1[1335:1328]} - {1'b0, layer_0_1[1335:1328]};
      top_1[1] = {1'b0,layer_1_1[1343:1336]} - {1'b0, layer_0_1[1343:1336]};
      top_1[2] = {1'b0,layer_1_1[1351:1344]} - {1'b0, layer_0_1[1351:1344]};
      top_2[0] = {1'b0,layer_1_2[1335:1328]} - {1'b0, layer_0_2[1335:1328]};
      top_2[1] = {1'b0,layer_1_2[1343:1336]} - {1'b0, layer_0_2[1343:1336]};
      top_2[2] = {1'b0,layer_1_2[1351:1344]} - {1'b0, layer_0_2[1351:1344]};
      mid_0[0] = {1'b0,layer_2_0[1335:1328]} - {1'b0, layer_1_0[1335:1328]};
      mid_0[1] = {1'b0,layer_2_0[1343:1336]} - {1'b0, layer_1_0[1343:1336]};
      mid_0[2] = {1'b0,layer_2_0[1351:1344]} - {1'b0, layer_1_0[1351:1344]};
      mid_1[0] = {1'b0,layer_2_1[1335:1328]} - {1'b0, layer_1_1[1335:1328]};
      mid_1[1] = {1'b0,layer_2_1[1343:1336]} - {1'b0, layer_1_1[1343:1336]};
      mid_1[2] = {1'b0,layer_2_1[1351:1344]} - {1'b0, layer_1_1[1351:1344]};
      mid_2[0] = {1'b0,layer_2_2[1335:1328]} - {1'b0, layer_1_2[1335:1328]};
      mid_2[1] = {1'b0,layer_2_2[1343:1336]} - {1'b0, layer_1_2[1343:1336]};
      mid_2[2] = {1'b0,layer_2_2[1351:1344]} - {1'b0, layer_1_2[1351:1344]};
      btm_0[0] = {1'b0,layer_3_0[1335:1328]} - {1'b0, layer_2_0[1335:1328]};
      btm_0[1] = {1'b0,layer_3_0[1343:1336]} - {1'b0, layer_2_0[1343:1336]};
      btm_0[2] = {1'b0,layer_3_0[1351:1344]} - {1'b0, layer_2_0[1351:1344]};
      btm_1[0] = {1'b0,layer_3_1[1335:1328]} - {1'b0, layer_2_1[1335:1328]};
      btm_1[1] = {1'b0,layer_3_1[1343:1336]} - {1'b0, layer_2_1[1343:1336]};
      btm_1[2] = {1'b0,layer_3_1[1351:1344]} - {1'b0, layer_2_1[1351:1344]};
      btm_2[0] = {1'b0,layer_3_2[1335:1328]} - {1'b0, layer_2_2[1335:1328]};
      btm_2[1] = {1'b0,layer_3_2[1343:1336]} - {1'b0, layer_2_2[1343:1336]};
      btm_2[2] = {1'b0,layer_3_2[1351:1344]} - {1'b0, layer_2_2[1351:1344]};
    end
    'd168: begin
      top_0[0] = {1'b0,layer_1_0[1343:1336]} - {1'b0, layer_0_0[1343:1336]};
      top_0[1] = {1'b0,layer_1_0[1351:1344]} - {1'b0, layer_0_0[1351:1344]};
      top_0[2] = {1'b0,layer_1_0[1359:1352]} - {1'b0, layer_0_0[1359:1352]};
      top_1[0] = {1'b0,layer_1_1[1343:1336]} - {1'b0, layer_0_1[1343:1336]};
      top_1[1] = {1'b0,layer_1_1[1351:1344]} - {1'b0, layer_0_1[1351:1344]};
      top_1[2] = {1'b0,layer_1_1[1359:1352]} - {1'b0, layer_0_1[1359:1352]};
      top_2[0] = {1'b0,layer_1_2[1343:1336]} - {1'b0, layer_0_2[1343:1336]};
      top_2[1] = {1'b0,layer_1_2[1351:1344]} - {1'b0, layer_0_2[1351:1344]};
      top_2[2] = {1'b0,layer_1_2[1359:1352]} - {1'b0, layer_0_2[1359:1352]};
      mid_0[0] = {1'b0,layer_2_0[1343:1336]} - {1'b0, layer_1_0[1343:1336]};
      mid_0[1] = {1'b0,layer_2_0[1351:1344]} - {1'b0, layer_1_0[1351:1344]};
      mid_0[2] = {1'b0,layer_2_0[1359:1352]} - {1'b0, layer_1_0[1359:1352]};
      mid_1[0] = {1'b0,layer_2_1[1343:1336]} - {1'b0, layer_1_1[1343:1336]};
      mid_1[1] = {1'b0,layer_2_1[1351:1344]} - {1'b0, layer_1_1[1351:1344]};
      mid_1[2] = {1'b0,layer_2_1[1359:1352]} - {1'b0, layer_1_1[1359:1352]};
      mid_2[0] = {1'b0,layer_2_2[1343:1336]} - {1'b0, layer_1_2[1343:1336]};
      mid_2[1] = {1'b0,layer_2_2[1351:1344]} - {1'b0, layer_1_2[1351:1344]};
      mid_2[2] = {1'b0,layer_2_2[1359:1352]} - {1'b0, layer_1_2[1359:1352]};
      btm_0[0] = {1'b0,layer_3_0[1343:1336]} - {1'b0, layer_2_0[1343:1336]};
      btm_0[1] = {1'b0,layer_3_0[1351:1344]} - {1'b0, layer_2_0[1351:1344]};
      btm_0[2] = {1'b0,layer_3_0[1359:1352]} - {1'b0, layer_2_0[1359:1352]};
      btm_1[0] = {1'b0,layer_3_1[1343:1336]} - {1'b0, layer_2_1[1343:1336]};
      btm_1[1] = {1'b0,layer_3_1[1351:1344]} - {1'b0, layer_2_1[1351:1344]};
      btm_1[2] = {1'b0,layer_3_1[1359:1352]} - {1'b0, layer_2_1[1359:1352]};
      btm_2[0] = {1'b0,layer_3_2[1343:1336]} - {1'b0, layer_2_2[1343:1336]};
      btm_2[1] = {1'b0,layer_3_2[1351:1344]} - {1'b0, layer_2_2[1351:1344]};
      btm_2[2] = {1'b0,layer_3_2[1359:1352]} - {1'b0, layer_2_2[1359:1352]};
    end
    'd169: begin
      top_0[0] = {1'b0,layer_1_0[1351:1344]} - {1'b0, layer_0_0[1351:1344]};
      top_0[1] = {1'b0,layer_1_0[1359:1352]} - {1'b0, layer_0_0[1359:1352]};
      top_0[2] = {1'b0,layer_1_0[1367:1360]} - {1'b0, layer_0_0[1367:1360]};
      top_1[0] = {1'b0,layer_1_1[1351:1344]} - {1'b0, layer_0_1[1351:1344]};
      top_1[1] = {1'b0,layer_1_1[1359:1352]} - {1'b0, layer_0_1[1359:1352]};
      top_1[2] = {1'b0,layer_1_1[1367:1360]} - {1'b0, layer_0_1[1367:1360]};
      top_2[0] = {1'b0,layer_1_2[1351:1344]} - {1'b0, layer_0_2[1351:1344]};
      top_2[1] = {1'b0,layer_1_2[1359:1352]} - {1'b0, layer_0_2[1359:1352]};
      top_2[2] = {1'b0,layer_1_2[1367:1360]} - {1'b0, layer_0_2[1367:1360]};
      mid_0[0] = {1'b0,layer_2_0[1351:1344]} - {1'b0, layer_1_0[1351:1344]};
      mid_0[1] = {1'b0,layer_2_0[1359:1352]} - {1'b0, layer_1_0[1359:1352]};
      mid_0[2] = {1'b0,layer_2_0[1367:1360]} - {1'b0, layer_1_0[1367:1360]};
      mid_1[0] = {1'b0,layer_2_1[1351:1344]} - {1'b0, layer_1_1[1351:1344]};
      mid_1[1] = {1'b0,layer_2_1[1359:1352]} - {1'b0, layer_1_1[1359:1352]};
      mid_1[2] = {1'b0,layer_2_1[1367:1360]} - {1'b0, layer_1_1[1367:1360]};
      mid_2[0] = {1'b0,layer_2_2[1351:1344]} - {1'b0, layer_1_2[1351:1344]};
      mid_2[1] = {1'b0,layer_2_2[1359:1352]} - {1'b0, layer_1_2[1359:1352]};
      mid_2[2] = {1'b0,layer_2_2[1367:1360]} - {1'b0, layer_1_2[1367:1360]};
      btm_0[0] = {1'b0,layer_3_0[1351:1344]} - {1'b0, layer_2_0[1351:1344]};
      btm_0[1] = {1'b0,layer_3_0[1359:1352]} - {1'b0, layer_2_0[1359:1352]};
      btm_0[2] = {1'b0,layer_3_0[1367:1360]} - {1'b0, layer_2_0[1367:1360]};
      btm_1[0] = {1'b0,layer_3_1[1351:1344]} - {1'b0, layer_2_1[1351:1344]};
      btm_1[1] = {1'b0,layer_3_1[1359:1352]} - {1'b0, layer_2_1[1359:1352]};
      btm_1[2] = {1'b0,layer_3_1[1367:1360]} - {1'b0, layer_2_1[1367:1360]};
      btm_2[0] = {1'b0,layer_3_2[1351:1344]} - {1'b0, layer_2_2[1351:1344]};
      btm_2[1] = {1'b0,layer_3_2[1359:1352]} - {1'b0, layer_2_2[1359:1352]};
      btm_2[2] = {1'b0,layer_3_2[1367:1360]} - {1'b0, layer_2_2[1367:1360]};
    end
    'd170: begin
      top_0[0] = {1'b0,layer_1_0[1359:1352]} - {1'b0, layer_0_0[1359:1352]};
      top_0[1] = {1'b0,layer_1_0[1367:1360]} - {1'b0, layer_0_0[1367:1360]};
      top_0[2] = {1'b0,layer_1_0[1375:1368]} - {1'b0, layer_0_0[1375:1368]};
      top_1[0] = {1'b0,layer_1_1[1359:1352]} - {1'b0, layer_0_1[1359:1352]};
      top_1[1] = {1'b0,layer_1_1[1367:1360]} - {1'b0, layer_0_1[1367:1360]};
      top_1[2] = {1'b0,layer_1_1[1375:1368]} - {1'b0, layer_0_1[1375:1368]};
      top_2[0] = {1'b0,layer_1_2[1359:1352]} - {1'b0, layer_0_2[1359:1352]};
      top_2[1] = {1'b0,layer_1_2[1367:1360]} - {1'b0, layer_0_2[1367:1360]};
      top_2[2] = {1'b0,layer_1_2[1375:1368]} - {1'b0, layer_0_2[1375:1368]};
      mid_0[0] = {1'b0,layer_2_0[1359:1352]} - {1'b0, layer_1_0[1359:1352]};
      mid_0[1] = {1'b0,layer_2_0[1367:1360]} - {1'b0, layer_1_0[1367:1360]};
      mid_0[2] = {1'b0,layer_2_0[1375:1368]} - {1'b0, layer_1_0[1375:1368]};
      mid_1[0] = {1'b0,layer_2_1[1359:1352]} - {1'b0, layer_1_1[1359:1352]};
      mid_1[1] = {1'b0,layer_2_1[1367:1360]} - {1'b0, layer_1_1[1367:1360]};
      mid_1[2] = {1'b0,layer_2_1[1375:1368]} - {1'b0, layer_1_1[1375:1368]};
      mid_2[0] = {1'b0,layer_2_2[1359:1352]} - {1'b0, layer_1_2[1359:1352]};
      mid_2[1] = {1'b0,layer_2_2[1367:1360]} - {1'b0, layer_1_2[1367:1360]};
      mid_2[2] = {1'b0,layer_2_2[1375:1368]} - {1'b0, layer_1_2[1375:1368]};
      btm_0[0] = {1'b0,layer_3_0[1359:1352]} - {1'b0, layer_2_0[1359:1352]};
      btm_0[1] = {1'b0,layer_3_0[1367:1360]} - {1'b0, layer_2_0[1367:1360]};
      btm_0[2] = {1'b0,layer_3_0[1375:1368]} - {1'b0, layer_2_0[1375:1368]};
      btm_1[0] = {1'b0,layer_3_1[1359:1352]} - {1'b0, layer_2_1[1359:1352]};
      btm_1[1] = {1'b0,layer_3_1[1367:1360]} - {1'b0, layer_2_1[1367:1360]};
      btm_1[2] = {1'b0,layer_3_1[1375:1368]} - {1'b0, layer_2_1[1375:1368]};
      btm_2[0] = {1'b0,layer_3_2[1359:1352]} - {1'b0, layer_2_2[1359:1352]};
      btm_2[1] = {1'b0,layer_3_2[1367:1360]} - {1'b0, layer_2_2[1367:1360]};
      btm_2[2] = {1'b0,layer_3_2[1375:1368]} - {1'b0, layer_2_2[1375:1368]};
    end
    'd171: begin
      top_0[0] = {1'b0,layer_1_0[1367:1360]} - {1'b0, layer_0_0[1367:1360]};
      top_0[1] = {1'b0,layer_1_0[1375:1368]} - {1'b0, layer_0_0[1375:1368]};
      top_0[2] = {1'b0,layer_1_0[1383:1376]} - {1'b0, layer_0_0[1383:1376]};
      top_1[0] = {1'b0,layer_1_1[1367:1360]} - {1'b0, layer_0_1[1367:1360]};
      top_1[1] = {1'b0,layer_1_1[1375:1368]} - {1'b0, layer_0_1[1375:1368]};
      top_1[2] = {1'b0,layer_1_1[1383:1376]} - {1'b0, layer_0_1[1383:1376]};
      top_2[0] = {1'b0,layer_1_2[1367:1360]} - {1'b0, layer_0_2[1367:1360]};
      top_2[1] = {1'b0,layer_1_2[1375:1368]} - {1'b0, layer_0_2[1375:1368]};
      top_2[2] = {1'b0,layer_1_2[1383:1376]} - {1'b0, layer_0_2[1383:1376]};
      mid_0[0] = {1'b0,layer_2_0[1367:1360]} - {1'b0, layer_1_0[1367:1360]};
      mid_0[1] = {1'b0,layer_2_0[1375:1368]} - {1'b0, layer_1_0[1375:1368]};
      mid_0[2] = {1'b0,layer_2_0[1383:1376]} - {1'b0, layer_1_0[1383:1376]};
      mid_1[0] = {1'b0,layer_2_1[1367:1360]} - {1'b0, layer_1_1[1367:1360]};
      mid_1[1] = {1'b0,layer_2_1[1375:1368]} - {1'b0, layer_1_1[1375:1368]};
      mid_1[2] = {1'b0,layer_2_1[1383:1376]} - {1'b0, layer_1_1[1383:1376]};
      mid_2[0] = {1'b0,layer_2_2[1367:1360]} - {1'b0, layer_1_2[1367:1360]};
      mid_2[1] = {1'b0,layer_2_2[1375:1368]} - {1'b0, layer_1_2[1375:1368]};
      mid_2[2] = {1'b0,layer_2_2[1383:1376]} - {1'b0, layer_1_2[1383:1376]};
      btm_0[0] = {1'b0,layer_3_0[1367:1360]} - {1'b0, layer_2_0[1367:1360]};
      btm_0[1] = {1'b0,layer_3_0[1375:1368]} - {1'b0, layer_2_0[1375:1368]};
      btm_0[2] = {1'b0,layer_3_0[1383:1376]} - {1'b0, layer_2_0[1383:1376]};
      btm_1[0] = {1'b0,layer_3_1[1367:1360]} - {1'b0, layer_2_1[1367:1360]};
      btm_1[1] = {1'b0,layer_3_1[1375:1368]} - {1'b0, layer_2_1[1375:1368]};
      btm_1[2] = {1'b0,layer_3_1[1383:1376]} - {1'b0, layer_2_1[1383:1376]};
      btm_2[0] = {1'b0,layer_3_2[1367:1360]} - {1'b0, layer_2_2[1367:1360]};
      btm_2[1] = {1'b0,layer_3_2[1375:1368]} - {1'b0, layer_2_2[1375:1368]};
      btm_2[2] = {1'b0,layer_3_2[1383:1376]} - {1'b0, layer_2_2[1383:1376]};
    end
    'd172: begin
      top_0[0] = {1'b0,layer_1_0[1375:1368]} - {1'b0, layer_0_0[1375:1368]};
      top_0[1] = {1'b0,layer_1_0[1383:1376]} - {1'b0, layer_0_0[1383:1376]};
      top_0[2] = {1'b0,layer_1_0[1391:1384]} - {1'b0, layer_0_0[1391:1384]};
      top_1[0] = {1'b0,layer_1_1[1375:1368]} - {1'b0, layer_0_1[1375:1368]};
      top_1[1] = {1'b0,layer_1_1[1383:1376]} - {1'b0, layer_0_1[1383:1376]};
      top_1[2] = {1'b0,layer_1_1[1391:1384]} - {1'b0, layer_0_1[1391:1384]};
      top_2[0] = {1'b0,layer_1_2[1375:1368]} - {1'b0, layer_0_2[1375:1368]};
      top_2[1] = {1'b0,layer_1_2[1383:1376]} - {1'b0, layer_0_2[1383:1376]};
      top_2[2] = {1'b0,layer_1_2[1391:1384]} - {1'b0, layer_0_2[1391:1384]};
      mid_0[0] = {1'b0,layer_2_0[1375:1368]} - {1'b0, layer_1_0[1375:1368]};
      mid_0[1] = {1'b0,layer_2_0[1383:1376]} - {1'b0, layer_1_0[1383:1376]};
      mid_0[2] = {1'b0,layer_2_0[1391:1384]} - {1'b0, layer_1_0[1391:1384]};
      mid_1[0] = {1'b0,layer_2_1[1375:1368]} - {1'b0, layer_1_1[1375:1368]};
      mid_1[1] = {1'b0,layer_2_1[1383:1376]} - {1'b0, layer_1_1[1383:1376]};
      mid_1[2] = {1'b0,layer_2_1[1391:1384]} - {1'b0, layer_1_1[1391:1384]};
      mid_2[0] = {1'b0,layer_2_2[1375:1368]} - {1'b0, layer_1_2[1375:1368]};
      mid_2[1] = {1'b0,layer_2_2[1383:1376]} - {1'b0, layer_1_2[1383:1376]};
      mid_2[2] = {1'b0,layer_2_2[1391:1384]} - {1'b0, layer_1_2[1391:1384]};
      btm_0[0] = {1'b0,layer_3_0[1375:1368]} - {1'b0, layer_2_0[1375:1368]};
      btm_0[1] = {1'b0,layer_3_0[1383:1376]} - {1'b0, layer_2_0[1383:1376]};
      btm_0[2] = {1'b0,layer_3_0[1391:1384]} - {1'b0, layer_2_0[1391:1384]};
      btm_1[0] = {1'b0,layer_3_1[1375:1368]} - {1'b0, layer_2_1[1375:1368]};
      btm_1[1] = {1'b0,layer_3_1[1383:1376]} - {1'b0, layer_2_1[1383:1376]};
      btm_1[2] = {1'b0,layer_3_1[1391:1384]} - {1'b0, layer_2_1[1391:1384]};
      btm_2[0] = {1'b0,layer_3_2[1375:1368]} - {1'b0, layer_2_2[1375:1368]};
      btm_2[1] = {1'b0,layer_3_2[1383:1376]} - {1'b0, layer_2_2[1383:1376]};
      btm_2[2] = {1'b0,layer_3_2[1391:1384]} - {1'b0, layer_2_2[1391:1384]};
    end
    'd173: begin
      top_0[0] = {1'b0,layer_1_0[1383:1376]} - {1'b0, layer_0_0[1383:1376]};
      top_0[1] = {1'b0,layer_1_0[1391:1384]} - {1'b0, layer_0_0[1391:1384]};
      top_0[2] = {1'b0,layer_1_0[1399:1392]} - {1'b0, layer_0_0[1399:1392]};
      top_1[0] = {1'b0,layer_1_1[1383:1376]} - {1'b0, layer_0_1[1383:1376]};
      top_1[1] = {1'b0,layer_1_1[1391:1384]} - {1'b0, layer_0_1[1391:1384]};
      top_1[2] = {1'b0,layer_1_1[1399:1392]} - {1'b0, layer_0_1[1399:1392]};
      top_2[0] = {1'b0,layer_1_2[1383:1376]} - {1'b0, layer_0_2[1383:1376]};
      top_2[1] = {1'b0,layer_1_2[1391:1384]} - {1'b0, layer_0_2[1391:1384]};
      top_2[2] = {1'b0,layer_1_2[1399:1392]} - {1'b0, layer_0_2[1399:1392]};
      mid_0[0] = {1'b0,layer_2_0[1383:1376]} - {1'b0, layer_1_0[1383:1376]};
      mid_0[1] = {1'b0,layer_2_0[1391:1384]} - {1'b0, layer_1_0[1391:1384]};
      mid_0[2] = {1'b0,layer_2_0[1399:1392]} - {1'b0, layer_1_0[1399:1392]};
      mid_1[0] = {1'b0,layer_2_1[1383:1376]} - {1'b0, layer_1_1[1383:1376]};
      mid_1[1] = {1'b0,layer_2_1[1391:1384]} - {1'b0, layer_1_1[1391:1384]};
      mid_1[2] = {1'b0,layer_2_1[1399:1392]} - {1'b0, layer_1_1[1399:1392]};
      mid_2[0] = {1'b0,layer_2_2[1383:1376]} - {1'b0, layer_1_2[1383:1376]};
      mid_2[1] = {1'b0,layer_2_2[1391:1384]} - {1'b0, layer_1_2[1391:1384]};
      mid_2[2] = {1'b0,layer_2_2[1399:1392]} - {1'b0, layer_1_2[1399:1392]};
      btm_0[0] = {1'b0,layer_3_0[1383:1376]} - {1'b0, layer_2_0[1383:1376]};
      btm_0[1] = {1'b0,layer_3_0[1391:1384]} - {1'b0, layer_2_0[1391:1384]};
      btm_0[2] = {1'b0,layer_3_0[1399:1392]} - {1'b0, layer_2_0[1399:1392]};
      btm_1[0] = {1'b0,layer_3_1[1383:1376]} - {1'b0, layer_2_1[1383:1376]};
      btm_1[1] = {1'b0,layer_3_1[1391:1384]} - {1'b0, layer_2_1[1391:1384]};
      btm_1[2] = {1'b0,layer_3_1[1399:1392]} - {1'b0, layer_2_1[1399:1392]};
      btm_2[0] = {1'b0,layer_3_2[1383:1376]} - {1'b0, layer_2_2[1383:1376]};
      btm_2[1] = {1'b0,layer_3_2[1391:1384]} - {1'b0, layer_2_2[1391:1384]};
      btm_2[2] = {1'b0,layer_3_2[1399:1392]} - {1'b0, layer_2_2[1399:1392]};
    end
    'd174: begin
      top_0[0] = {1'b0,layer_1_0[1391:1384]} - {1'b0, layer_0_0[1391:1384]};
      top_0[1] = {1'b0,layer_1_0[1399:1392]} - {1'b0, layer_0_0[1399:1392]};
      top_0[2] = {1'b0,layer_1_0[1407:1400]} - {1'b0, layer_0_0[1407:1400]};
      top_1[0] = {1'b0,layer_1_1[1391:1384]} - {1'b0, layer_0_1[1391:1384]};
      top_1[1] = {1'b0,layer_1_1[1399:1392]} - {1'b0, layer_0_1[1399:1392]};
      top_1[2] = {1'b0,layer_1_1[1407:1400]} - {1'b0, layer_0_1[1407:1400]};
      top_2[0] = {1'b0,layer_1_2[1391:1384]} - {1'b0, layer_0_2[1391:1384]};
      top_2[1] = {1'b0,layer_1_2[1399:1392]} - {1'b0, layer_0_2[1399:1392]};
      top_2[2] = {1'b0,layer_1_2[1407:1400]} - {1'b0, layer_0_2[1407:1400]};
      mid_0[0] = {1'b0,layer_2_0[1391:1384]} - {1'b0, layer_1_0[1391:1384]};
      mid_0[1] = {1'b0,layer_2_0[1399:1392]} - {1'b0, layer_1_0[1399:1392]};
      mid_0[2] = {1'b0,layer_2_0[1407:1400]} - {1'b0, layer_1_0[1407:1400]};
      mid_1[0] = {1'b0,layer_2_1[1391:1384]} - {1'b0, layer_1_1[1391:1384]};
      mid_1[1] = {1'b0,layer_2_1[1399:1392]} - {1'b0, layer_1_1[1399:1392]};
      mid_1[2] = {1'b0,layer_2_1[1407:1400]} - {1'b0, layer_1_1[1407:1400]};
      mid_2[0] = {1'b0,layer_2_2[1391:1384]} - {1'b0, layer_1_2[1391:1384]};
      mid_2[1] = {1'b0,layer_2_2[1399:1392]} - {1'b0, layer_1_2[1399:1392]};
      mid_2[2] = {1'b0,layer_2_2[1407:1400]} - {1'b0, layer_1_2[1407:1400]};
      btm_0[0] = {1'b0,layer_3_0[1391:1384]} - {1'b0, layer_2_0[1391:1384]};
      btm_0[1] = {1'b0,layer_3_0[1399:1392]} - {1'b0, layer_2_0[1399:1392]};
      btm_0[2] = {1'b0,layer_3_0[1407:1400]} - {1'b0, layer_2_0[1407:1400]};
      btm_1[0] = {1'b0,layer_3_1[1391:1384]} - {1'b0, layer_2_1[1391:1384]};
      btm_1[1] = {1'b0,layer_3_1[1399:1392]} - {1'b0, layer_2_1[1399:1392]};
      btm_1[2] = {1'b0,layer_3_1[1407:1400]} - {1'b0, layer_2_1[1407:1400]};
      btm_2[0] = {1'b0,layer_3_2[1391:1384]} - {1'b0, layer_2_2[1391:1384]};
      btm_2[1] = {1'b0,layer_3_2[1399:1392]} - {1'b0, layer_2_2[1399:1392]};
      btm_2[2] = {1'b0,layer_3_2[1407:1400]} - {1'b0, layer_2_2[1407:1400]};
    end
    'd175: begin
      top_0[0] = {1'b0,layer_1_0[1399:1392]} - {1'b0, layer_0_0[1399:1392]};
      top_0[1] = {1'b0,layer_1_0[1407:1400]} - {1'b0, layer_0_0[1407:1400]};
      top_0[2] = {1'b0,layer_1_0[1415:1408]} - {1'b0, layer_0_0[1415:1408]};
      top_1[0] = {1'b0,layer_1_1[1399:1392]} - {1'b0, layer_0_1[1399:1392]};
      top_1[1] = {1'b0,layer_1_1[1407:1400]} - {1'b0, layer_0_1[1407:1400]};
      top_1[2] = {1'b0,layer_1_1[1415:1408]} - {1'b0, layer_0_1[1415:1408]};
      top_2[0] = {1'b0,layer_1_2[1399:1392]} - {1'b0, layer_0_2[1399:1392]};
      top_2[1] = {1'b0,layer_1_2[1407:1400]} - {1'b0, layer_0_2[1407:1400]};
      top_2[2] = {1'b0,layer_1_2[1415:1408]} - {1'b0, layer_0_2[1415:1408]};
      mid_0[0] = {1'b0,layer_2_0[1399:1392]} - {1'b0, layer_1_0[1399:1392]};
      mid_0[1] = {1'b0,layer_2_0[1407:1400]} - {1'b0, layer_1_0[1407:1400]};
      mid_0[2] = {1'b0,layer_2_0[1415:1408]} - {1'b0, layer_1_0[1415:1408]};
      mid_1[0] = {1'b0,layer_2_1[1399:1392]} - {1'b0, layer_1_1[1399:1392]};
      mid_1[1] = {1'b0,layer_2_1[1407:1400]} - {1'b0, layer_1_1[1407:1400]};
      mid_1[2] = {1'b0,layer_2_1[1415:1408]} - {1'b0, layer_1_1[1415:1408]};
      mid_2[0] = {1'b0,layer_2_2[1399:1392]} - {1'b0, layer_1_2[1399:1392]};
      mid_2[1] = {1'b0,layer_2_2[1407:1400]} - {1'b0, layer_1_2[1407:1400]};
      mid_2[2] = {1'b0,layer_2_2[1415:1408]} - {1'b0, layer_1_2[1415:1408]};
      btm_0[0] = {1'b0,layer_3_0[1399:1392]} - {1'b0, layer_2_0[1399:1392]};
      btm_0[1] = {1'b0,layer_3_0[1407:1400]} - {1'b0, layer_2_0[1407:1400]};
      btm_0[2] = {1'b0,layer_3_0[1415:1408]} - {1'b0, layer_2_0[1415:1408]};
      btm_1[0] = {1'b0,layer_3_1[1399:1392]} - {1'b0, layer_2_1[1399:1392]};
      btm_1[1] = {1'b0,layer_3_1[1407:1400]} - {1'b0, layer_2_1[1407:1400]};
      btm_1[2] = {1'b0,layer_3_1[1415:1408]} - {1'b0, layer_2_1[1415:1408]};
      btm_2[0] = {1'b0,layer_3_2[1399:1392]} - {1'b0, layer_2_2[1399:1392]};
      btm_2[1] = {1'b0,layer_3_2[1407:1400]} - {1'b0, layer_2_2[1407:1400]};
      btm_2[2] = {1'b0,layer_3_2[1415:1408]} - {1'b0, layer_2_2[1415:1408]};
    end
    'd176: begin
      top_0[0] = {1'b0,layer_1_0[1407:1400]} - {1'b0, layer_0_0[1407:1400]};
      top_0[1] = {1'b0,layer_1_0[1415:1408]} - {1'b0, layer_0_0[1415:1408]};
      top_0[2] = {1'b0,layer_1_0[1423:1416]} - {1'b0, layer_0_0[1423:1416]};
      top_1[0] = {1'b0,layer_1_1[1407:1400]} - {1'b0, layer_0_1[1407:1400]};
      top_1[1] = {1'b0,layer_1_1[1415:1408]} - {1'b0, layer_0_1[1415:1408]};
      top_1[2] = {1'b0,layer_1_1[1423:1416]} - {1'b0, layer_0_1[1423:1416]};
      top_2[0] = {1'b0,layer_1_2[1407:1400]} - {1'b0, layer_0_2[1407:1400]};
      top_2[1] = {1'b0,layer_1_2[1415:1408]} - {1'b0, layer_0_2[1415:1408]};
      top_2[2] = {1'b0,layer_1_2[1423:1416]} - {1'b0, layer_0_2[1423:1416]};
      mid_0[0] = {1'b0,layer_2_0[1407:1400]} - {1'b0, layer_1_0[1407:1400]};
      mid_0[1] = {1'b0,layer_2_0[1415:1408]} - {1'b0, layer_1_0[1415:1408]};
      mid_0[2] = {1'b0,layer_2_0[1423:1416]} - {1'b0, layer_1_0[1423:1416]};
      mid_1[0] = {1'b0,layer_2_1[1407:1400]} - {1'b0, layer_1_1[1407:1400]};
      mid_1[1] = {1'b0,layer_2_1[1415:1408]} - {1'b0, layer_1_1[1415:1408]};
      mid_1[2] = {1'b0,layer_2_1[1423:1416]} - {1'b0, layer_1_1[1423:1416]};
      mid_2[0] = {1'b0,layer_2_2[1407:1400]} - {1'b0, layer_1_2[1407:1400]};
      mid_2[1] = {1'b0,layer_2_2[1415:1408]} - {1'b0, layer_1_2[1415:1408]};
      mid_2[2] = {1'b0,layer_2_2[1423:1416]} - {1'b0, layer_1_2[1423:1416]};
      btm_0[0] = {1'b0,layer_3_0[1407:1400]} - {1'b0, layer_2_0[1407:1400]};
      btm_0[1] = {1'b0,layer_3_0[1415:1408]} - {1'b0, layer_2_0[1415:1408]};
      btm_0[2] = {1'b0,layer_3_0[1423:1416]} - {1'b0, layer_2_0[1423:1416]};
      btm_1[0] = {1'b0,layer_3_1[1407:1400]} - {1'b0, layer_2_1[1407:1400]};
      btm_1[1] = {1'b0,layer_3_1[1415:1408]} - {1'b0, layer_2_1[1415:1408]};
      btm_1[2] = {1'b0,layer_3_1[1423:1416]} - {1'b0, layer_2_1[1423:1416]};
      btm_2[0] = {1'b0,layer_3_2[1407:1400]} - {1'b0, layer_2_2[1407:1400]};
      btm_2[1] = {1'b0,layer_3_2[1415:1408]} - {1'b0, layer_2_2[1415:1408]};
      btm_2[2] = {1'b0,layer_3_2[1423:1416]} - {1'b0, layer_2_2[1423:1416]};
    end
    'd177: begin
      top_0[0] = {1'b0,layer_1_0[1415:1408]} - {1'b0, layer_0_0[1415:1408]};
      top_0[1] = {1'b0,layer_1_0[1423:1416]} - {1'b0, layer_0_0[1423:1416]};
      top_0[2] = {1'b0,layer_1_0[1431:1424]} - {1'b0, layer_0_0[1431:1424]};
      top_1[0] = {1'b0,layer_1_1[1415:1408]} - {1'b0, layer_0_1[1415:1408]};
      top_1[1] = {1'b0,layer_1_1[1423:1416]} - {1'b0, layer_0_1[1423:1416]};
      top_1[2] = {1'b0,layer_1_1[1431:1424]} - {1'b0, layer_0_1[1431:1424]};
      top_2[0] = {1'b0,layer_1_2[1415:1408]} - {1'b0, layer_0_2[1415:1408]};
      top_2[1] = {1'b0,layer_1_2[1423:1416]} - {1'b0, layer_0_2[1423:1416]};
      top_2[2] = {1'b0,layer_1_2[1431:1424]} - {1'b0, layer_0_2[1431:1424]};
      mid_0[0] = {1'b0,layer_2_0[1415:1408]} - {1'b0, layer_1_0[1415:1408]};
      mid_0[1] = {1'b0,layer_2_0[1423:1416]} - {1'b0, layer_1_0[1423:1416]};
      mid_0[2] = {1'b0,layer_2_0[1431:1424]} - {1'b0, layer_1_0[1431:1424]};
      mid_1[0] = {1'b0,layer_2_1[1415:1408]} - {1'b0, layer_1_1[1415:1408]};
      mid_1[1] = {1'b0,layer_2_1[1423:1416]} - {1'b0, layer_1_1[1423:1416]};
      mid_1[2] = {1'b0,layer_2_1[1431:1424]} - {1'b0, layer_1_1[1431:1424]};
      mid_2[0] = {1'b0,layer_2_2[1415:1408]} - {1'b0, layer_1_2[1415:1408]};
      mid_2[1] = {1'b0,layer_2_2[1423:1416]} - {1'b0, layer_1_2[1423:1416]};
      mid_2[2] = {1'b0,layer_2_2[1431:1424]} - {1'b0, layer_1_2[1431:1424]};
      btm_0[0] = {1'b0,layer_3_0[1415:1408]} - {1'b0, layer_2_0[1415:1408]};
      btm_0[1] = {1'b0,layer_3_0[1423:1416]} - {1'b0, layer_2_0[1423:1416]};
      btm_0[2] = {1'b0,layer_3_0[1431:1424]} - {1'b0, layer_2_0[1431:1424]};
      btm_1[0] = {1'b0,layer_3_1[1415:1408]} - {1'b0, layer_2_1[1415:1408]};
      btm_1[1] = {1'b0,layer_3_1[1423:1416]} - {1'b0, layer_2_1[1423:1416]};
      btm_1[2] = {1'b0,layer_3_1[1431:1424]} - {1'b0, layer_2_1[1431:1424]};
      btm_2[0] = {1'b0,layer_3_2[1415:1408]} - {1'b0, layer_2_2[1415:1408]};
      btm_2[1] = {1'b0,layer_3_2[1423:1416]} - {1'b0, layer_2_2[1423:1416]};
      btm_2[2] = {1'b0,layer_3_2[1431:1424]} - {1'b0, layer_2_2[1431:1424]};
    end
    'd178: begin
      top_0[0] = {1'b0,layer_1_0[1423:1416]} - {1'b0, layer_0_0[1423:1416]};
      top_0[1] = {1'b0,layer_1_0[1431:1424]} - {1'b0, layer_0_0[1431:1424]};
      top_0[2] = {1'b0,layer_1_0[1439:1432]} - {1'b0, layer_0_0[1439:1432]};
      top_1[0] = {1'b0,layer_1_1[1423:1416]} - {1'b0, layer_0_1[1423:1416]};
      top_1[1] = {1'b0,layer_1_1[1431:1424]} - {1'b0, layer_0_1[1431:1424]};
      top_1[2] = {1'b0,layer_1_1[1439:1432]} - {1'b0, layer_0_1[1439:1432]};
      top_2[0] = {1'b0,layer_1_2[1423:1416]} - {1'b0, layer_0_2[1423:1416]};
      top_2[1] = {1'b0,layer_1_2[1431:1424]} - {1'b0, layer_0_2[1431:1424]};
      top_2[2] = {1'b0,layer_1_2[1439:1432]} - {1'b0, layer_0_2[1439:1432]};
      mid_0[0] = {1'b0,layer_2_0[1423:1416]} - {1'b0, layer_1_0[1423:1416]};
      mid_0[1] = {1'b0,layer_2_0[1431:1424]} - {1'b0, layer_1_0[1431:1424]};
      mid_0[2] = {1'b0,layer_2_0[1439:1432]} - {1'b0, layer_1_0[1439:1432]};
      mid_1[0] = {1'b0,layer_2_1[1423:1416]} - {1'b0, layer_1_1[1423:1416]};
      mid_1[1] = {1'b0,layer_2_1[1431:1424]} - {1'b0, layer_1_1[1431:1424]};
      mid_1[2] = {1'b0,layer_2_1[1439:1432]} - {1'b0, layer_1_1[1439:1432]};
      mid_2[0] = {1'b0,layer_2_2[1423:1416]} - {1'b0, layer_1_2[1423:1416]};
      mid_2[1] = {1'b0,layer_2_2[1431:1424]} - {1'b0, layer_1_2[1431:1424]};
      mid_2[2] = {1'b0,layer_2_2[1439:1432]} - {1'b0, layer_1_2[1439:1432]};
      btm_0[0] = {1'b0,layer_3_0[1423:1416]} - {1'b0, layer_2_0[1423:1416]};
      btm_0[1] = {1'b0,layer_3_0[1431:1424]} - {1'b0, layer_2_0[1431:1424]};
      btm_0[2] = {1'b0,layer_3_0[1439:1432]} - {1'b0, layer_2_0[1439:1432]};
      btm_1[0] = {1'b0,layer_3_1[1423:1416]} - {1'b0, layer_2_1[1423:1416]};
      btm_1[1] = {1'b0,layer_3_1[1431:1424]} - {1'b0, layer_2_1[1431:1424]};
      btm_1[2] = {1'b0,layer_3_1[1439:1432]} - {1'b0, layer_2_1[1439:1432]};
      btm_2[0] = {1'b0,layer_3_2[1423:1416]} - {1'b0, layer_2_2[1423:1416]};
      btm_2[1] = {1'b0,layer_3_2[1431:1424]} - {1'b0, layer_2_2[1431:1424]};
      btm_2[2] = {1'b0,layer_3_2[1439:1432]} - {1'b0, layer_2_2[1439:1432]};
    end
    'd179: begin
      top_0[0] = {1'b0,layer_1_0[1431:1424]} - {1'b0, layer_0_0[1431:1424]};
      top_0[1] = {1'b0,layer_1_0[1439:1432]} - {1'b0, layer_0_0[1439:1432]};
      top_0[2] = {1'b0,layer_1_0[1447:1440]} - {1'b0, layer_0_0[1447:1440]};
      top_1[0] = {1'b0,layer_1_1[1431:1424]} - {1'b0, layer_0_1[1431:1424]};
      top_1[1] = {1'b0,layer_1_1[1439:1432]} - {1'b0, layer_0_1[1439:1432]};
      top_1[2] = {1'b0,layer_1_1[1447:1440]} - {1'b0, layer_0_1[1447:1440]};
      top_2[0] = {1'b0,layer_1_2[1431:1424]} - {1'b0, layer_0_2[1431:1424]};
      top_2[1] = {1'b0,layer_1_2[1439:1432]} - {1'b0, layer_0_2[1439:1432]};
      top_2[2] = {1'b0,layer_1_2[1447:1440]} - {1'b0, layer_0_2[1447:1440]};
      mid_0[0] = {1'b0,layer_2_0[1431:1424]} - {1'b0, layer_1_0[1431:1424]};
      mid_0[1] = {1'b0,layer_2_0[1439:1432]} - {1'b0, layer_1_0[1439:1432]};
      mid_0[2] = {1'b0,layer_2_0[1447:1440]} - {1'b0, layer_1_0[1447:1440]};
      mid_1[0] = {1'b0,layer_2_1[1431:1424]} - {1'b0, layer_1_1[1431:1424]};
      mid_1[1] = {1'b0,layer_2_1[1439:1432]} - {1'b0, layer_1_1[1439:1432]};
      mid_1[2] = {1'b0,layer_2_1[1447:1440]} - {1'b0, layer_1_1[1447:1440]};
      mid_2[0] = {1'b0,layer_2_2[1431:1424]} - {1'b0, layer_1_2[1431:1424]};
      mid_2[1] = {1'b0,layer_2_2[1439:1432]} - {1'b0, layer_1_2[1439:1432]};
      mid_2[2] = {1'b0,layer_2_2[1447:1440]} - {1'b0, layer_1_2[1447:1440]};
      btm_0[0] = {1'b0,layer_3_0[1431:1424]} - {1'b0, layer_2_0[1431:1424]};
      btm_0[1] = {1'b0,layer_3_0[1439:1432]} - {1'b0, layer_2_0[1439:1432]};
      btm_0[2] = {1'b0,layer_3_0[1447:1440]} - {1'b0, layer_2_0[1447:1440]};
      btm_1[0] = {1'b0,layer_3_1[1431:1424]} - {1'b0, layer_2_1[1431:1424]};
      btm_1[1] = {1'b0,layer_3_1[1439:1432]} - {1'b0, layer_2_1[1439:1432]};
      btm_1[2] = {1'b0,layer_3_1[1447:1440]} - {1'b0, layer_2_1[1447:1440]};
      btm_2[0] = {1'b0,layer_3_2[1431:1424]} - {1'b0, layer_2_2[1431:1424]};
      btm_2[1] = {1'b0,layer_3_2[1439:1432]} - {1'b0, layer_2_2[1439:1432]};
      btm_2[2] = {1'b0,layer_3_2[1447:1440]} - {1'b0, layer_2_2[1447:1440]};
    end
    'd180: begin
      top_0[0] = {1'b0,layer_1_0[1439:1432]} - {1'b0, layer_0_0[1439:1432]};
      top_0[1] = {1'b0,layer_1_0[1447:1440]} - {1'b0, layer_0_0[1447:1440]};
      top_0[2] = {1'b0,layer_1_0[1455:1448]} - {1'b0, layer_0_0[1455:1448]};
      top_1[0] = {1'b0,layer_1_1[1439:1432]} - {1'b0, layer_0_1[1439:1432]};
      top_1[1] = {1'b0,layer_1_1[1447:1440]} - {1'b0, layer_0_1[1447:1440]};
      top_1[2] = {1'b0,layer_1_1[1455:1448]} - {1'b0, layer_0_1[1455:1448]};
      top_2[0] = {1'b0,layer_1_2[1439:1432]} - {1'b0, layer_0_2[1439:1432]};
      top_2[1] = {1'b0,layer_1_2[1447:1440]} - {1'b0, layer_0_2[1447:1440]};
      top_2[2] = {1'b0,layer_1_2[1455:1448]} - {1'b0, layer_0_2[1455:1448]};
      mid_0[0] = {1'b0,layer_2_0[1439:1432]} - {1'b0, layer_1_0[1439:1432]};
      mid_0[1] = {1'b0,layer_2_0[1447:1440]} - {1'b0, layer_1_0[1447:1440]};
      mid_0[2] = {1'b0,layer_2_0[1455:1448]} - {1'b0, layer_1_0[1455:1448]};
      mid_1[0] = {1'b0,layer_2_1[1439:1432]} - {1'b0, layer_1_1[1439:1432]};
      mid_1[1] = {1'b0,layer_2_1[1447:1440]} - {1'b0, layer_1_1[1447:1440]};
      mid_1[2] = {1'b0,layer_2_1[1455:1448]} - {1'b0, layer_1_1[1455:1448]};
      mid_2[0] = {1'b0,layer_2_2[1439:1432]} - {1'b0, layer_1_2[1439:1432]};
      mid_2[1] = {1'b0,layer_2_2[1447:1440]} - {1'b0, layer_1_2[1447:1440]};
      mid_2[2] = {1'b0,layer_2_2[1455:1448]} - {1'b0, layer_1_2[1455:1448]};
      btm_0[0] = {1'b0,layer_3_0[1439:1432]} - {1'b0, layer_2_0[1439:1432]};
      btm_0[1] = {1'b0,layer_3_0[1447:1440]} - {1'b0, layer_2_0[1447:1440]};
      btm_0[2] = {1'b0,layer_3_0[1455:1448]} - {1'b0, layer_2_0[1455:1448]};
      btm_1[0] = {1'b0,layer_3_1[1439:1432]} - {1'b0, layer_2_1[1439:1432]};
      btm_1[1] = {1'b0,layer_3_1[1447:1440]} - {1'b0, layer_2_1[1447:1440]};
      btm_1[2] = {1'b0,layer_3_1[1455:1448]} - {1'b0, layer_2_1[1455:1448]};
      btm_2[0] = {1'b0,layer_3_2[1439:1432]} - {1'b0, layer_2_2[1439:1432]};
      btm_2[1] = {1'b0,layer_3_2[1447:1440]} - {1'b0, layer_2_2[1447:1440]};
      btm_2[2] = {1'b0,layer_3_2[1455:1448]} - {1'b0, layer_2_2[1455:1448]};
    end
    'd181: begin
      top_0[0] = {1'b0,layer_1_0[1447:1440]} - {1'b0, layer_0_0[1447:1440]};
      top_0[1] = {1'b0,layer_1_0[1455:1448]} - {1'b0, layer_0_0[1455:1448]};
      top_0[2] = {1'b0,layer_1_0[1463:1456]} - {1'b0, layer_0_0[1463:1456]};
      top_1[0] = {1'b0,layer_1_1[1447:1440]} - {1'b0, layer_0_1[1447:1440]};
      top_1[1] = {1'b0,layer_1_1[1455:1448]} - {1'b0, layer_0_1[1455:1448]};
      top_1[2] = {1'b0,layer_1_1[1463:1456]} - {1'b0, layer_0_1[1463:1456]};
      top_2[0] = {1'b0,layer_1_2[1447:1440]} - {1'b0, layer_0_2[1447:1440]};
      top_2[1] = {1'b0,layer_1_2[1455:1448]} - {1'b0, layer_0_2[1455:1448]};
      top_2[2] = {1'b0,layer_1_2[1463:1456]} - {1'b0, layer_0_2[1463:1456]};
      mid_0[0] = {1'b0,layer_2_0[1447:1440]} - {1'b0, layer_1_0[1447:1440]};
      mid_0[1] = {1'b0,layer_2_0[1455:1448]} - {1'b0, layer_1_0[1455:1448]};
      mid_0[2] = {1'b0,layer_2_0[1463:1456]} - {1'b0, layer_1_0[1463:1456]};
      mid_1[0] = {1'b0,layer_2_1[1447:1440]} - {1'b0, layer_1_1[1447:1440]};
      mid_1[1] = {1'b0,layer_2_1[1455:1448]} - {1'b0, layer_1_1[1455:1448]};
      mid_1[2] = {1'b0,layer_2_1[1463:1456]} - {1'b0, layer_1_1[1463:1456]};
      mid_2[0] = {1'b0,layer_2_2[1447:1440]} - {1'b0, layer_1_2[1447:1440]};
      mid_2[1] = {1'b0,layer_2_2[1455:1448]} - {1'b0, layer_1_2[1455:1448]};
      mid_2[2] = {1'b0,layer_2_2[1463:1456]} - {1'b0, layer_1_2[1463:1456]};
      btm_0[0] = {1'b0,layer_3_0[1447:1440]} - {1'b0, layer_2_0[1447:1440]};
      btm_0[1] = {1'b0,layer_3_0[1455:1448]} - {1'b0, layer_2_0[1455:1448]};
      btm_0[2] = {1'b0,layer_3_0[1463:1456]} - {1'b0, layer_2_0[1463:1456]};
      btm_1[0] = {1'b0,layer_3_1[1447:1440]} - {1'b0, layer_2_1[1447:1440]};
      btm_1[1] = {1'b0,layer_3_1[1455:1448]} - {1'b0, layer_2_1[1455:1448]};
      btm_1[2] = {1'b0,layer_3_1[1463:1456]} - {1'b0, layer_2_1[1463:1456]};
      btm_2[0] = {1'b0,layer_3_2[1447:1440]} - {1'b0, layer_2_2[1447:1440]};
      btm_2[1] = {1'b0,layer_3_2[1455:1448]} - {1'b0, layer_2_2[1455:1448]};
      btm_2[2] = {1'b0,layer_3_2[1463:1456]} - {1'b0, layer_2_2[1463:1456]};
    end
    'd182: begin
      top_0[0] = {1'b0,layer_1_0[1455:1448]} - {1'b0, layer_0_0[1455:1448]};
      top_0[1] = {1'b0,layer_1_0[1463:1456]} - {1'b0, layer_0_0[1463:1456]};
      top_0[2] = {1'b0,layer_1_0[1471:1464]} - {1'b0, layer_0_0[1471:1464]};
      top_1[0] = {1'b0,layer_1_1[1455:1448]} - {1'b0, layer_0_1[1455:1448]};
      top_1[1] = {1'b0,layer_1_1[1463:1456]} - {1'b0, layer_0_1[1463:1456]};
      top_1[2] = {1'b0,layer_1_1[1471:1464]} - {1'b0, layer_0_1[1471:1464]};
      top_2[0] = {1'b0,layer_1_2[1455:1448]} - {1'b0, layer_0_2[1455:1448]};
      top_2[1] = {1'b0,layer_1_2[1463:1456]} - {1'b0, layer_0_2[1463:1456]};
      top_2[2] = {1'b0,layer_1_2[1471:1464]} - {1'b0, layer_0_2[1471:1464]};
      mid_0[0] = {1'b0,layer_2_0[1455:1448]} - {1'b0, layer_1_0[1455:1448]};
      mid_0[1] = {1'b0,layer_2_0[1463:1456]} - {1'b0, layer_1_0[1463:1456]};
      mid_0[2] = {1'b0,layer_2_0[1471:1464]} - {1'b0, layer_1_0[1471:1464]};
      mid_1[0] = {1'b0,layer_2_1[1455:1448]} - {1'b0, layer_1_1[1455:1448]};
      mid_1[1] = {1'b0,layer_2_1[1463:1456]} - {1'b0, layer_1_1[1463:1456]};
      mid_1[2] = {1'b0,layer_2_1[1471:1464]} - {1'b0, layer_1_1[1471:1464]};
      mid_2[0] = {1'b0,layer_2_2[1455:1448]} - {1'b0, layer_1_2[1455:1448]};
      mid_2[1] = {1'b0,layer_2_2[1463:1456]} - {1'b0, layer_1_2[1463:1456]};
      mid_2[2] = {1'b0,layer_2_2[1471:1464]} - {1'b0, layer_1_2[1471:1464]};
      btm_0[0] = {1'b0,layer_3_0[1455:1448]} - {1'b0, layer_2_0[1455:1448]};
      btm_0[1] = {1'b0,layer_3_0[1463:1456]} - {1'b0, layer_2_0[1463:1456]};
      btm_0[2] = {1'b0,layer_3_0[1471:1464]} - {1'b0, layer_2_0[1471:1464]};
      btm_1[0] = {1'b0,layer_3_1[1455:1448]} - {1'b0, layer_2_1[1455:1448]};
      btm_1[1] = {1'b0,layer_3_1[1463:1456]} - {1'b0, layer_2_1[1463:1456]};
      btm_1[2] = {1'b0,layer_3_1[1471:1464]} - {1'b0, layer_2_1[1471:1464]};
      btm_2[0] = {1'b0,layer_3_2[1455:1448]} - {1'b0, layer_2_2[1455:1448]};
      btm_2[1] = {1'b0,layer_3_2[1463:1456]} - {1'b0, layer_2_2[1463:1456]};
      btm_2[2] = {1'b0,layer_3_2[1471:1464]} - {1'b0, layer_2_2[1471:1464]};
    end
    'd183: begin
      top_0[0] = {1'b0,layer_1_0[1463:1456]} - {1'b0, layer_0_0[1463:1456]};
      top_0[1] = {1'b0,layer_1_0[1471:1464]} - {1'b0, layer_0_0[1471:1464]};
      top_0[2] = {1'b0,layer_1_0[1479:1472]} - {1'b0, layer_0_0[1479:1472]};
      top_1[0] = {1'b0,layer_1_1[1463:1456]} - {1'b0, layer_0_1[1463:1456]};
      top_1[1] = {1'b0,layer_1_1[1471:1464]} - {1'b0, layer_0_1[1471:1464]};
      top_1[2] = {1'b0,layer_1_1[1479:1472]} - {1'b0, layer_0_1[1479:1472]};
      top_2[0] = {1'b0,layer_1_2[1463:1456]} - {1'b0, layer_0_2[1463:1456]};
      top_2[1] = {1'b0,layer_1_2[1471:1464]} - {1'b0, layer_0_2[1471:1464]};
      top_2[2] = {1'b0,layer_1_2[1479:1472]} - {1'b0, layer_0_2[1479:1472]};
      mid_0[0] = {1'b0,layer_2_0[1463:1456]} - {1'b0, layer_1_0[1463:1456]};
      mid_0[1] = {1'b0,layer_2_0[1471:1464]} - {1'b0, layer_1_0[1471:1464]};
      mid_0[2] = {1'b0,layer_2_0[1479:1472]} - {1'b0, layer_1_0[1479:1472]};
      mid_1[0] = {1'b0,layer_2_1[1463:1456]} - {1'b0, layer_1_1[1463:1456]};
      mid_1[1] = {1'b0,layer_2_1[1471:1464]} - {1'b0, layer_1_1[1471:1464]};
      mid_1[2] = {1'b0,layer_2_1[1479:1472]} - {1'b0, layer_1_1[1479:1472]};
      mid_2[0] = {1'b0,layer_2_2[1463:1456]} - {1'b0, layer_1_2[1463:1456]};
      mid_2[1] = {1'b0,layer_2_2[1471:1464]} - {1'b0, layer_1_2[1471:1464]};
      mid_2[2] = {1'b0,layer_2_2[1479:1472]} - {1'b0, layer_1_2[1479:1472]};
      btm_0[0] = {1'b0,layer_3_0[1463:1456]} - {1'b0, layer_2_0[1463:1456]};
      btm_0[1] = {1'b0,layer_3_0[1471:1464]} - {1'b0, layer_2_0[1471:1464]};
      btm_0[2] = {1'b0,layer_3_0[1479:1472]} - {1'b0, layer_2_0[1479:1472]};
      btm_1[0] = {1'b0,layer_3_1[1463:1456]} - {1'b0, layer_2_1[1463:1456]};
      btm_1[1] = {1'b0,layer_3_1[1471:1464]} - {1'b0, layer_2_1[1471:1464]};
      btm_1[2] = {1'b0,layer_3_1[1479:1472]} - {1'b0, layer_2_1[1479:1472]};
      btm_2[0] = {1'b0,layer_3_2[1463:1456]} - {1'b0, layer_2_2[1463:1456]};
      btm_2[1] = {1'b0,layer_3_2[1471:1464]} - {1'b0, layer_2_2[1471:1464]};
      btm_2[2] = {1'b0,layer_3_2[1479:1472]} - {1'b0, layer_2_2[1479:1472]};
    end
    'd184: begin
      top_0[0] = {1'b0,layer_1_0[1471:1464]} - {1'b0, layer_0_0[1471:1464]};
      top_0[1] = {1'b0,layer_1_0[1479:1472]} - {1'b0, layer_0_0[1479:1472]};
      top_0[2] = {1'b0,layer_1_0[1487:1480]} - {1'b0, layer_0_0[1487:1480]};
      top_1[0] = {1'b0,layer_1_1[1471:1464]} - {1'b0, layer_0_1[1471:1464]};
      top_1[1] = {1'b0,layer_1_1[1479:1472]} - {1'b0, layer_0_1[1479:1472]};
      top_1[2] = {1'b0,layer_1_1[1487:1480]} - {1'b0, layer_0_1[1487:1480]};
      top_2[0] = {1'b0,layer_1_2[1471:1464]} - {1'b0, layer_0_2[1471:1464]};
      top_2[1] = {1'b0,layer_1_2[1479:1472]} - {1'b0, layer_0_2[1479:1472]};
      top_2[2] = {1'b0,layer_1_2[1487:1480]} - {1'b0, layer_0_2[1487:1480]};
      mid_0[0] = {1'b0,layer_2_0[1471:1464]} - {1'b0, layer_1_0[1471:1464]};
      mid_0[1] = {1'b0,layer_2_0[1479:1472]} - {1'b0, layer_1_0[1479:1472]};
      mid_0[2] = {1'b0,layer_2_0[1487:1480]} - {1'b0, layer_1_0[1487:1480]};
      mid_1[0] = {1'b0,layer_2_1[1471:1464]} - {1'b0, layer_1_1[1471:1464]};
      mid_1[1] = {1'b0,layer_2_1[1479:1472]} - {1'b0, layer_1_1[1479:1472]};
      mid_1[2] = {1'b0,layer_2_1[1487:1480]} - {1'b0, layer_1_1[1487:1480]};
      mid_2[0] = {1'b0,layer_2_2[1471:1464]} - {1'b0, layer_1_2[1471:1464]};
      mid_2[1] = {1'b0,layer_2_2[1479:1472]} - {1'b0, layer_1_2[1479:1472]};
      mid_2[2] = {1'b0,layer_2_2[1487:1480]} - {1'b0, layer_1_2[1487:1480]};
      btm_0[0] = {1'b0,layer_3_0[1471:1464]} - {1'b0, layer_2_0[1471:1464]};
      btm_0[1] = {1'b0,layer_3_0[1479:1472]} - {1'b0, layer_2_0[1479:1472]};
      btm_0[2] = {1'b0,layer_3_0[1487:1480]} - {1'b0, layer_2_0[1487:1480]};
      btm_1[0] = {1'b0,layer_3_1[1471:1464]} - {1'b0, layer_2_1[1471:1464]};
      btm_1[1] = {1'b0,layer_3_1[1479:1472]} - {1'b0, layer_2_1[1479:1472]};
      btm_1[2] = {1'b0,layer_3_1[1487:1480]} - {1'b0, layer_2_1[1487:1480]};
      btm_2[0] = {1'b0,layer_3_2[1471:1464]} - {1'b0, layer_2_2[1471:1464]};
      btm_2[1] = {1'b0,layer_3_2[1479:1472]} - {1'b0, layer_2_2[1479:1472]};
      btm_2[2] = {1'b0,layer_3_2[1487:1480]} - {1'b0, layer_2_2[1487:1480]};
    end
    'd185: begin
      top_0[0] = {1'b0,layer_1_0[1479:1472]} - {1'b0, layer_0_0[1479:1472]};
      top_0[1] = {1'b0,layer_1_0[1487:1480]} - {1'b0, layer_0_0[1487:1480]};
      top_0[2] = {1'b0,layer_1_0[1495:1488]} - {1'b0, layer_0_0[1495:1488]};
      top_1[0] = {1'b0,layer_1_1[1479:1472]} - {1'b0, layer_0_1[1479:1472]};
      top_1[1] = {1'b0,layer_1_1[1487:1480]} - {1'b0, layer_0_1[1487:1480]};
      top_1[2] = {1'b0,layer_1_1[1495:1488]} - {1'b0, layer_0_1[1495:1488]};
      top_2[0] = {1'b0,layer_1_2[1479:1472]} - {1'b0, layer_0_2[1479:1472]};
      top_2[1] = {1'b0,layer_1_2[1487:1480]} - {1'b0, layer_0_2[1487:1480]};
      top_2[2] = {1'b0,layer_1_2[1495:1488]} - {1'b0, layer_0_2[1495:1488]};
      mid_0[0] = {1'b0,layer_2_0[1479:1472]} - {1'b0, layer_1_0[1479:1472]};
      mid_0[1] = {1'b0,layer_2_0[1487:1480]} - {1'b0, layer_1_0[1487:1480]};
      mid_0[2] = {1'b0,layer_2_0[1495:1488]} - {1'b0, layer_1_0[1495:1488]};
      mid_1[0] = {1'b0,layer_2_1[1479:1472]} - {1'b0, layer_1_1[1479:1472]};
      mid_1[1] = {1'b0,layer_2_1[1487:1480]} - {1'b0, layer_1_1[1487:1480]};
      mid_1[2] = {1'b0,layer_2_1[1495:1488]} - {1'b0, layer_1_1[1495:1488]};
      mid_2[0] = {1'b0,layer_2_2[1479:1472]} - {1'b0, layer_1_2[1479:1472]};
      mid_2[1] = {1'b0,layer_2_2[1487:1480]} - {1'b0, layer_1_2[1487:1480]};
      mid_2[2] = {1'b0,layer_2_2[1495:1488]} - {1'b0, layer_1_2[1495:1488]};
      btm_0[0] = {1'b0,layer_3_0[1479:1472]} - {1'b0, layer_2_0[1479:1472]};
      btm_0[1] = {1'b0,layer_3_0[1487:1480]} - {1'b0, layer_2_0[1487:1480]};
      btm_0[2] = {1'b0,layer_3_0[1495:1488]} - {1'b0, layer_2_0[1495:1488]};
      btm_1[0] = {1'b0,layer_3_1[1479:1472]} - {1'b0, layer_2_1[1479:1472]};
      btm_1[1] = {1'b0,layer_3_1[1487:1480]} - {1'b0, layer_2_1[1487:1480]};
      btm_1[2] = {1'b0,layer_3_1[1495:1488]} - {1'b0, layer_2_1[1495:1488]};
      btm_2[0] = {1'b0,layer_3_2[1479:1472]} - {1'b0, layer_2_2[1479:1472]};
      btm_2[1] = {1'b0,layer_3_2[1487:1480]} - {1'b0, layer_2_2[1487:1480]};
      btm_2[2] = {1'b0,layer_3_2[1495:1488]} - {1'b0, layer_2_2[1495:1488]};
    end
    'd186: begin
      top_0[0] = {1'b0,layer_1_0[1487:1480]} - {1'b0, layer_0_0[1487:1480]};
      top_0[1] = {1'b0,layer_1_0[1495:1488]} - {1'b0, layer_0_0[1495:1488]};
      top_0[2] = {1'b0,layer_1_0[1503:1496]} - {1'b0, layer_0_0[1503:1496]};
      top_1[0] = {1'b0,layer_1_1[1487:1480]} - {1'b0, layer_0_1[1487:1480]};
      top_1[1] = {1'b0,layer_1_1[1495:1488]} - {1'b0, layer_0_1[1495:1488]};
      top_1[2] = {1'b0,layer_1_1[1503:1496]} - {1'b0, layer_0_1[1503:1496]};
      top_2[0] = {1'b0,layer_1_2[1487:1480]} - {1'b0, layer_0_2[1487:1480]};
      top_2[1] = {1'b0,layer_1_2[1495:1488]} - {1'b0, layer_0_2[1495:1488]};
      top_2[2] = {1'b0,layer_1_2[1503:1496]} - {1'b0, layer_0_2[1503:1496]};
      mid_0[0] = {1'b0,layer_2_0[1487:1480]} - {1'b0, layer_1_0[1487:1480]};
      mid_0[1] = {1'b0,layer_2_0[1495:1488]} - {1'b0, layer_1_0[1495:1488]};
      mid_0[2] = {1'b0,layer_2_0[1503:1496]} - {1'b0, layer_1_0[1503:1496]};
      mid_1[0] = {1'b0,layer_2_1[1487:1480]} - {1'b0, layer_1_1[1487:1480]};
      mid_1[1] = {1'b0,layer_2_1[1495:1488]} - {1'b0, layer_1_1[1495:1488]};
      mid_1[2] = {1'b0,layer_2_1[1503:1496]} - {1'b0, layer_1_1[1503:1496]};
      mid_2[0] = {1'b0,layer_2_2[1487:1480]} - {1'b0, layer_1_2[1487:1480]};
      mid_2[1] = {1'b0,layer_2_2[1495:1488]} - {1'b0, layer_1_2[1495:1488]};
      mid_2[2] = {1'b0,layer_2_2[1503:1496]} - {1'b0, layer_1_2[1503:1496]};
      btm_0[0] = {1'b0,layer_3_0[1487:1480]} - {1'b0, layer_2_0[1487:1480]};
      btm_0[1] = {1'b0,layer_3_0[1495:1488]} - {1'b0, layer_2_0[1495:1488]};
      btm_0[2] = {1'b0,layer_3_0[1503:1496]} - {1'b0, layer_2_0[1503:1496]};
      btm_1[0] = {1'b0,layer_3_1[1487:1480]} - {1'b0, layer_2_1[1487:1480]};
      btm_1[1] = {1'b0,layer_3_1[1495:1488]} - {1'b0, layer_2_1[1495:1488]};
      btm_1[2] = {1'b0,layer_3_1[1503:1496]} - {1'b0, layer_2_1[1503:1496]};
      btm_2[0] = {1'b0,layer_3_2[1487:1480]} - {1'b0, layer_2_2[1487:1480]};
      btm_2[1] = {1'b0,layer_3_2[1495:1488]} - {1'b0, layer_2_2[1495:1488]};
      btm_2[2] = {1'b0,layer_3_2[1503:1496]} - {1'b0, layer_2_2[1503:1496]};
    end
    'd187: begin
      top_0[0] = {1'b0,layer_1_0[1495:1488]} - {1'b0, layer_0_0[1495:1488]};
      top_0[1] = {1'b0,layer_1_0[1503:1496]} - {1'b0, layer_0_0[1503:1496]};
      top_0[2] = {1'b0,layer_1_0[1511:1504]} - {1'b0, layer_0_0[1511:1504]};
      top_1[0] = {1'b0,layer_1_1[1495:1488]} - {1'b0, layer_0_1[1495:1488]};
      top_1[1] = {1'b0,layer_1_1[1503:1496]} - {1'b0, layer_0_1[1503:1496]};
      top_1[2] = {1'b0,layer_1_1[1511:1504]} - {1'b0, layer_0_1[1511:1504]};
      top_2[0] = {1'b0,layer_1_2[1495:1488]} - {1'b0, layer_0_2[1495:1488]};
      top_2[1] = {1'b0,layer_1_2[1503:1496]} - {1'b0, layer_0_2[1503:1496]};
      top_2[2] = {1'b0,layer_1_2[1511:1504]} - {1'b0, layer_0_2[1511:1504]};
      mid_0[0] = {1'b0,layer_2_0[1495:1488]} - {1'b0, layer_1_0[1495:1488]};
      mid_0[1] = {1'b0,layer_2_0[1503:1496]} - {1'b0, layer_1_0[1503:1496]};
      mid_0[2] = {1'b0,layer_2_0[1511:1504]} - {1'b0, layer_1_0[1511:1504]};
      mid_1[0] = {1'b0,layer_2_1[1495:1488]} - {1'b0, layer_1_1[1495:1488]};
      mid_1[1] = {1'b0,layer_2_1[1503:1496]} - {1'b0, layer_1_1[1503:1496]};
      mid_1[2] = {1'b0,layer_2_1[1511:1504]} - {1'b0, layer_1_1[1511:1504]};
      mid_2[0] = {1'b0,layer_2_2[1495:1488]} - {1'b0, layer_1_2[1495:1488]};
      mid_2[1] = {1'b0,layer_2_2[1503:1496]} - {1'b0, layer_1_2[1503:1496]};
      mid_2[2] = {1'b0,layer_2_2[1511:1504]} - {1'b0, layer_1_2[1511:1504]};
      btm_0[0] = {1'b0,layer_3_0[1495:1488]} - {1'b0, layer_2_0[1495:1488]};
      btm_0[1] = {1'b0,layer_3_0[1503:1496]} - {1'b0, layer_2_0[1503:1496]};
      btm_0[2] = {1'b0,layer_3_0[1511:1504]} - {1'b0, layer_2_0[1511:1504]};
      btm_1[0] = {1'b0,layer_3_1[1495:1488]} - {1'b0, layer_2_1[1495:1488]};
      btm_1[1] = {1'b0,layer_3_1[1503:1496]} - {1'b0, layer_2_1[1503:1496]};
      btm_1[2] = {1'b0,layer_3_1[1511:1504]} - {1'b0, layer_2_1[1511:1504]};
      btm_2[0] = {1'b0,layer_3_2[1495:1488]} - {1'b0, layer_2_2[1495:1488]};
      btm_2[1] = {1'b0,layer_3_2[1503:1496]} - {1'b0, layer_2_2[1503:1496]};
      btm_2[2] = {1'b0,layer_3_2[1511:1504]} - {1'b0, layer_2_2[1511:1504]};
    end
    'd188: begin
      top_0[0] = {1'b0,layer_1_0[1503:1496]} - {1'b0, layer_0_0[1503:1496]};
      top_0[1] = {1'b0,layer_1_0[1511:1504]} - {1'b0, layer_0_0[1511:1504]};
      top_0[2] = {1'b0,layer_1_0[1519:1512]} - {1'b0, layer_0_0[1519:1512]};
      top_1[0] = {1'b0,layer_1_1[1503:1496]} - {1'b0, layer_0_1[1503:1496]};
      top_1[1] = {1'b0,layer_1_1[1511:1504]} - {1'b0, layer_0_1[1511:1504]};
      top_1[2] = {1'b0,layer_1_1[1519:1512]} - {1'b0, layer_0_1[1519:1512]};
      top_2[0] = {1'b0,layer_1_2[1503:1496]} - {1'b0, layer_0_2[1503:1496]};
      top_2[1] = {1'b0,layer_1_2[1511:1504]} - {1'b0, layer_0_2[1511:1504]};
      top_2[2] = {1'b0,layer_1_2[1519:1512]} - {1'b0, layer_0_2[1519:1512]};
      mid_0[0] = {1'b0,layer_2_0[1503:1496]} - {1'b0, layer_1_0[1503:1496]};
      mid_0[1] = {1'b0,layer_2_0[1511:1504]} - {1'b0, layer_1_0[1511:1504]};
      mid_0[2] = {1'b0,layer_2_0[1519:1512]} - {1'b0, layer_1_0[1519:1512]};
      mid_1[0] = {1'b0,layer_2_1[1503:1496]} - {1'b0, layer_1_1[1503:1496]};
      mid_1[1] = {1'b0,layer_2_1[1511:1504]} - {1'b0, layer_1_1[1511:1504]};
      mid_1[2] = {1'b0,layer_2_1[1519:1512]} - {1'b0, layer_1_1[1519:1512]};
      mid_2[0] = {1'b0,layer_2_2[1503:1496]} - {1'b0, layer_1_2[1503:1496]};
      mid_2[1] = {1'b0,layer_2_2[1511:1504]} - {1'b0, layer_1_2[1511:1504]};
      mid_2[2] = {1'b0,layer_2_2[1519:1512]} - {1'b0, layer_1_2[1519:1512]};
      btm_0[0] = {1'b0,layer_3_0[1503:1496]} - {1'b0, layer_2_0[1503:1496]};
      btm_0[1] = {1'b0,layer_3_0[1511:1504]} - {1'b0, layer_2_0[1511:1504]};
      btm_0[2] = {1'b0,layer_3_0[1519:1512]} - {1'b0, layer_2_0[1519:1512]};
      btm_1[0] = {1'b0,layer_3_1[1503:1496]} - {1'b0, layer_2_1[1503:1496]};
      btm_1[1] = {1'b0,layer_3_1[1511:1504]} - {1'b0, layer_2_1[1511:1504]};
      btm_1[2] = {1'b0,layer_3_1[1519:1512]} - {1'b0, layer_2_1[1519:1512]};
      btm_2[0] = {1'b0,layer_3_2[1503:1496]} - {1'b0, layer_2_2[1503:1496]};
      btm_2[1] = {1'b0,layer_3_2[1511:1504]} - {1'b0, layer_2_2[1511:1504]};
      btm_2[2] = {1'b0,layer_3_2[1519:1512]} - {1'b0, layer_2_2[1519:1512]};
    end
    'd189: begin
      top_0[0] = {1'b0,layer_1_0[1511:1504]} - {1'b0, layer_0_0[1511:1504]};
      top_0[1] = {1'b0,layer_1_0[1519:1512]} - {1'b0, layer_0_0[1519:1512]};
      top_0[2] = {1'b0,layer_1_0[1527:1520]} - {1'b0, layer_0_0[1527:1520]};
      top_1[0] = {1'b0,layer_1_1[1511:1504]} - {1'b0, layer_0_1[1511:1504]};
      top_1[1] = {1'b0,layer_1_1[1519:1512]} - {1'b0, layer_0_1[1519:1512]};
      top_1[2] = {1'b0,layer_1_1[1527:1520]} - {1'b0, layer_0_1[1527:1520]};
      top_2[0] = {1'b0,layer_1_2[1511:1504]} - {1'b0, layer_0_2[1511:1504]};
      top_2[1] = {1'b0,layer_1_2[1519:1512]} - {1'b0, layer_0_2[1519:1512]};
      top_2[2] = {1'b0,layer_1_2[1527:1520]} - {1'b0, layer_0_2[1527:1520]};
      mid_0[0] = {1'b0,layer_2_0[1511:1504]} - {1'b0, layer_1_0[1511:1504]};
      mid_0[1] = {1'b0,layer_2_0[1519:1512]} - {1'b0, layer_1_0[1519:1512]};
      mid_0[2] = {1'b0,layer_2_0[1527:1520]} - {1'b0, layer_1_0[1527:1520]};
      mid_1[0] = {1'b0,layer_2_1[1511:1504]} - {1'b0, layer_1_1[1511:1504]};
      mid_1[1] = {1'b0,layer_2_1[1519:1512]} - {1'b0, layer_1_1[1519:1512]};
      mid_1[2] = {1'b0,layer_2_1[1527:1520]} - {1'b0, layer_1_1[1527:1520]};
      mid_2[0] = {1'b0,layer_2_2[1511:1504]} - {1'b0, layer_1_2[1511:1504]};
      mid_2[1] = {1'b0,layer_2_2[1519:1512]} - {1'b0, layer_1_2[1519:1512]};
      mid_2[2] = {1'b0,layer_2_2[1527:1520]} - {1'b0, layer_1_2[1527:1520]};
      btm_0[0] = {1'b0,layer_3_0[1511:1504]} - {1'b0, layer_2_0[1511:1504]};
      btm_0[1] = {1'b0,layer_3_0[1519:1512]} - {1'b0, layer_2_0[1519:1512]};
      btm_0[2] = {1'b0,layer_3_0[1527:1520]} - {1'b0, layer_2_0[1527:1520]};
      btm_1[0] = {1'b0,layer_3_1[1511:1504]} - {1'b0, layer_2_1[1511:1504]};
      btm_1[1] = {1'b0,layer_3_1[1519:1512]} - {1'b0, layer_2_1[1519:1512]};
      btm_1[2] = {1'b0,layer_3_1[1527:1520]} - {1'b0, layer_2_1[1527:1520]};
      btm_2[0] = {1'b0,layer_3_2[1511:1504]} - {1'b0, layer_2_2[1511:1504]};
      btm_2[1] = {1'b0,layer_3_2[1519:1512]} - {1'b0, layer_2_2[1519:1512]};
      btm_2[2] = {1'b0,layer_3_2[1527:1520]} - {1'b0, layer_2_2[1527:1520]};
    end
    'd190: begin
      top_0[0] = {1'b0,layer_1_0[1519:1512]} - {1'b0, layer_0_0[1519:1512]};
      top_0[1] = {1'b0,layer_1_0[1527:1520]} - {1'b0, layer_0_0[1527:1520]};
      top_0[2] = {1'b0,layer_1_0[1535:1528]} - {1'b0, layer_0_0[1535:1528]};
      top_1[0] = {1'b0,layer_1_1[1519:1512]} - {1'b0, layer_0_1[1519:1512]};
      top_1[1] = {1'b0,layer_1_1[1527:1520]} - {1'b0, layer_0_1[1527:1520]};
      top_1[2] = {1'b0,layer_1_1[1535:1528]} - {1'b0, layer_0_1[1535:1528]};
      top_2[0] = {1'b0,layer_1_2[1519:1512]} - {1'b0, layer_0_2[1519:1512]};
      top_2[1] = {1'b0,layer_1_2[1527:1520]} - {1'b0, layer_0_2[1527:1520]};
      top_2[2] = {1'b0,layer_1_2[1535:1528]} - {1'b0, layer_0_2[1535:1528]};
      mid_0[0] = {1'b0,layer_2_0[1519:1512]} - {1'b0, layer_1_0[1519:1512]};
      mid_0[1] = {1'b0,layer_2_0[1527:1520]} - {1'b0, layer_1_0[1527:1520]};
      mid_0[2] = {1'b0,layer_2_0[1535:1528]} - {1'b0, layer_1_0[1535:1528]};
      mid_1[0] = {1'b0,layer_2_1[1519:1512]} - {1'b0, layer_1_1[1519:1512]};
      mid_1[1] = {1'b0,layer_2_1[1527:1520]} - {1'b0, layer_1_1[1527:1520]};
      mid_1[2] = {1'b0,layer_2_1[1535:1528]} - {1'b0, layer_1_1[1535:1528]};
      mid_2[0] = {1'b0,layer_2_2[1519:1512]} - {1'b0, layer_1_2[1519:1512]};
      mid_2[1] = {1'b0,layer_2_2[1527:1520]} - {1'b0, layer_1_2[1527:1520]};
      mid_2[2] = {1'b0,layer_2_2[1535:1528]} - {1'b0, layer_1_2[1535:1528]};
      btm_0[0] = {1'b0,layer_3_0[1519:1512]} - {1'b0, layer_2_0[1519:1512]};
      btm_0[1] = {1'b0,layer_3_0[1527:1520]} - {1'b0, layer_2_0[1527:1520]};
      btm_0[2] = {1'b0,layer_3_0[1535:1528]} - {1'b0, layer_2_0[1535:1528]};
      btm_1[0] = {1'b0,layer_3_1[1519:1512]} - {1'b0, layer_2_1[1519:1512]};
      btm_1[1] = {1'b0,layer_3_1[1527:1520]} - {1'b0, layer_2_1[1527:1520]};
      btm_1[2] = {1'b0,layer_3_1[1535:1528]} - {1'b0, layer_2_1[1535:1528]};
      btm_2[0] = {1'b0,layer_3_2[1519:1512]} - {1'b0, layer_2_2[1519:1512]};
      btm_2[1] = {1'b0,layer_3_2[1527:1520]} - {1'b0, layer_2_2[1527:1520]};
      btm_2[2] = {1'b0,layer_3_2[1535:1528]} - {1'b0, layer_2_2[1535:1528]};
    end
    'd191: begin
      top_0[0] = {1'b0,layer_1_0[1527:1520]} - {1'b0, layer_0_0[1527:1520]};
      top_0[1] = {1'b0,layer_1_0[1535:1528]} - {1'b0, layer_0_0[1535:1528]};
      top_0[2] = {1'b0,layer_1_0[1543:1536]} - {1'b0, layer_0_0[1543:1536]};
      top_1[0] = {1'b0,layer_1_1[1527:1520]} - {1'b0, layer_0_1[1527:1520]};
      top_1[1] = {1'b0,layer_1_1[1535:1528]} - {1'b0, layer_0_1[1535:1528]};
      top_1[2] = {1'b0,layer_1_1[1543:1536]} - {1'b0, layer_0_1[1543:1536]};
      top_2[0] = {1'b0,layer_1_2[1527:1520]} - {1'b0, layer_0_2[1527:1520]};
      top_2[1] = {1'b0,layer_1_2[1535:1528]} - {1'b0, layer_0_2[1535:1528]};
      top_2[2] = {1'b0,layer_1_2[1543:1536]} - {1'b0, layer_0_2[1543:1536]};
      mid_0[0] = {1'b0,layer_2_0[1527:1520]} - {1'b0, layer_1_0[1527:1520]};
      mid_0[1] = {1'b0,layer_2_0[1535:1528]} - {1'b0, layer_1_0[1535:1528]};
      mid_0[2] = {1'b0,layer_2_0[1543:1536]} - {1'b0, layer_1_0[1543:1536]};
      mid_1[0] = {1'b0,layer_2_1[1527:1520]} - {1'b0, layer_1_1[1527:1520]};
      mid_1[1] = {1'b0,layer_2_1[1535:1528]} - {1'b0, layer_1_1[1535:1528]};
      mid_1[2] = {1'b0,layer_2_1[1543:1536]} - {1'b0, layer_1_1[1543:1536]};
      mid_2[0] = {1'b0,layer_2_2[1527:1520]} - {1'b0, layer_1_2[1527:1520]};
      mid_2[1] = {1'b0,layer_2_2[1535:1528]} - {1'b0, layer_1_2[1535:1528]};
      mid_2[2] = {1'b0,layer_2_2[1543:1536]} - {1'b0, layer_1_2[1543:1536]};
      btm_0[0] = {1'b0,layer_3_0[1527:1520]} - {1'b0, layer_2_0[1527:1520]};
      btm_0[1] = {1'b0,layer_3_0[1535:1528]} - {1'b0, layer_2_0[1535:1528]};
      btm_0[2] = {1'b0,layer_3_0[1543:1536]} - {1'b0, layer_2_0[1543:1536]};
      btm_1[0] = {1'b0,layer_3_1[1527:1520]} - {1'b0, layer_2_1[1527:1520]};
      btm_1[1] = {1'b0,layer_3_1[1535:1528]} - {1'b0, layer_2_1[1535:1528]};
      btm_1[2] = {1'b0,layer_3_1[1543:1536]} - {1'b0, layer_2_1[1543:1536]};
      btm_2[0] = {1'b0,layer_3_2[1527:1520]} - {1'b0, layer_2_2[1527:1520]};
      btm_2[1] = {1'b0,layer_3_2[1535:1528]} - {1'b0, layer_2_2[1535:1528]};
      btm_2[2] = {1'b0,layer_3_2[1543:1536]} - {1'b0, layer_2_2[1543:1536]};
    end
    'd192: begin
      top_0[0] = {1'b0,layer_1_0[1535:1528]} - {1'b0, layer_0_0[1535:1528]};
      top_0[1] = {1'b0,layer_1_0[1543:1536]} - {1'b0, layer_0_0[1543:1536]};
      top_0[2] = {1'b0,layer_1_0[1551:1544]} - {1'b0, layer_0_0[1551:1544]};
      top_1[0] = {1'b0,layer_1_1[1535:1528]} - {1'b0, layer_0_1[1535:1528]};
      top_1[1] = {1'b0,layer_1_1[1543:1536]} - {1'b0, layer_0_1[1543:1536]};
      top_1[2] = {1'b0,layer_1_1[1551:1544]} - {1'b0, layer_0_1[1551:1544]};
      top_2[0] = {1'b0,layer_1_2[1535:1528]} - {1'b0, layer_0_2[1535:1528]};
      top_2[1] = {1'b0,layer_1_2[1543:1536]} - {1'b0, layer_0_2[1543:1536]};
      top_2[2] = {1'b0,layer_1_2[1551:1544]} - {1'b0, layer_0_2[1551:1544]};
      mid_0[0] = {1'b0,layer_2_0[1535:1528]} - {1'b0, layer_1_0[1535:1528]};
      mid_0[1] = {1'b0,layer_2_0[1543:1536]} - {1'b0, layer_1_0[1543:1536]};
      mid_0[2] = {1'b0,layer_2_0[1551:1544]} - {1'b0, layer_1_0[1551:1544]};
      mid_1[0] = {1'b0,layer_2_1[1535:1528]} - {1'b0, layer_1_1[1535:1528]};
      mid_1[1] = {1'b0,layer_2_1[1543:1536]} - {1'b0, layer_1_1[1543:1536]};
      mid_1[2] = {1'b0,layer_2_1[1551:1544]} - {1'b0, layer_1_1[1551:1544]};
      mid_2[0] = {1'b0,layer_2_2[1535:1528]} - {1'b0, layer_1_2[1535:1528]};
      mid_2[1] = {1'b0,layer_2_2[1543:1536]} - {1'b0, layer_1_2[1543:1536]};
      mid_2[2] = {1'b0,layer_2_2[1551:1544]} - {1'b0, layer_1_2[1551:1544]};
      btm_0[0] = {1'b0,layer_3_0[1535:1528]} - {1'b0, layer_2_0[1535:1528]};
      btm_0[1] = {1'b0,layer_3_0[1543:1536]} - {1'b0, layer_2_0[1543:1536]};
      btm_0[2] = {1'b0,layer_3_0[1551:1544]} - {1'b0, layer_2_0[1551:1544]};
      btm_1[0] = {1'b0,layer_3_1[1535:1528]} - {1'b0, layer_2_1[1535:1528]};
      btm_1[1] = {1'b0,layer_3_1[1543:1536]} - {1'b0, layer_2_1[1543:1536]};
      btm_1[2] = {1'b0,layer_3_1[1551:1544]} - {1'b0, layer_2_1[1551:1544]};
      btm_2[0] = {1'b0,layer_3_2[1535:1528]} - {1'b0, layer_2_2[1535:1528]};
      btm_2[1] = {1'b0,layer_3_2[1543:1536]} - {1'b0, layer_2_2[1543:1536]};
      btm_2[2] = {1'b0,layer_3_2[1551:1544]} - {1'b0, layer_2_2[1551:1544]};
    end
    'd193: begin
      top_0[0] = {1'b0,layer_1_0[1543:1536]} - {1'b0, layer_0_0[1543:1536]};
      top_0[1] = {1'b0,layer_1_0[1551:1544]} - {1'b0, layer_0_0[1551:1544]};
      top_0[2] = {1'b0,layer_1_0[1559:1552]} - {1'b0, layer_0_0[1559:1552]};
      top_1[0] = {1'b0,layer_1_1[1543:1536]} - {1'b0, layer_0_1[1543:1536]};
      top_1[1] = {1'b0,layer_1_1[1551:1544]} - {1'b0, layer_0_1[1551:1544]};
      top_1[2] = {1'b0,layer_1_1[1559:1552]} - {1'b0, layer_0_1[1559:1552]};
      top_2[0] = {1'b0,layer_1_2[1543:1536]} - {1'b0, layer_0_2[1543:1536]};
      top_2[1] = {1'b0,layer_1_2[1551:1544]} - {1'b0, layer_0_2[1551:1544]};
      top_2[2] = {1'b0,layer_1_2[1559:1552]} - {1'b0, layer_0_2[1559:1552]};
      mid_0[0] = {1'b0,layer_2_0[1543:1536]} - {1'b0, layer_1_0[1543:1536]};
      mid_0[1] = {1'b0,layer_2_0[1551:1544]} - {1'b0, layer_1_0[1551:1544]};
      mid_0[2] = {1'b0,layer_2_0[1559:1552]} - {1'b0, layer_1_0[1559:1552]};
      mid_1[0] = {1'b0,layer_2_1[1543:1536]} - {1'b0, layer_1_1[1543:1536]};
      mid_1[1] = {1'b0,layer_2_1[1551:1544]} - {1'b0, layer_1_1[1551:1544]};
      mid_1[2] = {1'b0,layer_2_1[1559:1552]} - {1'b0, layer_1_1[1559:1552]};
      mid_2[0] = {1'b0,layer_2_2[1543:1536]} - {1'b0, layer_1_2[1543:1536]};
      mid_2[1] = {1'b0,layer_2_2[1551:1544]} - {1'b0, layer_1_2[1551:1544]};
      mid_2[2] = {1'b0,layer_2_2[1559:1552]} - {1'b0, layer_1_2[1559:1552]};
      btm_0[0] = {1'b0,layer_3_0[1543:1536]} - {1'b0, layer_2_0[1543:1536]};
      btm_0[1] = {1'b0,layer_3_0[1551:1544]} - {1'b0, layer_2_0[1551:1544]};
      btm_0[2] = {1'b0,layer_3_0[1559:1552]} - {1'b0, layer_2_0[1559:1552]};
      btm_1[0] = {1'b0,layer_3_1[1543:1536]} - {1'b0, layer_2_1[1543:1536]};
      btm_1[1] = {1'b0,layer_3_1[1551:1544]} - {1'b0, layer_2_1[1551:1544]};
      btm_1[2] = {1'b0,layer_3_1[1559:1552]} - {1'b0, layer_2_1[1559:1552]};
      btm_2[0] = {1'b0,layer_3_2[1543:1536]} - {1'b0, layer_2_2[1543:1536]};
      btm_2[1] = {1'b0,layer_3_2[1551:1544]} - {1'b0, layer_2_2[1551:1544]};
      btm_2[2] = {1'b0,layer_3_2[1559:1552]} - {1'b0, layer_2_2[1559:1552]};
    end
    'd194: begin
      top_0[0] = {1'b0,layer_1_0[1551:1544]} - {1'b0, layer_0_0[1551:1544]};
      top_0[1] = {1'b0,layer_1_0[1559:1552]} - {1'b0, layer_0_0[1559:1552]};
      top_0[2] = {1'b0,layer_1_0[1567:1560]} - {1'b0, layer_0_0[1567:1560]};
      top_1[0] = {1'b0,layer_1_1[1551:1544]} - {1'b0, layer_0_1[1551:1544]};
      top_1[1] = {1'b0,layer_1_1[1559:1552]} - {1'b0, layer_0_1[1559:1552]};
      top_1[2] = {1'b0,layer_1_1[1567:1560]} - {1'b0, layer_0_1[1567:1560]};
      top_2[0] = {1'b0,layer_1_2[1551:1544]} - {1'b0, layer_0_2[1551:1544]};
      top_2[1] = {1'b0,layer_1_2[1559:1552]} - {1'b0, layer_0_2[1559:1552]};
      top_2[2] = {1'b0,layer_1_2[1567:1560]} - {1'b0, layer_0_2[1567:1560]};
      mid_0[0] = {1'b0,layer_2_0[1551:1544]} - {1'b0, layer_1_0[1551:1544]};
      mid_0[1] = {1'b0,layer_2_0[1559:1552]} - {1'b0, layer_1_0[1559:1552]};
      mid_0[2] = {1'b0,layer_2_0[1567:1560]} - {1'b0, layer_1_0[1567:1560]};
      mid_1[0] = {1'b0,layer_2_1[1551:1544]} - {1'b0, layer_1_1[1551:1544]};
      mid_1[1] = {1'b0,layer_2_1[1559:1552]} - {1'b0, layer_1_1[1559:1552]};
      mid_1[2] = {1'b0,layer_2_1[1567:1560]} - {1'b0, layer_1_1[1567:1560]};
      mid_2[0] = {1'b0,layer_2_2[1551:1544]} - {1'b0, layer_1_2[1551:1544]};
      mid_2[1] = {1'b0,layer_2_2[1559:1552]} - {1'b0, layer_1_2[1559:1552]};
      mid_2[2] = {1'b0,layer_2_2[1567:1560]} - {1'b0, layer_1_2[1567:1560]};
      btm_0[0] = {1'b0,layer_3_0[1551:1544]} - {1'b0, layer_2_0[1551:1544]};
      btm_0[1] = {1'b0,layer_3_0[1559:1552]} - {1'b0, layer_2_0[1559:1552]};
      btm_0[2] = {1'b0,layer_3_0[1567:1560]} - {1'b0, layer_2_0[1567:1560]};
      btm_1[0] = {1'b0,layer_3_1[1551:1544]} - {1'b0, layer_2_1[1551:1544]};
      btm_1[1] = {1'b0,layer_3_1[1559:1552]} - {1'b0, layer_2_1[1559:1552]};
      btm_1[2] = {1'b0,layer_3_1[1567:1560]} - {1'b0, layer_2_1[1567:1560]};
      btm_2[0] = {1'b0,layer_3_2[1551:1544]} - {1'b0, layer_2_2[1551:1544]};
      btm_2[1] = {1'b0,layer_3_2[1559:1552]} - {1'b0, layer_2_2[1559:1552]};
      btm_2[2] = {1'b0,layer_3_2[1567:1560]} - {1'b0, layer_2_2[1567:1560]};
    end
    'd195: begin
      top_0[0] = {1'b0,layer_1_0[1559:1552]} - {1'b0, layer_0_0[1559:1552]};
      top_0[1] = {1'b0,layer_1_0[1567:1560]} - {1'b0, layer_0_0[1567:1560]};
      top_0[2] = {1'b0,layer_1_0[1575:1568]} - {1'b0, layer_0_0[1575:1568]};
      top_1[0] = {1'b0,layer_1_1[1559:1552]} - {1'b0, layer_0_1[1559:1552]};
      top_1[1] = {1'b0,layer_1_1[1567:1560]} - {1'b0, layer_0_1[1567:1560]};
      top_1[2] = {1'b0,layer_1_1[1575:1568]} - {1'b0, layer_0_1[1575:1568]};
      top_2[0] = {1'b0,layer_1_2[1559:1552]} - {1'b0, layer_0_2[1559:1552]};
      top_2[1] = {1'b0,layer_1_2[1567:1560]} - {1'b0, layer_0_2[1567:1560]};
      top_2[2] = {1'b0,layer_1_2[1575:1568]} - {1'b0, layer_0_2[1575:1568]};
      mid_0[0] = {1'b0,layer_2_0[1559:1552]} - {1'b0, layer_1_0[1559:1552]};
      mid_0[1] = {1'b0,layer_2_0[1567:1560]} - {1'b0, layer_1_0[1567:1560]};
      mid_0[2] = {1'b0,layer_2_0[1575:1568]} - {1'b0, layer_1_0[1575:1568]};
      mid_1[0] = {1'b0,layer_2_1[1559:1552]} - {1'b0, layer_1_1[1559:1552]};
      mid_1[1] = {1'b0,layer_2_1[1567:1560]} - {1'b0, layer_1_1[1567:1560]};
      mid_1[2] = {1'b0,layer_2_1[1575:1568]} - {1'b0, layer_1_1[1575:1568]};
      mid_2[0] = {1'b0,layer_2_2[1559:1552]} - {1'b0, layer_1_2[1559:1552]};
      mid_2[1] = {1'b0,layer_2_2[1567:1560]} - {1'b0, layer_1_2[1567:1560]};
      mid_2[2] = {1'b0,layer_2_2[1575:1568]} - {1'b0, layer_1_2[1575:1568]};
      btm_0[0] = {1'b0,layer_3_0[1559:1552]} - {1'b0, layer_2_0[1559:1552]};
      btm_0[1] = {1'b0,layer_3_0[1567:1560]} - {1'b0, layer_2_0[1567:1560]};
      btm_0[2] = {1'b0,layer_3_0[1575:1568]} - {1'b0, layer_2_0[1575:1568]};
      btm_1[0] = {1'b0,layer_3_1[1559:1552]} - {1'b0, layer_2_1[1559:1552]};
      btm_1[1] = {1'b0,layer_3_1[1567:1560]} - {1'b0, layer_2_1[1567:1560]};
      btm_1[2] = {1'b0,layer_3_1[1575:1568]} - {1'b0, layer_2_1[1575:1568]};
      btm_2[0] = {1'b0,layer_3_2[1559:1552]} - {1'b0, layer_2_2[1559:1552]};
      btm_2[1] = {1'b0,layer_3_2[1567:1560]} - {1'b0, layer_2_2[1567:1560]};
      btm_2[2] = {1'b0,layer_3_2[1575:1568]} - {1'b0, layer_2_2[1575:1568]};
    end
    'd196: begin
      top_0[0] = {1'b0,layer_1_0[1567:1560]} - {1'b0, layer_0_0[1567:1560]};
      top_0[1] = {1'b0,layer_1_0[1575:1568]} - {1'b0, layer_0_0[1575:1568]};
      top_0[2] = {1'b0,layer_1_0[1583:1576]} - {1'b0, layer_0_0[1583:1576]};
      top_1[0] = {1'b0,layer_1_1[1567:1560]} - {1'b0, layer_0_1[1567:1560]};
      top_1[1] = {1'b0,layer_1_1[1575:1568]} - {1'b0, layer_0_1[1575:1568]};
      top_1[2] = {1'b0,layer_1_1[1583:1576]} - {1'b0, layer_0_1[1583:1576]};
      top_2[0] = {1'b0,layer_1_2[1567:1560]} - {1'b0, layer_0_2[1567:1560]};
      top_2[1] = {1'b0,layer_1_2[1575:1568]} - {1'b0, layer_0_2[1575:1568]};
      top_2[2] = {1'b0,layer_1_2[1583:1576]} - {1'b0, layer_0_2[1583:1576]};
      mid_0[0] = {1'b0,layer_2_0[1567:1560]} - {1'b0, layer_1_0[1567:1560]};
      mid_0[1] = {1'b0,layer_2_0[1575:1568]} - {1'b0, layer_1_0[1575:1568]};
      mid_0[2] = {1'b0,layer_2_0[1583:1576]} - {1'b0, layer_1_0[1583:1576]};
      mid_1[0] = {1'b0,layer_2_1[1567:1560]} - {1'b0, layer_1_1[1567:1560]};
      mid_1[1] = {1'b0,layer_2_1[1575:1568]} - {1'b0, layer_1_1[1575:1568]};
      mid_1[2] = {1'b0,layer_2_1[1583:1576]} - {1'b0, layer_1_1[1583:1576]};
      mid_2[0] = {1'b0,layer_2_2[1567:1560]} - {1'b0, layer_1_2[1567:1560]};
      mid_2[1] = {1'b0,layer_2_2[1575:1568]} - {1'b0, layer_1_2[1575:1568]};
      mid_2[2] = {1'b0,layer_2_2[1583:1576]} - {1'b0, layer_1_2[1583:1576]};
      btm_0[0] = {1'b0,layer_3_0[1567:1560]} - {1'b0, layer_2_0[1567:1560]};
      btm_0[1] = {1'b0,layer_3_0[1575:1568]} - {1'b0, layer_2_0[1575:1568]};
      btm_0[2] = {1'b0,layer_3_0[1583:1576]} - {1'b0, layer_2_0[1583:1576]};
      btm_1[0] = {1'b0,layer_3_1[1567:1560]} - {1'b0, layer_2_1[1567:1560]};
      btm_1[1] = {1'b0,layer_3_1[1575:1568]} - {1'b0, layer_2_1[1575:1568]};
      btm_1[2] = {1'b0,layer_3_1[1583:1576]} - {1'b0, layer_2_1[1583:1576]};
      btm_2[0] = {1'b0,layer_3_2[1567:1560]} - {1'b0, layer_2_2[1567:1560]};
      btm_2[1] = {1'b0,layer_3_2[1575:1568]} - {1'b0, layer_2_2[1575:1568]};
      btm_2[2] = {1'b0,layer_3_2[1583:1576]} - {1'b0, layer_2_2[1583:1576]};
    end
    'd197: begin
      top_0[0] = {1'b0,layer_1_0[1575:1568]} - {1'b0, layer_0_0[1575:1568]};
      top_0[1] = {1'b0,layer_1_0[1583:1576]} - {1'b0, layer_0_0[1583:1576]};
      top_0[2] = {1'b0,layer_1_0[1591:1584]} - {1'b0, layer_0_0[1591:1584]};
      top_1[0] = {1'b0,layer_1_1[1575:1568]} - {1'b0, layer_0_1[1575:1568]};
      top_1[1] = {1'b0,layer_1_1[1583:1576]} - {1'b0, layer_0_1[1583:1576]};
      top_1[2] = {1'b0,layer_1_1[1591:1584]} - {1'b0, layer_0_1[1591:1584]};
      top_2[0] = {1'b0,layer_1_2[1575:1568]} - {1'b0, layer_0_2[1575:1568]};
      top_2[1] = {1'b0,layer_1_2[1583:1576]} - {1'b0, layer_0_2[1583:1576]};
      top_2[2] = {1'b0,layer_1_2[1591:1584]} - {1'b0, layer_0_2[1591:1584]};
      mid_0[0] = {1'b0,layer_2_0[1575:1568]} - {1'b0, layer_1_0[1575:1568]};
      mid_0[1] = {1'b0,layer_2_0[1583:1576]} - {1'b0, layer_1_0[1583:1576]};
      mid_0[2] = {1'b0,layer_2_0[1591:1584]} - {1'b0, layer_1_0[1591:1584]};
      mid_1[0] = {1'b0,layer_2_1[1575:1568]} - {1'b0, layer_1_1[1575:1568]};
      mid_1[1] = {1'b0,layer_2_1[1583:1576]} - {1'b0, layer_1_1[1583:1576]};
      mid_1[2] = {1'b0,layer_2_1[1591:1584]} - {1'b0, layer_1_1[1591:1584]};
      mid_2[0] = {1'b0,layer_2_2[1575:1568]} - {1'b0, layer_1_2[1575:1568]};
      mid_2[1] = {1'b0,layer_2_2[1583:1576]} - {1'b0, layer_1_2[1583:1576]};
      mid_2[2] = {1'b0,layer_2_2[1591:1584]} - {1'b0, layer_1_2[1591:1584]};
      btm_0[0] = {1'b0,layer_3_0[1575:1568]} - {1'b0, layer_2_0[1575:1568]};
      btm_0[1] = {1'b0,layer_3_0[1583:1576]} - {1'b0, layer_2_0[1583:1576]};
      btm_0[2] = {1'b0,layer_3_0[1591:1584]} - {1'b0, layer_2_0[1591:1584]};
      btm_1[0] = {1'b0,layer_3_1[1575:1568]} - {1'b0, layer_2_1[1575:1568]};
      btm_1[1] = {1'b0,layer_3_1[1583:1576]} - {1'b0, layer_2_1[1583:1576]};
      btm_1[2] = {1'b0,layer_3_1[1591:1584]} - {1'b0, layer_2_1[1591:1584]};
      btm_2[0] = {1'b0,layer_3_2[1575:1568]} - {1'b0, layer_2_2[1575:1568]};
      btm_2[1] = {1'b0,layer_3_2[1583:1576]} - {1'b0, layer_2_2[1583:1576]};
      btm_2[2] = {1'b0,layer_3_2[1591:1584]} - {1'b0, layer_2_2[1591:1584]};
    end
    'd198: begin
      top_0[0] = {1'b0,layer_1_0[1583:1576]} - {1'b0, layer_0_0[1583:1576]};
      top_0[1] = {1'b0,layer_1_0[1591:1584]} - {1'b0, layer_0_0[1591:1584]};
      top_0[2] = {1'b0,layer_1_0[1599:1592]} - {1'b0, layer_0_0[1599:1592]};
      top_1[0] = {1'b0,layer_1_1[1583:1576]} - {1'b0, layer_0_1[1583:1576]};
      top_1[1] = {1'b0,layer_1_1[1591:1584]} - {1'b0, layer_0_1[1591:1584]};
      top_1[2] = {1'b0,layer_1_1[1599:1592]} - {1'b0, layer_0_1[1599:1592]};
      top_2[0] = {1'b0,layer_1_2[1583:1576]} - {1'b0, layer_0_2[1583:1576]};
      top_2[1] = {1'b0,layer_1_2[1591:1584]} - {1'b0, layer_0_2[1591:1584]};
      top_2[2] = {1'b0,layer_1_2[1599:1592]} - {1'b0, layer_0_2[1599:1592]};
      mid_0[0] = {1'b0,layer_2_0[1583:1576]} - {1'b0, layer_1_0[1583:1576]};
      mid_0[1] = {1'b0,layer_2_0[1591:1584]} - {1'b0, layer_1_0[1591:1584]};
      mid_0[2] = {1'b0,layer_2_0[1599:1592]} - {1'b0, layer_1_0[1599:1592]};
      mid_1[0] = {1'b0,layer_2_1[1583:1576]} - {1'b0, layer_1_1[1583:1576]};
      mid_1[1] = {1'b0,layer_2_1[1591:1584]} - {1'b0, layer_1_1[1591:1584]};
      mid_1[2] = {1'b0,layer_2_1[1599:1592]} - {1'b0, layer_1_1[1599:1592]};
      mid_2[0] = {1'b0,layer_2_2[1583:1576]} - {1'b0, layer_1_2[1583:1576]};
      mid_2[1] = {1'b0,layer_2_2[1591:1584]} - {1'b0, layer_1_2[1591:1584]};
      mid_2[2] = {1'b0,layer_2_2[1599:1592]} - {1'b0, layer_1_2[1599:1592]};
      btm_0[0] = {1'b0,layer_3_0[1583:1576]} - {1'b0, layer_2_0[1583:1576]};
      btm_0[1] = {1'b0,layer_3_0[1591:1584]} - {1'b0, layer_2_0[1591:1584]};
      btm_0[2] = {1'b0,layer_3_0[1599:1592]} - {1'b0, layer_2_0[1599:1592]};
      btm_1[0] = {1'b0,layer_3_1[1583:1576]} - {1'b0, layer_2_1[1583:1576]};
      btm_1[1] = {1'b0,layer_3_1[1591:1584]} - {1'b0, layer_2_1[1591:1584]};
      btm_1[2] = {1'b0,layer_3_1[1599:1592]} - {1'b0, layer_2_1[1599:1592]};
      btm_2[0] = {1'b0,layer_3_2[1583:1576]} - {1'b0, layer_2_2[1583:1576]};
      btm_2[1] = {1'b0,layer_3_2[1591:1584]} - {1'b0, layer_2_2[1591:1584]};
      btm_2[2] = {1'b0,layer_3_2[1599:1592]} - {1'b0, layer_2_2[1599:1592]};
    end
    'd199: begin
      top_0[0] = {1'b0,layer_1_0[1591:1584]} - {1'b0, layer_0_0[1591:1584]};
      top_0[1] = {1'b0,layer_1_0[1599:1592]} - {1'b0, layer_0_0[1599:1592]};
      top_0[2] = {1'b0,layer_1_0[1607:1600]} - {1'b0, layer_0_0[1607:1600]};
      top_1[0] = {1'b0,layer_1_1[1591:1584]} - {1'b0, layer_0_1[1591:1584]};
      top_1[1] = {1'b0,layer_1_1[1599:1592]} - {1'b0, layer_0_1[1599:1592]};
      top_1[2] = {1'b0,layer_1_1[1607:1600]} - {1'b0, layer_0_1[1607:1600]};
      top_2[0] = {1'b0,layer_1_2[1591:1584]} - {1'b0, layer_0_2[1591:1584]};
      top_2[1] = {1'b0,layer_1_2[1599:1592]} - {1'b0, layer_0_2[1599:1592]};
      top_2[2] = {1'b0,layer_1_2[1607:1600]} - {1'b0, layer_0_2[1607:1600]};
      mid_0[0] = {1'b0,layer_2_0[1591:1584]} - {1'b0, layer_1_0[1591:1584]};
      mid_0[1] = {1'b0,layer_2_0[1599:1592]} - {1'b0, layer_1_0[1599:1592]};
      mid_0[2] = {1'b0,layer_2_0[1607:1600]} - {1'b0, layer_1_0[1607:1600]};
      mid_1[0] = {1'b0,layer_2_1[1591:1584]} - {1'b0, layer_1_1[1591:1584]};
      mid_1[1] = {1'b0,layer_2_1[1599:1592]} - {1'b0, layer_1_1[1599:1592]};
      mid_1[2] = {1'b0,layer_2_1[1607:1600]} - {1'b0, layer_1_1[1607:1600]};
      mid_2[0] = {1'b0,layer_2_2[1591:1584]} - {1'b0, layer_1_2[1591:1584]};
      mid_2[1] = {1'b0,layer_2_2[1599:1592]} - {1'b0, layer_1_2[1599:1592]};
      mid_2[2] = {1'b0,layer_2_2[1607:1600]} - {1'b0, layer_1_2[1607:1600]};
      btm_0[0] = {1'b0,layer_3_0[1591:1584]} - {1'b0, layer_2_0[1591:1584]};
      btm_0[1] = {1'b0,layer_3_0[1599:1592]} - {1'b0, layer_2_0[1599:1592]};
      btm_0[2] = {1'b0,layer_3_0[1607:1600]} - {1'b0, layer_2_0[1607:1600]};
      btm_1[0] = {1'b0,layer_3_1[1591:1584]} - {1'b0, layer_2_1[1591:1584]};
      btm_1[1] = {1'b0,layer_3_1[1599:1592]} - {1'b0, layer_2_1[1599:1592]};
      btm_1[2] = {1'b0,layer_3_1[1607:1600]} - {1'b0, layer_2_1[1607:1600]};
      btm_2[0] = {1'b0,layer_3_2[1591:1584]} - {1'b0, layer_2_2[1591:1584]};
      btm_2[1] = {1'b0,layer_3_2[1599:1592]} - {1'b0, layer_2_2[1599:1592]};
      btm_2[2] = {1'b0,layer_3_2[1607:1600]} - {1'b0, layer_2_2[1607:1600]};
    end
    'd200: begin
      top_0[0] = {1'b0,layer_1_0[1599:1592]} - {1'b0, layer_0_0[1599:1592]};
      top_0[1] = {1'b0,layer_1_0[1607:1600]} - {1'b0, layer_0_0[1607:1600]};
      top_0[2] = {1'b0,layer_1_0[1615:1608]} - {1'b0, layer_0_0[1615:1608]};
      top_1[0] = {1'b0,layer_1_1[1599:1592]} - {1'b0, layer_0_1[1599:1592]};
      top_1[1] = {1'b0,layer_1_1[1607:1600]} - {1'b0, layer_0_1[1607:1600]};
      top_1[2] = {1'b0,layer_1_1[1615:1608]} - {1'b0, layer_0_1[1615:1608]};
      top_2[0] = {1'b0,layer_1_2[1599:1592]} - {1'b0, layer_0_2[1599:1592]};
      top_2[1] = {1'b0,layer_1_2[1607:1600]} - {1'b0, layer_0_2[1607:1600]};
      top_2[2] = {1'b0,layer_1_2[1615:1608]} - {1'b0, layer_0_2[1615:1608]};
      mid_0[0] = {1'b0,layer_2_0[1599:1592]} - {1'b0, layer_1_0[1599:1592]};
      mid_0[1] = {1'b0,layer_2_0[1607:1600]} - {1'b0, layer_1_0[1607:1600]};
      mid_0[2] = {1'b0,layer_2_0[1615:1608]} - {1'b0, layer_1_0[1615:1608]};
      mid_1[0] = {1'b0,layer_2_1[1599:1592]} - {1'b0, layer_1_1[1599:1592]};
      mid_1[1] = {1'b0,layer_2_1[1607:1600]} - {1'b0, layer_1_1[1607:1600]};
      mid_1[2] = {1'b0,layer_2_1[1615:1608]} - {1'b0, layer_1_1[1615:1608]};
      mid_2[0] = {1'b0,layer_2_2[1599:1592]} - {1'b0, layer_1_2[1599:1592]};
      mid_2[1] = {1'b0,layer_2_2[1607:1600]} - {1'b0, layer_1_2[1607:1600]};
      mid_2[2] = {1'b0,layer_2_2[1615:1608]} - {1'b0, layer_1_2[1615:1608]};
      btm_0[0] = {1'b0,layer_3_0[1599:1592]} - {1'b0, layer_2_0[1599:1592]};
      btm_0[1] = {1'b0,layer_3_0[1607:1600]} - {1'b0, layer_2_0[1607:1600]};
      btm_0[2] = {1'b0,layer_3_0[1615:1608]} - {1'b0, layer_2_0[1615:1608]};
      btm_1[0] = {1'b0,layer_3_1[1599:1592]} - {1'b0, layer_2_1[1599:1592]};
      btm_1[1] = {1'b0,layer_3_1[1607:1600]} - {1'b0, layer_2_1[1607:1600]};
      btm_1[2] = {1'b0,layer_3_1[1615:1608]} - {1'b0, layer_2_1[1615:1608]};
      btm_2[0] = {1'b0,layer_3_2[1599:1592]} - {1'b0, layer_2_2[1599:1592]};
      btm_2[1] = {1'b0,layer_3_2[1607:1600]} - {1'b0, layer_2_2[1607:1600]};
      btm_2[2] = {1'b0,layer_3_2[1615:1608]} - {1'b0, layer_2_2[1615:1608]};
    end
    'd201: begin
      top_0[0] = {1'b0,layer_1_0[1607:1600]} - {1'b0, layer_0_0[1607:1600]};
      top_0[1] = {1'b0,layer_1_0[1615:1608]} - {1'b0, layer_0_0[1615:1608]};
      top_0[2] = {1'b0,layer_1_0[1623:1616]} - {1'b0, layer_0_0[1623:1616]};
      top_1[0] = {1'b0,layer_1_1[1607:1600]} - {1'b0, layer_0_1[1607:1600]};
      top_1[1] = {1'b0,layer_1_1[1615:1608]} - {1'b0, layer_0_1[1615:1608]};
      top_1[2] = {1'b0,layer_1_1[1623:1616]} - {1'b0, layer_0_1[1623:1616]};
      top_2[0] = {1'b0,layer_1_2[1607:1600]} - {1'b0, layer_0_2[1607:1600]};
      top_2[1] = {1'b0,layer_1_2[1615:1608]} - {1'b0, layer_0_2[1615:1608]};
      top_2[2] = {1'b0,layer_1_2[1623:1616]} - {1'b0, layer_0_2[1623:1616]};
      mid_0[0] = {1'b0,layer_2_0[1607:1600]} - {1'b0, layer_1_0[1607:1600]};
      mid_0[1] = {1'b0,layer_2_0[1615:1608]} - {1'b0, layer_1_0[1615:1608]};
      mid_0[2] = {1'b0,layer_2_0[1623:1616]} - {1'b0, layer_1_0[1623:1616]};
      mid_1[0] = {1'b0,layer_2_1[1607:1600]} - {1'b0, layer_1_1[1607:1600]};
      mid_1[1] = {1'b0,layer_2_1[1615:1608]} - {1'b0, layer_1_1[1615:1608]};
      mid_1[2] = {1'b0,layer_2_1[1623:1616]} - {1'b0, layer_1_1[1623:1616]};
      mid_2[0] = {1'b0,layer_2_2[1607:1600]} - {1'b0, layer_1_2[1607:1600]};
      mid_2[1] = {1'b0,layer_2_2[1615:1608]} - {1'b0, layer_1_2[1615:1608]};
      mid_2[2] = {1'b0,layer_2_2[1623:1616]} - {1'b0, layer_1_2[1623:1616]};
      btm_0[0] = {1'b0,layer_3_0[1607:1600]} - {1'b0, layer_2_0[1607:1600]};
      btm_0[1] = {1'b0,layer_3_0[1615:1608]} - {1'b0, layer_2_0[1615:1608]};
      btm_0[2] = {1'b0,layer_3_0[1623:1616]} - {1'b0, layer_2_0[1623:1616]};
      btm_1[0] = {1'b0,layer_3_1[1607:1600]} - {1'b0, layer_2_1[1607:1600]};
      btm_1[1] = {1'b0,layer_3_1[1615:1608]} - {1'b0, layer_2_1[1615:1608]};
      btm_1[2] = {1'b0,layer_3_1[1623:1616]} - {1'b0, layer_2_1[1623:1616]};
      btm_2[0] = {1'b0,layer_3_2[1607:1600]} - {1'b0, layer_2_2[1607:1600]};
      btm_2[1] = {1'b0,layer_3_2[1615:1608]} - {1'b0, layer_2_2[1615:1608]};
      btm_2[2] = {1'b0,layer_3_2[1623:1616]} - {1'b0, layer_2_2[1623:1616]};
    end
    'd202: begin
      top_0[0] = {1'b0,layer_1_0[1615:1608]} - {1'b0, layer_0_0[1615:1608]};
      top_0[1] = {1'b0,layer_1_0[1623:1616]} - {1'b0, layer_0_0[1623:1616]};
      top_0[2] = {1'b0,layer_1_0[1631:1624]} - {1'b0, layer_0_0[1631:1624]};
      top_1[0] = {1'b0,layer_1_1[1615:1608]} - {1'b0, layer_0_1[1615:1608]};
      top_1[1] = {1'b0,layer_1_1[1623:1616]} - {1'b0, layer_0_1[1623:1616]};
      top_1[2] = {1'b0,layer_1_1[1631:1624]} - {1'b0, layer_0_1[1631:1624]};
      top_2[0] = {1'b0,layer_1_2[1615:1608]} - {1'b0, layer_0_2[1615:1608]};
      top_2[1] = {1'b0,layer_1_2[1623:1616]} - {1'b0, layer_0_2[1623:1616]};
      top_2[2] = {1'b0,layer_1_2[1631:1624]} - {1'b0, layer_0_2[1631:1624]};
      mid_0[0] = {1'b0,layer_2_0[1615:1608]} - {1'b0, layer_1_0[1615:1608]};
      mid_0[1] = {1'b0,layer_2_0[1623:1616]} - {1'b0, layer_1_0[1623:1616]};
      mid_0[2] = {1'b0,layer_2_0[1631:1624]} - {1'b0, layer_1_0[1631:1624]};
      mid_1[0] = {1'b0,layer_2_1[1615:1608]} - {1'b0, layer_1_1[1615:1608]};
      mid_1[1] = {1'b0,layer_2_1[1623:1616]} - {1'b0, layer_1_1[1623:1616]};
      mid_1[2] = {1'b0,layer_2_1[1631:1624]} - {1'b0, layer_1_1[1631:1624]};
      mid_2[0] = {1'b0,layer_2_2[1615:1608]} - {1'b0, layer_1_2[1615:1608]};
      mid_2[1] = {1'b0,layer_2_2[1623:1616]} - {1'b0, layer_1_2[1623:1616]};
      mid_2[2] = {1'b0,layer_2_2[1631:1624]} - {1'b0, layer_1_2[1631:1624]};
      btm_0[0] = {1'b0,layer_3_0[1615:1608]} - {1'b0, layer_2_0[1615:1608]};
      btm_0[1] = {1'b0,layer_3_0[1623:1616]} - {1'b0, layer_2_0[1623:1616]};
      btm_0[2] = {1'b0,layer_3_0[1631:1624]} - {1'b0, layer_2_0[1631:1624]};
      btm_1[0] = {1'b0,layer_3_1[1615:1608]} - {1'b0, layer_2_1[1615:1608]};
      btm_1[1] = {1'b0,layer_3_1[1623:1616]} - {1'b0, layer_2_1[1623:1616]};
      btm_1[2] = {1'b0,layer_3_1[1631:1624]} - {1'b0, layer_2_1[1631:1624]};
      btm_2[0] = {1'b0,layer_3_2[1615:1608]} - {1'b0, layer_2_2[1615:1608]};
      btm_2[1] = {1'b0,layer_3_2[1623:1616]} - {1'b0, layer_2_2[1623:1616]};
      btm_2[2] = {1'b0,layer_3_2[1631:1624]} - {1'b0, layer_2_2[1631:1624]};
    end
    'd203: begin
      top_0[0] = {1'b0,layer_1_0[1623:1616]} - {1'b0, layer_0_0[1623:1616]};
      top_0[1] = {1'b0,layer_1_0[1631:1624]} - {1'b0, layer_0_0[1631:1624]};
      top_0[2] = {1'b0,layer_1_0[1639:1632]} - {1'b0, layer_0_0[1639:1632]};
      top_1[0] = {1'b0,layer_1_1[1623:1616]} - {1'b0, layer_0_1[1623:1616]};
      top_1[1] = {1'b0,layer_1_1[1631:1624]} - {1'b0, layer_0_1[1631:1624]};
      top_1[2] = {1'b0,layer_1_1[1639:1632]} - {1'b0, layer_0_1[1639:1632]};
      top_2[0] = {1'b0,layer_1_2[1623:1616]} - {1'b0, layer_0_2[1623:1616]};
      top_2[1] = {1'b0,layer_1_2[1631:1624]} - {1'b0, layer_0_2[1631:1624]};
      top_2[2] = {1'b0,layer_1_2[1639:1632]} - {1'b0, layer_0_2[1639:1632]};
      mid_0[0] = {1'b0,layer_2_0[1623:1616]} - {1'b0, layer_1_0[1623:1616]};
      mid_0[1] = {1'b0,layer_2_0[1631:1624]} - {1'b0, layer_1_0[1631:1624]};
      mid_0[2] = {1'b0,layer_2_0[1639:1632]} - {1'b0, layer_1_0[1639:1632]};
      mid_1[0] = {1'b0,layer_2_1[1623:1616]} - {1'b0, layer_1_1[1623:1616]};
      mid_1[1] = {1'b0,layer_2_1[1631:1624]} - {1'b0, layer_1_1[1631:1624]};
      mid_1[2] = {1'b0,layer_2_1[1639:1632]} - {1'b0, layer_1_1[1639:1632]};
      mid_2[0] = {1'b0,layer_2_2[1623:1616]} - {1'b0, layer_1_2[1623:1616]};
      mid_2[1] = {1'b0,layer_2_2[1631:1624]} - {1'b0, layer_1_2[1631:1624]};
      mid_2[2] = {1'b0,layer_2_2[1639:1632]} - {1'b0, layer_1_2[1639:1632]};
      btm_0[0] = {1'b0,layer_3_0[1623:1616]} - {1'b0, layer_2_0[1623:1616]};
      btm_0[1] = {1'b0,layer_3_0[1631:1624]} - {1'b0, layer_2_0[1631:1624]};
      btm_0[2] = {1'b0,layer_3_0[1639:1632]} - {1'b0, layer_2_0[1639:1632]};
      btm_1[0] = {1'b0,layer_3_1[1623:1616]} - {1'b0, layer_2_1[1623:1616]};
      btm_1[1] = {1'b0,layer_3_1[1631:1624]} - {1'b0, layer_2_1[1631:1624]};
      btm_1[2] = {1'b0,layer_3_1[1639:1632]} - {1'b0, layer_2_1[1639:1632]};
      btm_2[0] = {1'b0,layer_3_2[1623:1616]} - {1'b0, layer_2_2[1623:1616]};
      btm_2[1] = {1'b0,layer_3_2[1631:1624]} - {1'b0, layer_2_2[1631:1624]};
      btm_2[2] = {1'b0,layer_3_2[1639:1632]} - {1'b0, layer_2_2[1639:1632]};
    end
    'd204: begin
      top_0[0] = {1'b0,layer_1_0[1631:1624]} - {1'b0, layer_0_0[1631:1624]};
      top_0[1] = {1'b0,layer_1_0[1639:1632]} - {1'b0, layer_0_0[1639:1632]};
      top_0[2] = {1'b0,layer_1_0[1647:1640]} - {1'b0, layer_0_0[1647:1640]};
      top_1[0] = {1'b0,layer_1_1[1631:1624]} - {1'b0, layer_0_1[1631:1624]};
      top_1[1] = {1'b0,layer_1_1[1639:1632]} - {1'b0, layer_0_1[1639:1632]};
      top_1[2] = {1'b0,layer_1_1[1647:1640]} - {1'b0, layer_0_1[1647:1640]};
      top_2[0] = {1'b0,layer_1_2[1631:1624]} - {1'b0, layer_0_2[1631:1624]};
      top_2[1] = {1'b0,layer_1_2[1639:1632]} - {1'b0, layer_0_2[1639:1632]};
      top_2[2] = {1'b0,layer_1_2[1647:1640]} - {1'b0, layer_0_2[1647:1640]};
      mid_0[0] = {1'b0,layer_2_0[1631:1624]} - {1'b0, layer_1_0[1631:1624]};
      mid_0[1] = {1'b0,layer_2_0[1639:1632]} - {1'b0, layer_1_0[1639:1632]};
      mid_0[2] = {1'b0,layer_2_0[1647:1640]} - {1'b0, layer_1_0[1647:1640]};
      mid_1[0] = {1'b0,layer_2_1[1631:1624]} - {1'b0, layer_1_1[1631:1624]};
      mid_1[1] = {1'b0,layer_2_1[1639:1632]} - {1'b0, layer_1_1[1639:1632]};
      mid_1[2] = {1'b0,layer_2_1[1647:1640]} - {1'b0, layer_1_1[1647:1640]};
      mid_2[0] = {1'b0,layer_2_2[1631:1624]} - {1'b0, layer_1_2[1631:1624]};
      mid_2[1] = {1'b0,layer_2_2[1639:1632]} - {1'b0, layer_1_2[1639:1632]};
      mid_2[2] = {1'b0,layer_2_2[1647:1640]} - {1'b0, layer_1_2[1647:1640]};
      btm_0[0] = {1'b0,layer_3_0[1631:1624]} - {1'b0, layer_2_0[1631:1624]};
      btm_0[1] = {1'b0,layer_3_0[1639:1632]} - {1'b0, layer_2_0[1639:1632]};
      btm_0[2] = {1'b0,layer_3_0[1647:1640]} - {1'b0, layer_2_0[1647:1640]};
      btm_1[0] = {1'b0,layer_3_1[1631:1624]} - {1'b0, layer_2_1[1631:1624]};
      btm_1[1] = {1'b0,layer_3_1[1639:1632]} - {1'b0, layer_2_1[1639:1632]};
      btm_1[2] = {1'b0,layer_3_1[1647:1640]} - {1'b0, layer_2_1[1647:1640]};
      btm_2[0] = {1'b0,layer_3_2[1631:1624]} - {1'b0, layer_2_2[1631:1624]};
      btm_2[1] = {1'b0,layer_3_2[1639:1632]} - {1'b0, layer_2_2[1639:1632]};
      btm_2[2] = {1'b0,layer_3_2[1647:1640]} - {1'b0, layer_2_2[1647:1640]};
    end
    'd205: begin
      top_0[0] = {1'b0,layer_1_0[1639:1632]} - {1'b0, layer_0_0[1639:1632]};
      top_0[1] = {1'b0,layer_1_0[1647:1640]} - {1'b0, layer_0_0[1647:1640]};
      top_0[2] = {1'b0,layer_1_0[1655:1648]} - {1'b0, layer_0_0[1655:1648]};
      top_1[0] = {1'b0,layer_1_1[1639:1632]} - {1'b0, layer_0_1[1639:1632]};
      top_1[1] = {1'b0,layer_1_1[1647:1640]} - {1'b0, layer_0_1[1647:1640]};
      top_1[2] = {1'b0,layer_1_1[1655:1648]} - {1'b0, layer_0_1[1655:1648]};
      top_2[0] = {1'b0,layer_1_2[1639:1632]} - {1'b0, layer_0_2[1639:1632]};
      top_2[1] = {1'b0,layer_1_2[1647:1640]} - {1'b0, layer_0_2[1647:1640]};
      top_2[2] = {1'b0,layer_1_2[1655:1648]} - {1'b0, layer_0_2[1655:1648]};
      mid_0[0] = {1'b0,layer_2_0[1639:1632]} - {1'b0, layer_1_0[1639:1632]};
      mid_0[1] = {1'b0,layer_2_0[1647:1640]} - {1'b0, layer_1_0[1647:1640]};
      mid_0[2] = {1'b0,layer_2_0[1655:1648]} - {1'b0, layer_1_0[1655:1648]};
      mid_1[0] = {1'b0,layer_2_1[1639:1632]} - {1'b0, layer_1_1[1639:1632]};
      mid_1[1] = {1'b0,layer_2_1[1647:1640]} - {1'b0, layer_1_1[1647:1640]};
      mid_1[2] = {1'b0,layer_2_1[1655:1648]} - {1'b0, layer_1_1[1655:1648]};
      mid_2[0] = {1'b0,layer_2_2[1639:1632]} - {1'b0, layer_1_2[1639:1632]};
      mid_2[1] = {1'b0,layer_2_2[1647:1640]} - {1'b0, layer_1_2[1647:1640]};
      mid_2[2] = {1'b0,layer_2_2[1655:1648]} - {1'b0, layer_1_2[1655:1648]};
      btm_0[0] = {1'b0,layer_3_0[1639:1632]} - {1'b0, layer_2_0[1639:1632]};
      btm_0[1] = {1'b0,layer_3_0[1647:1640]} - {1'b0, layer_2_0[1647:1640]};
      btm_0[2] = {1'b0,layer_3_0[1655:1648]} - {1'b0, layer_2_0[1655:1648]};
      btm_1[0] = {1'b0,layer_3_1[1639:1632]} - {1'b0, layer_2_1[1639:1632]};
      btm_1[1] = {1'b0,layer_3_1[1647:1640]} - {1'b0, layer_2_1[1647:1640]};
      btm_1[2] = {1'b0,layer_3_1[1655:1648]} - {1'b0, layer_2_1[1655:1648]};
      btm_2[0] = {1'b0,layer_3_2[1639:1632]} - {1'b0, layer_2_2[1639:1632]};
      btm_2[1] = {1'b0,layer_3_2[1647:1640]} - {1'b0, layer_2_2[1647:1640]};
      btm_2[2] = {1'b0,layer_3_2[1655:1648]} - {1'b0, layer_2_2[1655:1648]};
    end
    'd206: begin
      top_0[0] = {1'b0,layer_1_0[1647:1640]} - {1'b0, layer_0_0[1647:1640]};
      top_0[1] = {1'b0,layer_1_0[1655:1648]} - {1'b0, layer_0_0[1655:1648]};
      top_0[2] = {1'b0,layer_1_0[1663:1656]} - {1'b0, layer_0_0[1663:1656]};
      top_1[0] = {1'b0,layer_1_1[1647:1640]} - {1'b0, layer_0_1[1647:1640]};
      top_1[1] = {1'b0,layer_1_1[1655:1648]} - {1'b0, layer_0_1[1655:1648]};
      top_1[2] = {1'b0,layer_1_1[1663:1656]} - {1'b0, layer_0_1[1663:1656]};
      top_2[0] = {1'b0,layer_1_2[1647:1640]} - {1'b0, layer_0_2[1647:1640]};
      top_2[1] = {1'b0,layer_1_2[1655:1648]} - {1'b0, layer_0_2[1655:1648]};
      top_2[2] = {1'b0,layer_1_2[1663:1656]} - {1'b0, layer_0_2[1663:1656]};
      mid_0[0] = {1'b0,layer_2_0[1647:1640]} - {1'b0, layer_1_0[1647:1640]};
      mid_0[1] = {1'b0,layer_2_0[1655:1648]} - {1'b0, layer_1_0[1655:1648]};
      mid_0[2] = {1'b0,layer_2_0[1663:1656]} - {1'b0, layer_1_0[1663:1656]};
      mid_1[0] = {1'b0,layer_2_1[1647:1640]} - {1'b0, layer_1_1[1647:1640]};
      mid_1[1] = {1'b0,layer_2_1[1655:1648]} - {1'b0, layer_1_1[1655:1648]};
      mid_1[2] = {1'b0,layer_2_1[1663:1656]} - {1'b0, layer_1_1[1663:1656]};
      mid_2[0] = {1'b0,layer_2_2[1647:1640]} - {1'b0, layer_1_2[1647:1640]};
      mid_2[1] = {1'b0,layer_2_2[1655:1648]} - {1'b0, layer_1_2[1655:1648]};
      mid_2[2] = {1'b0,layer_2_2[1663:1656]} - {1'b0, layer_1_2[1663:1656]};
      btm_0[0] = {1'b0,layer_3_0[1647:1640]} - {1'b0, layer_2_0[1647:1640]};
      btm_0[1] = {1'b0,layer_3_0[1655:1648]} - {1'b0, layer_2_0[1655:1648]};
      btm_0[2] = {1'b0,layer_3_0[1663:1656]} - {1'b0, layer_2_0[1663:1656]};
      btm_1[0] = {1'b0,layer_3_1[1647:1640]} - {1'b0, layer_2_1[1647:1640]};
      btm_1[1] = {1'b0,layer_3_1[1655:1648]} - {1'b0, layer_2_1[1655:1648]};
      btm_1[2] = {1'b0,layer_3_1[1663:1656]} - {1'b0, layer_2_1[1663:1656]};
      btm_2[0] = {1'b0,layer_3_2[1647:1640]} - {1'b0, layer_2_2[1647:1640]};
      btm_2[1] = {1'b0,layer_3_2[1655:1648]} - {1'b0, layer_2_2[1655:1648]};
      btm_2[2] = {1'b0,layer_3_2[1663:1656]} - {1'b0, layer_2_2[1663:1656]};
    end
    'd207: begin
      top_0[0] = {1'b0,layer_1_0[1655:1648]} - {1'b0, layer_0_0[1655:1648]};
      top_0[1] = {1'b0,layer_1_0[1663:1656]} - {1'b0, layer_0_0[1663:1656]};
      top_0[2] = {1'b0,layer_1_0[1671:1664]} - {1'b0, layer_0_0[1671:1664]};
      top_1[0] = {1'b0,layer_1_1[1655:1648]} - {1'b0, layer_0_1[1655:1648]};
      top_1[1] = {1'b0,layer_1_1[1663:1656]} - {1'b0, layer_0_1[1663:1656]};
      top_1[2] = {1'b0,layer_1_1[1671:1664]} - {1'b0, layer_0_1[1671:1664]};
      top_2[0] = {1'b0,layer_1_2[1655:1648]} - {1'b0, layer_0_2[1655:1648]};
      top_2[1] = {1'b0,layer_1_2[1663:1656]} - {1'b0, layer_0_2[1663:1656]};
      top_2[2] = {1'b0,layer_1_2[1671:1664]} - {1'b0, layer_0_2[1671:1664]};
      mid_0[0] = {1'b0,layer_2_0[1655:1648]} - {1'b0, layer_1_0[1655:1648]};
      mid_0[1] = {1'b0,layer_2_0[1663:1656]} - {1'b0, layer_1_0[1663:1656]};
      mid_0[2] = {1'b0,layer_2_0[1671:1664]} - {1'b0, layer_1_0[1671:1664]};
      mid_1[0] = {1'b0,layer_2_1[1655:1648]} - {1'b0, layer_1_1[1655:1648]};
      mid_1[1] = {1'b0,layer_2_1[1663:1656]} - {1'b0, layer_1_1[1663:1656]};
      mid_1[2] = {1'b0,layer_2_1[1671:1664]} - {1'b0, layer_1_1[1671:1664]};
      mid_2[0] = {1'b0,layer_2_2[1655:1648]} - {1'b0, layer_1_2[1655:1648]};
      mid_2[1] = {1'b0,layer_2_2[1663:1656]} - {1'b0, layer_1_2[1663:1656]};
      mid_2[2] = {1'b0,layer_2_2[1671:1664]} - {1'b0, layer_1_2[1671:1664]};
      btm_0[0] = {1'b0,layer_3_0[1655:1648]} - {1'b0, layer_2_0[1655:1648]};
      btm_0[1] = {1'b0,layer_3_0[1663:1656]} - {1'b0, layer_2_0[1663:1656]};
      btm_0[2] = {1'b0,layer_3_0[1671:1664]} - {1'b0, layer_2_0[1671:1664]};
      btm_1[0] = {1'b0,layer_3_1[1655:1648]} - {1'b0, layer_2_1[1655:1648]};
      btm_1[1] = {1'b0,layer_3_1[1663:1656]} - {1'b0, layer_2_1[1663:1656]};
      btm_1[2] = {1'b0,layer_3_1[1671:1664]} - {1'b0, layer_2_1[1671:1664]};
      btm_2[0] = {1'b0,layer_3_2[1655:1648]} - {1'b0, layer_2_2[1655:1648]};
      btm_2[1] = {1'b0,layer_3_2[1663:1656]} - {1'b0, layer_2_2[1663:1656]};
      btm_2[2] = {1'b0,layer_3_2[1671:1664]} - {1'b0, layer_2_2[1671:1664]};
    end
    'd208: begin
      top_0[0] = {1'b0,layer_1_0[1663:1656]} - {1'b0, layer_0_0[1663:1656]};
      top_0[1] = {1'b0,layer_1_0[1671:1664]} - {1'b0, layer_0_0[1671:1664]};
      top_0[2] = {1'b0,layer_1_0[1679:1672]} - {1'b0, layer_0_0[1679:1672]};
      top_1[0] = {1'b0,layer_1_1[1663:1656]} - {1'b0, layer_0_1[1663:1656]};
      top_1[1] = {1'b0,layer_1_1[1671:1664]} - {1'b0, layer_0_1[1671:1664]};
      top_1[2] = {1'b0,layer_1_1[1679:1672]} - {1'b0, layer_0_1[1679:1672]};
      top_2[0] = {1'b0,layer_1_2[1663:1656]} - {1'b0, layer_0_2[1663:1656]};
      top_2[1] = {1'b0,layer_1_2[1671:1664]} - {1'b0, layer_0_2[1671:1664]};
      top_2[2] = {1'b0,layer_1_2[1679:1672]} - {1'b0, layer_0_2[1679:1672]};
      mid_0[0] = {1'b0,layer_2_0[1663:1656]} - {1'b0, layer_1_0[1663:1656]};
      mid_0[1] = {1'b0,layer_2_0[1671:1664]} - {1'b0, layer_1_0[1671:1664]};
      mid_0[2] = {1'b0,layer_2_0[1679:1672]} - {1'b0, layer_1_0[1679:1672]};
      mid_1[0] = {1'b0,layer_2_1[1663:1656]} - {1'b0, layer_1_1[1663:1656]};
      mid_1[1] = {1'b0,layer_2_1[1671:1664]} - {1'b0, layer_1_1[1671:1664]};
      mid_1[2] = {1'b0,layer_2_1[1679:1672]} - {1'b0, layer_1_1[1679:1672]};
      mid_2[0] = {1'b0,layer_2_2[1663:1656]} - {1'b0, layer_1_2[1663:1656]};
      mid_2[1] = {1'b0,layer_2_2[1671:1664]} - {1'b0, layer_1_2[1671:1664]};
      mid_2[2] = {1'b0,layer_2_2[1679:1672]} - {1'b0, layer_1_2[1679:1672]};
      btm_0[0] = {1'b0,layer_3_0[1663:1656]} - {1'b0, layer_2_0[1663:1656]};
      btm_0[1] = {1'b0,layer_3_0[1671:1664]} - {1'b0, layer_2_0[1671:1664]};
      btm_0[2] = {1'b0,layer_3_0[1679:1672]} - {1'b0, layer_2_0[1679:1672]};
      btm_1[0] = {1'b0,layer_3_1[1663:1656]} - {1'b0, layer_2_1[1663:1656]};
      btm_1[1] = {1'b0,layer_3_1[1671:1664]} - {1'b0, layer_2_1[1671:1664]};
      btm_1[2] = {1'b0,layer_3_1[1679:1672]} - {1'b0, layer_2_1[1679:1672]};
      btm_2[0] = {1'b0,layer_3_2[1663:1656]} - {1'b0, layer_2_2[1663:1656]};
      btm_2[1] = {1'b0,layer_3_2[1671:1664]} - {1'b0, layer_2_2[1671:1664]};
      btm_2[2] = {1'b0,layer_3_2[1679:1672]} - {1'b0, layer_2_2[1679:1672]};
    end
    'd209: begin
      top_0[0] = {1'b0,layer_1_0[1671:1664]} - {1'b0, layer_0_0[1671:1664]};
      top_0[1] = {1'b0,layer_1_0[1679:1672]} - {1'b0, layer_0_0[1679:1672]};
      top_0[2] = {1'b0,layer_1_0[1687:1680]} - {1'b0, layer_0_0[1687:1680]};
      top_1[0] = {1'b0,layer_1_1[1671:1664]} - {1'b0, layer_0_1[1671:1664]};
      top_1[1] = {1'b0,layer_1_1[1679:1672]} - {1'b0, layer_0_1[1679:1672]};
      top_1[2] = {1'b0,layer_1_1[1687:1680]} - {1'b0, layer_0_1[1687:1680]};
      top_2[0] = {1'b0,layer_1_2[1671:1664]} - {1'b0, layer_0_2[1671:1664]};
      top_2[1] = {1'b0,layer_1_2[1679:1672]} - {1'b0, layer_0_2[1679:1672]};
      top_2[2] = {1'b0,layer_1_2[1687:1680]} - {1'b0, layer_0_2[1687:1680]};
      mid_0[0] = {1'b0,layer_2_0[1671:1664]} - {1'b0, layer_1_0[1671:1664]};
      mid_0[1] = {1'b0,layer_2_0[1679:1672]} - {1'b0, layer_1_0[1679:1672]};
      mid_0[2] = {1'b0,layer_2_0[1687:1680]} - {1'b0, layer_1_0[1687:1680]};
      mid_1[0] = {1'b0,layer_2_1[1671:1664]} - {1'b0, layer_1_1[1671:1664]};
      mid_1[1] = {1'b0,layer_2_1[1679:1672]} - {1'b0, layer_1_1[1679:1672]};
      mid_1[2] = {1'b0,layer_2_1[1687:1680]} - {1'b0, layer_1_1[1687:1680]};
      mid_2[0] = {1'b0,layer_2_2[1671:1664]} - {1'b0, layer_1_2[1671:1664]};
      mid_2[1] = {1'b0,layer_2_2[1679:1672]} - {1'b0, layer_1_2[1679:1672]};
      mid_2[2] = {1'b0,layer_2_2[1687:1680]} - {1'b0, layer_1_2[1687:1680]};
      btm_0[0] = {1'b0,layer_3_0[1671:1664]} - {1'b0, layer_2_0[1671:1664]};
      btm_0[1] = {1'b0,layer_3_0[1679:1672]} - {1'b0, layer_2_0[1679:1672]};
      btm_0[2] = {1'b0,layer_3_0[1687:1680]} - {1'b0, layer_2_0[1687:1680]};
      btm_1[0] = {1'b0,layer_3_1[1671:1664]} - {1'b0, layer_2_1[1671:1664]};
      btm_1[1] = {1'b0,layer_3_1[1679:1672]} - {1'b0, layer_2_1[1679:1672]};
      btm_1[2] = {1'b0,layer_3_1[1687:1680]} - {1'b0, layer_2_1[1687:1680]};
      btm_2[0] = {1'b0,layer_3_2[1671:1664]} - {1'b0, layer_2_2[1671:1664]};
      btm_2[1] = {1'b0,layer_3_2[1679:1672]} - {1'b0, layer_2_2[1679:1672]};
      btm_2[2] = {1'b0,layer_3_2[1687:1680]} - {1'b0, layer_2_2[1687:1680]};
    end
    'd210: begin
      top_0[0] = {1'b0,layer_1_0[1679:1672]} - {1'b0, layer_0_0[1679:1672]};
      top_0[1] = {1'b0,layer_1_0[1687:1680]} - {1'b0, layer_0_0[1687:1680]};
      top_0[2] = {1'b0,layer_1_0[1695:1688]} - {1'b0, layer_0_0[1695:1688]};
      top_1[0] = {1'b0,layer_1_1[1679:1672]} - {1'b0, layer_0_1[1679:1672]};
      top_1[1] = {1'b0,layer_1_1[1687:1680]} - {1'b0, layer_0_1[1687:1680]};
      top_1[2] = {1'b0,layer_1_1[1695:1688]} - {1'b0, layer_0_1[1695:1688]};
      top_2[0] = {1'b0,layer_1_2[1679:1672]} - {1'b0, layer_0_2[1679:1672]};
      top_2[1] = {1'b0,layer_1_2[1687:1680]} - {1'b0, layer_0_2[1687:1680]};
      top_2[2] = {1'b0,layer_1_2[1695:1688]} - {1'b0, layer_0_2[1695:1688]};
      mid_0[0] = {1'b0,layer_2_0[1679:1672]} - {1'b0, layer_1_0[1679:1672]};
      mid_0[1] = {1'b0,layer_2_0[1687:1680]} - {1'b0, layer_1_0[1687:1680]};
      mid_0[2] = {1'b0,layer_2_0[1695:1688]} - {1'b0, layer_1_0[1695:1688]};
      mid_1[0] = {1'b0,layer_2_1[1679:1672]} - {1'b0, layer_1_1[1679:1672]};
      mid_1[1] = {1'b0,layer_2_1[1687:1680]} - {1'b0, layer_1_1[1687:1680]};
      mid_1[2] = {1'b0,layer_2_1[1695:1688]} - {1'b0, layer_1_1[1695:1688]};
      mid_2[0] = {1'b0,layer_2_2[1679:1672]} - {1'b0, layer_1_2[1679:1672]};
      mid_2[1] = {1'b0,layer_2_2[1687:1680]} - {1'b0, layer_1_2[1687:1680]};
      mid_2[2] = {1'b0,layer_2_2[1695:1688]} - {1'b0, layer_1_2[1695:1688]};
      btm_0[0] = {1'b0,layer_3_0[1679:1672]} - {1'b0, layer_2_0[1679:1672]};
      btm_0[1] = {1'b0,layer_3_0[1687:1680]} - {1'b0, layer_2_0[1687:1680]};
      btm_0[2] = {1'b0,layer_3_0[1695:1688]} - {1'b0, layer_2_0[1695:1688]};
      btm_1[0] = {1'b0,layer_3_1[1679:1672]} - {1'b0, layer_2_1[1679:1672]};
      btm_1[1] = {1'b0,layer_3_1[1687:1680]} - {1'b0, layer_2_1[1687:1680]};
      btm_1[2] = {1'b0,layer_3_1[1695:1688]} - {1'b0, layer_2_1[1695:1688]};
      btm_2[0] = {1'b0,layer_3_2[1679:1672]} - {1'b0, layer_2_2[1679:1672]};
      btm_2[1] = {1'b0,layer_3_2[1687:1680]} - {1'b0, layer_2_2[1687:1680]};
      btm_2[2] = {1'b0,layer_3_2[1695:1688]} - {1'b0, layer_2_2[1695:1688]};
    end
    'd211: begin
      top_0[0] = {1'b0,layer_1_0[1687:1680]} - {1'b0, layer_0_0[1687:1680]};
      top_0[1] = {1'b0,layer_1_0[1695:1688]} - {1'b0, layer_0_0[1695:1688]};
      top_0[2] = {1'b0,layer_1_0[1703:1696]} - {1'b0, layer_0_0[1703:1696]};
      top_1[0] = {1'b0,layer_1_1[1687:1680]} - {1'b0, layer_0_1[1687:1680]};
      top_1[1] = {1'b0,layer_1_1[1695:1688]} - {1'b0, layer_0_1[1695:1688]};
      top_1[2] = {1'b0,layer_1_1[1703:1696]} - {1'b0, layer_0_1[1703:1696]};
      top_2[0] = {1'b0,layer_1_2[1687:1680]} - {1'b0, layer_0_2[1687:1680]};
      top_2[1] = {1'b0,layer_1_2[1695:1688]} - {1'b0, layer_0_2[1695:1688]};
      top_2[2] = {1'b0,layer_1_2[1703:1696]} - {1'b0, layer_0_2[1703:1696]};
      mid_0[0] = {1'b0,layer_2_0[1687:1680]} - {1'b0, layer_1_0[1687:1680]};
      mid_0[1] = {1'b0,layer_2_0[1695:1688]} - {1'b0, layer_1_0[1695:1688]};
      mid_0[2] = {1'b0,layer_2_0[1703:1696]} - {1'b0, layer_1_0[1703:1696]};
      mid_1[0] = {1'b0,layer_2_1[1687:1680]} - {1'b0, layer_1_1[1687:1680]};
      mid_1[1] = {1'b0,layer_2_1[1695:1688]} - {1'b0, layer_1_1[1695:1688]};
      mid_1[2] = {1'b0,layer_2_1[1703:1696]} - {1'b0, layer_1_1[1703:1696]};
      mid_2[0] = {1'b0,layer_2_2[1687:1680]} - {1'b0, layer_1_2[1687:1680]};
      mid_2[1] = {1'b0,layer_2_2[1695:1688]} - {1'b0, layer_1_2[1695:1688]};
      mid_2[2] = {1'b0,layer_2_2[1703:1696]} - {1'b0, layer_1_2[1703:1696]};
      btm_0[0] = {1'b0,layer_3_0[1687:1680]} - {1'b0, layer_2_0[1687:1680]};
      btm_0[1] = {1'b0,layer_3_0[1695:1688]} - {1'b0, layer_2_0[1695:1688]};
      btm_0[2] = {1'b0,layer_3_0[1703:1696]} - {1'b0, layer_2_0[1703:1696]};
      btm_1[0] = {1'b0,layer_3_1[1687:1680]} - {1'b0, layer_2_1[1687:1680]};
      btm_1[1] = {1'b0,layer_3_1[1695:1688]} - {1'b0, layer_2_1[1695:1688]};
      btm_1[2] = {1'b0,layer_3_1[1703:1696]} - {1'b0, layer_2_1[1703:1696]};
      btm_2[0] = {1'b0,layer_3_2[1687:1680]} - {1'b0, layer_2_2[1687:1680]};
      btm_2[1] = {1'b0,layer_3_2[1695:1688]} - {1'b0, layer_2_2[1695:1688]};
      btm_2[2] = {1'b0,layer_3_2[1703:1696]} - {1'b0, layer_2_2[1703:1696]};
    end
    'd212: begin
      top_0[0] = {1'b0,layer_1_0[1695:1688]} - {1'b0, layer_0_0[1695:1688]};
      top_0[1] = {1'b0,layer_1_0[1703:1696]} - {1'b0, layer_0_0[1703:1696]};
      top_0[2] = {1'b0,layer_1_0[1711:1704]} - {1'b0, layer_0_0[1711:1704]};
      top_1[0] = {1'b0,layer_1_1[1695:1688]} - {1'b0, layer_0_1[1695:1688]};
      top_1[1] = {1'b0,layer_1_1[1703:1696]} - {1'b0, layer_0_1[1703:1696]};
      top_1[2] = {1'b0,layer_1_1[1711:1704]} - {1'b0, layer_0_1[1711:1704]};
      top_2[0] = {1'b0,layer_1_2[1695:1688]} - {1'b0, layer_0_2[1695:1688]};
      top_2[1] = {1'b0,layer_1_2[1703:1696]} - {1'b0, layer_0_2[1703:1696]};
      top_2[2] = {1'b0,layer_1_2[1711:1704]} - {1'b0, layer_0_2[1711:1704]};
      mid_0[0] = {1'b0,layer_2_0[1695:1688]} - {1'b0, layer_1_0[1695:1688]};
      mid_0[1] = {1'b0,layer_2_0[1703:1696]} - {1'b0, layer_1_0[1703:1696]};
      mid_0[2] = {1'b0,layer_2_0[1711:1704]} - {1'b0, layer_1_0[1711:1704]};
      mid_1[0] = {1'b0,layer_2_1[1695:1688]} - {1'b0, layer_1_1[1695:1688]};
      mid_1[1] = {1'b0,layer_2_1[1703:1696]} - {1'b0, layer_1_1[1703:1696]};
      mid_1[2] = {1'b0,layer_2_1[1711:1704]} - {1'b0, layer_1_1[1711:1704]};
      mid_2[0] = {1'b0,layer_2_2[1695:1688]} - {1'b0, layer_1_2[1695:1688]};
      mid_2[1] = {1'b0,layer_2_2[1703:1696]} - {1'b0, layer_1_2[1703:1696]};
      mid_2[2] = {1'b0,layer_2_2[1711:1704]} - {1'b0, layer_1_2[1711:1704]};
      btm_0[0] = {1'b0,layer_3_0[1695:1688]} - {1'b0, layer_2_0[1695:1688]};
      btm_0[1] = {1'b0,layer_3_0[1703:1696]} - {1'b0, layer_2_0[1703:1696]};
      btm_0[2] = {1'b0,layer_3_0[1711:1704]} - {1'b0, layer_2_0[1711:1704]};
      btm_1[0] = {1'b0,layer_3_1[1695:1688]} - {1'b0, layer_2_1[1695:1688]};
      btm_1[1] = {1'b0,layer_3_1[1703:1696]} - {1'b0, layer_2_1[1703:1696]};
      btm_1[2] = {1'b0,layer_3_1[1711:1704]} - {1'b0, layer_2_1[1711:1704]};
      btm_2[0] = {1'b0,layer_3_2[1695:1688]} - {1'b0, layer_2_2[1695:1688]};
      btm_2[1] = {1'b0,layer_3_2[1703:1696]} - {1'b0, layer_2_2[1703:1696]};
      btm_2[2] = {1'b0,layer_3_2[1711:1704]} - {1'b0, layer_2_2[1711:1704]};
    end
    'd213: begin
      top_0[0] = {1'b0,layer_1_0[1703:1696]} - {1'b0, layer_0_0[1703:1696]};
      top_0[1] = {1'b0,layer_1_0[1711:1704]} - {1'b0, layer_0_0[1711:1704]};
      top_0[2] = {1'b0,layer_1_0[1719:1712]} - {1'b0, layer_0_0[1719:1712]};
      top_1[0] = {1'b0,layer_1_1[1703:1696]} - {1'b0, layer_0_1[1703:1696]};
      top_1[1] = {1'b0,layer_1_1[1711:1704]} - {1'b0, layer_0_1[1711:1704]};
      top_1[2] = {1'b0,layer_1_1[1719:1712]} - {1'b0, layer_0_1[1719:1712]};
      top_2[0] = {1'b0,layer_1_2[1703:1696]} - {1'b0, layer_0_2[1703:1696]};
      top_2[1] = {1'b0,layer_1_2[1711:1704]} - {1'b0, layer_0_2[1711:1704]};
      top_2[2] = {1'b0,layer_1_2[1719:1712]} - {1'b0, layer_0_2[1719:1712]};
      mid_0[0] = {1'b0,layer_2_0[1703:1696]} - {1'b0, layer_1_0[1703:1696]};
      mid_0[1] = {1'b0,layer_2_0[1711:1704]} - {1'b0, layer_1_0[1711:1704]};
      mid_0[2] = {1'b0,layer_2_0[1719:1712]} - {1'b0, layer_1_0[1719:1712]};
      mid_1[0] = {1'b0,layer_2_1[1703:1696]} - {1'b0, layer_1_1[1703:1696]};
      mid_1[1] = {1'b0,layer_2_1[1711:1704]} - {1'b0, layer_1_1[1711:1704]};
      mid_1[2] = {1'b0,layer_2_1[1719:1712]} - {1'b0, layer_1_1[1719:1712]};
      mid_2[0] = {1'b0,layer_2_2[1703:1696]} - {1'b0, layer_1_2[1703:1696]};
      mid_2[1] = {1'b0,layer_2_2[1711:1704]} - {1'b0, layer_1_2[1711:1704]};
      mid_2[2] = {1'b0,layer_2_2[1719:1712]} - {1'b0, layer_1_2[1719:1712]};
      btm_0[0] = {1'b0,layer_3_0[1703:1696]} - {1'b0, layer_2_0[1703:1696]};
      btm_0[1] = {1'b0,layer_3_0[1711:1704]} - {1'b0, layer_2_0[1711:1704]};
      btm_0[2] = {1'b0,layer_3_0[1719:1712]} - {1'b0, layer_2_0[1719:1712]};
      btm_1[0] = {1'b0,layer_3_1[1703:1696]} - {1'b0, layer_2_1[1703:1696]};
      btm_1[1] = {1'b0,layer_3_1[1711:1704]} - {1'b0, layer_2_1[1711:1704]};
      btm_1[2] = {1'b0,layer_3_1[1719:1712]} - {1'b0, layer_2_1[1719:1712]};
      btm_2[0] = {1'b0,layer_3_2[1703:1696]} - {1'b0, layer_2_2[1703:1696]};
      btm_2[1] = {1'b0,layer_3_2[1711:1704]} - {1'b0, layer_2_2[1711:1704]};
      btm_2[2] = {1'b0,layer_3_2[1719:1712]} - {1'b0, layer_2_2[1719:1712]};
    end
    'd214: begin
      top_0[0] = {1'b0,layer_1_0[1711:1704]} - {1'b0, layer_0_0[1711:1704]};
      top_0[1] = {1'b0,layer_1_0[1719:1712]} - {1'b0, layer_0_0[1719:1712]};
      top_0[2] = {1'b0,layer_1_0[1727:1720]} - {1'b0, layer_0_0[1727:1720]};
      top_1[0] = {1'b0,layer_1_1[1711:1704]} - {1'b0, layer_0_1[1711:1704]};
      top_1[1] = {1'b0,layer_1_1[1719:1712]} - {1'b0, layer_0_1[1719:1712]};
      top_1[2] = {1'b0,layer_1_1[1727:1720]} - {1'b0, layer_0_1[1727:1720]};
      top_2[0] = {1'b0,layer_1_2[1711:1704]} - {1'b0, layer_0_2[1711:1704]};
      top_2[1] = {1'b0,layer_1_2[1719:1712]} - {1'b0, layer_0_2[1719:1712]};
      top_2[2] = {1'b0,layer_1_2[1727:1720]} - {1'b0, layer_0_2[1727:1720]};
      mid_0[0] = {1'b0,layer_2_0[1711:1704]} - {1'b0, layer_1_0[1711:1704]};
      mid_0[1] = {1'b0,layer_2_0[1719:1712]} - {1'b0, layer_1_0[1719:1712]};
      mid_0[2] = {1'b0,layer_2_0[1727:1720]} - {1'b0, layer_1_0[1727:1720]};
      mid_1[0] = {1'b0,layer_2_1[1711:1704]} - {1'b0, layer_1_1[1711:1704]};
      mid_1[1] = {1'b0,layer_2_1[1719:1712]} - {1'b0, layer_1_1[1719:1712]};
      mid_1[2] = {1'b0,layer_2_1[1727:1720]} - {1'b0, layer_1_1[1727:1720]};
      mid_2[0] = {1'b0,layer_2_2[1711:1704]} - {1'b0, layer_1_2[1711:1704]};
      mid_2[1] = {1'b0,layer_2_2[1719:1712]} - {1'b0, layer_1_2[1719:1712]};
      mid_2[2] = {1'b0,layer_2_2[1727:1720]} - {1'b0, layer_1_2[1727:1720]};
      btm_0[0] = {1'b0,layer_3_0[1711:1704]} - {1'b0, layer_2_0[1711:1704]};
      btm_0[1] = {1'b0,layer_3_0[1719:1712]} - {1'b0, layer_2_0[1719:1712]};
      btm_0[2] = {1'b0,layer_3_0[1727:1720]} - {1'b0, layer_2_0[1727:1720]};
      btm_1[0] = {1'b0,layer_3_1[1711:1704]} - {1'b0, layer_2_1[1711:1704]};
      btm_1[1] = {1'b0,layer_3_1[1719:1712]} - {1'b0, layer_2_1[1719:1712]};
      btm_1[2] = {1'b0,layer_3_1[1727:1720]} - {1'b0, layer_2_1[1727:1720]};
      btm_2[0] = {1'b0,layer_3_2[1711:1704]} - {1'b0, layer_2_2[1711:1704]};
      btm_2[1] = {1'b0,layer_3_2[1719:1712]} - {1'b0, layer_2_2[1719:1712]};
      btm_2[2] = {1'b0,layer_3_2[1727:1720]} - {1'b0, layer_2_2[1727:1720]};
    end
    'd215: begin
      top_0[0] = {1'b0,layer_1_0[1719:1712]} - {1'b0, layer_0_0[1719:1712]};
      top_0[1] = {1'b0,layer_1_0[1727:1720]} - {1'b0, layer_0_0[1727:1720]};
      top_0[2] = {1'b0,layer_1_0[1735:1728]} - {1'b0, layer_0_0[1735:1728]};
      top_1[0] = {1'b0,layer_1_1[1719:1712]} - {1'b0, layer_0_1[1719:1712]};
      top_1[1] = {1'b0,layer_1_1[1727:1720]} - {1'b0, layer_0_1[1727:1720]};
      top_1[2] = {1'b0,layer_1_1[1735:1728]} - {1'b0, layer_0_1[1735:1728]};
      top_2[0] = {1'b0,layer_1_2[1719:1712]} - {1'b0, layer_0_2[1719:1712]};
      top_2[1] = {1'b0,layer_1_2[1727:1720]} - {1'b0, layer_0_2[1727:1720]};
      top_2[2] = {1'b0,layer_1_2[1735:1728]} - {1'b0, layer_0_2[1735:1728]};
      mid_0[0] = {1'b0,layer_2_0[1719:1712]} - {1'b0, layer_1_0[1719:1712]};
      mid_0[1] = {1'b0,layer_2_0[1727:1720]} - {1'b0, layer_1_0[1727:1720]};
      mid_0[2] = {1'b0,layer_2_0[1735:1728]} - {1'b0, layer_1_0[1735:1728]};
      mid_1[0] = {1'b0,layer_2_1[1719:1712]} - {1'b0, layer_1_1[1719:1712]};
      mid_1[1] = {1'b0,layer_2_1[1727:1720]} - {1'b0, layer_1_1[1727:1720]};
      mid_1[2] = {1'b0,layer_2_1[1735:1728]} - {1'b0, layer_1_1[1735:1728]};
      mid_2[0] = {1'b0,layer_2_2[1719:1712]} - {1'b0, layer_1_2[1719:1712]};
      mid_2[1] = {1'b0,layer_2_2[1727:1720]} - {1'b0, layer_1_2[1727:1720]};
      mid_2[2] = {1'b0,layer_2_2[1735:1728]} - {1'b0, layer_1_2[1735:1728]};
      btm_0[0] = {1'b0,layer_3_0[1719:1712]} - {1'b0, layer_2_0[1719:1712]};
      btm_0[1] = {1'b0,layer_3_0[1727:1720]} - {1'b0, layer_2_0[1727:1720]};
      btm_0[2] = {1'b0,layer_3_0[1735:1728]} - {1'b0, layer_2_0[1735:1728]};
      btm_1[0] = {1'b0,layer_3_1[1719:1712]} - {1'b0, layer_2_1[1719:1712]};
      btm_1[1] = {1'b0,layer_3_1[1727:1720]} - {1'b0, layer_2_1[1727:1720]};
      btm_1[2] = {1'b0,layer_3_1[1735:1728]} - {1'b0, layer_2_1[1735:1728]};
      btm_2[0] = {1'b0,layer_3_2[1719:1712]} - {1'b0, layer_2_2[1719:1712]};
      btm_2[1] = {1'b0,layer_3_2[1727:1720]} - {1'b0, layer_2_2[1727:1720]};
      btm_2[2] = {1'b0,layer_3_2[1735:1728]} - {1'b0, layer_2_2[1735:1728]};
    end
    'd216: begin
      top_0[0] = {1'b0,layer_1_0[1727:1720]} - {1'b0, layer_0_0[1727:1720]};
      top_0[1] = {1'b0,layer_1_0[1735:1728]} - {1'b0, layer_0_0[1735:1728]};
      top_0[2] = {1'b0,layer_1_0[1743:1736]} - {1'b0, layer_0_0[1743:1736]};
      top_1[0] = {1'b0,layer_1_1[1727:1720]} - {1'b0, layer_0_1[1727:1720]};
      top_1[1] = {1'b0,layer_1_1[1735:1728]} - {1'b0, layer_0_1[1735:1728]};
      top_1[2] = {1'b0,layer_1_1[1743:1736]} - {1'b0, layer_0_1[1743:1736]};
      top_2[0] = {1'b0,layer_1_2[1727:1720]} - {1'b0, layer_0_2[1727:1720]};
      top_2[1] = {1'b0,layer_1_2[1735:1728]} - {1'b0, layer_0_2[1735:1728]};
      top_2[2] = {1'b0,layer_1_2[1743:1736]} - {1'b0, layer_0_2[1743:1736]};
      mid_0[0] = {1'b0,layer_2_0[1727:1720]} - {1'b0, layer_1_0[1727:1720]};
      mid_0[1] = {1'b0,layer_2_0[1735:1728]} - {1'b0, layer_1_0[1735:1728]};
      mid_0[2] = {1'b0,layer_2_0[1743:1736]} - {1'b0, layer_1_0[1743:1736]};
      mid_1[0] = {1'b0,layer_2_1[1727:1720]} - {1'b0, layer_1_1[1727:1720]};
      mid_1[1] = {1'b0,layer_2_1[1735:1728]} - {1'b0, layer_1_1[1735:1728]};
      mid_1[2] = {1'b0,layer_2_1[1743:1736]} - {1'b0, layer_1_1[1743:1736]};
      mid_2[0] = {1'b0,layer_2_2[1727:1720]} - {1'b0, layer_1_2[1727:1720]};
      mid_2[1] = {1'b0,layer_2_2[1735:1728]} - {1'b0, layer_1_2[1735:1728]};
      mid_2[2] = {1'b0,layer_2_2[1743:1736]} - {1'b0, layer_1_2[1743:1736]};
      btm_0[0] = {1'b0,layer_3_0[1727:1720]} - {1'b0, layer_2_0[1727:1720]};
      btm_0[1] = {1'b0,layer_3_0[1735:1728]} - {1'b0, layer_2_0[1735:1728]};
      btm_0[2] = {1'b0,layer_3_0[1743:1736]} - {1'b0, layer_2_0[1743:1736]};
      btm_1[0] = {1'b0,layer_3_1[1727:1720]} - {1'b0, layer_2_1[1727:1720]};
      btm_1[1] = {1'b0,layer_3_1[1735:1728]} - {1'b0, layer_2_1[1735:1728]};
      btm_1[2] = {1'b0,layer_3_1[1743:1736]} - {1'b0, layer_2_1[1743:1736]};
      btm_2[0] = {1'b0,layer_3_2[1727:1720]} - {1'b0, layer_2_2[1727:1720]};
      btm_2[1] = {1'b0,layer_3_2[1735:1728]} - {1'b0, layer_2_2[1735:1728]};
      btm_2[2] = {1'b0,layer_3_2[1743:1736]} - {1'b0, layer_2_2[1743:1736]};
    end
    'd217: begin
      top_0[0] = {1'b0,layer_1_0[1735:1728]} - {1'b0, layer_0_0[1735:1728]};
      top_0[1] = {1'b0,layer_1_0[1743:1736]} - {1'b0, layer_0_0[1743:1736]};
      top_0[2] = {1'b0,layer_1_0[1751:1744]} - {1'b0, layer_0_0[1751:1744]};
      top_1[0] = {1'b0,layer_1_1[1735:1728]} - {1'b0, layer_0_1[1735:1728]};
      top_1[1] = {1'b0,layer_1_1[1743:1736]} - {1'b0, layer_0_1[1743:1736]};
      top_1[2] = {1'b0,layer_1_1[1751:1744]} - {1'b0, layer_0_1[1751:1744]};
      top_2[0] = {1'b0,layer_1_2[1735:1728]} - {1'b0, layer_0_2[1735:1728]};
      top_2[1] = {1'b0,layer_1_2[1743:1736]} - {1'b0, layer_0_2[1743:1736]};
      top_2[2] = {1'b0,layer_1_2[1751:1744]} - {1'b0, layer_0_2[1751:1744]};
      mid_0[0] = {1'b0,layer_2_0[1735:1728]} - {1'b0, layer_1_0[1735:1728]};
      mid_0[1] = {1'b0,layer_2_0[1743:1736]} - {1'b0, layer_1_0[1743:1736]};
      mid_0[2] = {1'b0,layer_2_0[1751:1744]} - {1'b0, layer_1_0[1751:1744]};
      mid_1[0] = {1'b0,layer_2_1[1735:1728]} - {1'b0, layer_1_1[1735:1728]};
      mid_1[1] = {1'b0,layer_2_1[1743:1736]} - {1'b0, layer_1_1[1743:1736]};
      mid_1[2] = {1'b0,layer_2_1[1751:1744]} - {1'b0, layer_1_1[1751:1744]};
      mid_2[0] = {1'b0,layer_2_2[1735:1728]} - {1'b0, layer_1_2[1735:1728]};
      mid_2[1] = {1'b0,layer_2_2[1743:1736]} - {1'b0, layer_1_2[1743:1736]};
      mid_2[2] = {1'b0,layer_2_2[1751:1744]} - {1'b0, layer_1_2[1751:1744]};
      btm_0[0] = {1'b0,layer_3_0[1735:1728]} - {1'b0, layer_2_0[1735:1728]};
      btm_0[1] = {1'b0,layer_3_0[1743:1736]} - {1'b0, layer_2_0[1743:1736]};
      btm_0[2] = {1'b0,layer_3_0[1751:1744]} - {1'b0, layer_2_0[1751:1744]};
      btm_1[0] = {1'b0,layer_3_1[1735:1728]} - {1'b0, layer_2_1[1735:1728]};
      btm_1[1] = {1'b0,layer_3_1[1743:1736]} - {1'b0, layer_2_1[1743:1736]};
      btm_1[2] = {1'b0,layer_3_1[1751:1744]} - {1'b0, layer_2_1[1751:1744]};
      btm_2[0] = {1'b0,layer_3_2[1735:1728]} - {1'b0, layer_2_2[1735:1728]};
      btm_2[1] = {1'b0,layer_3_2[1743:1736]} - {1'b0, layer_2_2[1743:1736]};
      btm_2[2] = {1'b0,layer_3_2[1751:1744]} - {1'b0, layer_2_2[1751:1744]};
    end
    'd218: begin
      top_0[0] = {1'b0,layer_1_0[1743:1736]} - {1'b0, layer_0_0[1743:1736]};
      top_0[1] = {1'b0,layer_1_0[1751:1744]} - {1'b0, layer_0_0[1751:1744]};
      top_0[2] = {1'b0,layer_1_0[1759:1752]} - {1'b0, layer_0_0[1759:1752]};
      top_1[0] = {1'b0,layer_1_1[1743:1736]} - {1'b0, layer_0_1[1743:1736]};
      top_1[1] = {1'b0,layer_1_1[1751:1744]} - {1'b0, layer_0_1[1751:1744]};
      top_1[2] = {1'b0,layer_1_1[1759:1752]} - {1'b0, layer_0_1[1759:1752]};
      top_2[0] = {1'b0,layer_1_2[1743:1736]} - {1'b0, layer_0_2[1743:1736]};
      top_2[1] = {1'b0,layer_1_2[1751:1744]} - {1'b0, layer_0_2[1751:1744]};
      top_2[2] = {1'b0,layer_1_2[1759:1752]} - {1'b0, layer_0_2[1759:1752]};
      mid_0[0] = {1'b0,layer_2_0[1743:1736]} - {1'b0, layer_1_0[1743:1736]};
      mid_0[1] = {1'b0,layer_2_0[1751:1744]} - {1'b0, layer_1_0[1751:1744]};
      mid_0[2] = {1'b0,layer_2_0[1759:1752]} - {1'b0, layer_1_0[1759:1752]};
      mid_1[0] = {1'b0,layer_2_1[1743:1736]} - {1'b0, layer_1_1[1743:1736]};
      mid_1[1] = {1'b0,layer_2_1[1751:1744]} - {1'b0, layer_1_1[1751:1744]};
      mid_1[2] = {1'b0,layer_2_1[1759:1752]} - {1'b0, layer_1_1[1759:1752]};
      mid_2[0] = {1'b0,layer_2_2[1743:1736]} - {1'b0, layer_1_2[1743:1736]};
      mid_2[1] = {1'b0,layer_2_2[1751:1744]} - {1'b0, layer_1_2[1751:1744]};
      mid_2[2] = {1'b0,layer_2_2[1759:1752]} - {1'b0, layer_1_2[1759:1752]};
      btm_0[0] = {1'b0,layer_3_0[1743:1736]} - {1'b0, layer_2_0[1743:1736]};
      btm_0[1] = {1'b0,layer_3_0[1751:1744]} - {1'b0, layer_2_0[1751:1744]};
      btm_0[2] = {1'b0,layer_3_0[1759:1752]} - {1'b0, layer_2_0[1759:1752]};
      btm_1[0] = {1'b0,layer_3_1[1743:1736]} - {1'b0, layer_2_1[1743:1736]};
      btm_1[1] = {1'b0,layer_3_1[1751:1744]} - {1'b0, layer_2_1[1751:1744]};
      btm_1[2] = {1'b0,layer_3_1[1759:1752]} - {1'b0, layer_2_1[1759:1752]};
      btm_2[0] = {1'b0,layer_3_2[1743:1736]} - {1'b0, layer_2_2[1743:1736]};
      btm_2[1] = {1'b0,layer_3_2[1751:1744]} - {1'b0, layer_2_2[1751:1744]};
      btm_2[2] = {1'b0,layer_3_2[1759:1752]} - {1'b0, layer_2_2[1759:1752]};
    end
    'd219: begin
      top_0[0] = {1'b0,layer_1_0[1751:1744]} - {1'b0, layer_0_0[1751:1744]};
      top_0[1] = {1'b0,layer_1_0[1759:1752]} - {1'b0, layer_0_0[1759:1752]};
      top_0[2] = {1'b0,layer_1_0[1767:1760]} - {1'b0, layer_0_0[1767:1760]};
      top_1[0] = {1'b0,layer_1_1[1751:1744]} - {1'b0, layer_0_1[1751:1744]};
      top_1[1] = {1'b0,layer_1_1[1759:1752]} - {1'b0, layer_0_1[1759:1752]};
      top_1[2] = {1'b0,layer_1_1[1767:1760]} - {1'b0, layer_0_1[1767:1760]};
      top_2[0] = {1'b0,layer_1_2[1751:1744]} - {1'b0, layer_0_2[1751:1744]};
      top_2[1] = {1'b0,layer_1_2[1759:1752]} - {1'b0, layer_0_2[1759:1752]};
      top_2[2] = {1'b0,layer_1_2[1767:1760]} - {1'b0, layer_0_2[1767:1760]};
      mid_0[0] = {1'b0,layer_2_0[1751:1744]} - {1'b0, layer_1_0[1751:1744]};
      mid_0[1] = {1'b0,layer_2_0[1759:1752]} - {1'b0, layer_1_0[1759:1752]};
      mid_0[2] = {1'b0,layer_2_0[1767:1760]} - {1'b0, layer_1_0[1767:1760]};
      mid_1[0] = {1'b0,layer_2_1[1751:1744]} - {1'b0, layer_1_1[1751:1744]};
      mid_1[1] = {1'b0,layer_2_1[1759:1752]} - {1'b0, layer_1_1[1759:1752]};
      mid_1[2] = {1'b0,layer_2_1[1767:1760]} - {1'b0, layer_1_1[1767:1760]};
      mid_2[0] = {1'b0,layer_2_2[1751:1744]} - {1'b0, layer_1_2[1751:1744]};
      mid_2[1] = {1'b0,layer_2_2[1759:1752]} - {1'b0, layer_1_2[1759:1752]};
      mid_2[2] = {1'b0,layer_2_2[1767:1760]} - {1'b0, layer_1_2[1767:1760]};
      btm_0[0] = {1'b0,layer_3_0[1751:1744]} - {1'b0, layer_2_0[1751:1744]};
      btm_0[1] = {1'b0,layer_3_0[1759:1752]} - {1'b0, layer_2_0[1759:1752]};
      btm_0[2] = {1'b0,layer_3_0[1767:1760]} - {1'b0, layer_2_0[1767:1760]};
      btm_1[0] = {1'b0,layer_3_1[1751:1744]} - {1'b0, layer_2_1[1751:1744]};
      btm_1[1] = {1'b0,layer_3_1[1759:1752]} - {1'b0, layer_2_1[1759:1752]};
      btm_1[2] = {1'b0,layer_3_1[1767:1760]} - {1'b0, layer_2_1[1767:1760]};
      btm_2[0] = {1'b0,layer_3_2[1751:1744]} - {1'b0, layer_2_2[1751:1744]};
      btm_2[1] = {1'b0,layer_3_2[1759:1752]} - {1'b0, layer_2_2[1759:1752]};
      btm_2[2] = {1'b0,layer_3_2[1767:1760]} - {1'b0, layer_2_2[1767:1760]};
    end
    'd220: begin
      top_0[0] = {1'b0,layer_1_0[1759:1752]} - {1'b0, layer_0_0[1759:1752]};
      top_0[1] = {1'b0,layer_1_0[1767:1760]} - {1'b0, layer_0_0[1767:1760]};
      top_0[2] = {1'b0,layer_1_0[1775:1768]} - {1'b0, layer_0_0[1775:1768]};
      top_1[0] = {1'b0,layer_1_1[1759:1752]} - {1'b0, layer_0_1[1759:1752]};
      top_1[1] = {1'b0,layer_1_1[1767:1760]} - {1'b0, layer_0_1[1767:1760]};
      top_1[2] = {1'b0,layer_1_1[1775:1768]} - {1'b0, layer_0_1[1775:1768]};
      top_2[0] = {1'b0,layer_1_2[1759:1752]} - {1'b0, layer_0_2[1759:1752]};
      top_2[1] = {1'b0,layer_1_2[1767:1760]} - {1'b0, layer_0_2[1767:1760]};
      top_2[2] = {1'b0,layer_1_2[1775:1768]} - {1'b0, layer_0_2[1775:1768]};
      mid_0[0] = {1'b0,layer_2_0[1759:1752]} - {1'b0, layer_1_0[1759:1752]};
      mid_0[1] = {1'b0,layer_2_0[1767:1760]} - {1'b0, layer_1_0[1767:1760]};
      mid_0[2] = {1'b0,layer_2_0[1775:1768]} - {1'b0, layer_1_0[1775:1768]};
      mid_1[0] = {1'b0,layer_2_1[1759:1752]} - {1'b0, layer_1_1[1759:1752]};
      mid_1[1] = {1'b0,layer_2_1[1767:1760]} - {1'b0, layer_1_1[1767:1760]};
      mid_1[2] = {1'b0,layer_2_1[1775:1768]} - {1'b0, layer_1_1[1775:1768]};
      mid_2[0] = {1'b0,layer_2_2[1759:1752]} - {1'b0, layer_1_2[1759:1752]};
      mid_2[1] = {1'b0,layer_2_2[1767:1760]} - {1'b0, layer_1_2[1767:1760]};
      mid_2[2] = {1'b0,layer_2_2[1775:1768]} - {1'b0, layer_1_2[1775:1768]};
      btm_0[0] = {1'b0,layer_3_0[1759:1752]} - {1'b0, layer_2_0[1759:1752]};
      btm_0[1] = {1'b0,layer_3_0[1767:1760]} - {1'b0, layer_2_0[1767:1760]};
      btm_0[2] = {1'b0,layer_3_0[1775:1768]} - {1'b0, layer_2_0[1775:1768]};
      btm_1[0] = {1'b0,layer_3_1[1759:1752]} - {1'b0, layer_2_1[1759:1752]};
      btm_1[1] = {1'b0,layer_3_1[1767:1760]} - {1'b0, layer_2_1[1767:1760]};
      btm_1[2] = {1'b0,layer_3_1[1775:1768]} - {1'b0, layer_2_1[1775:1768]};
      btm_2[0] = {1'b0,layer_3_2[1759:1752]} - {1'b0, layer_2_2[1759:1752]};
      btm_2[1] = {1'b0,layer_3_2[1767:1760]} - {1'b0, layer_2_2[1767:1760]};
      btm_2[2] = {1'b0,layer_3_2[1775:1768]} - {1'b0, layer_2_2[1775:1768]};
    end
    'd221: begin
      top_0[0] = {1'b0,layer_1_0[1767:1760]} - {1'b0, layer_0_0[1767:1760]};
      top_0[1] = {1'b0,layer_1_0[1775:1768]} - {1'b0, layer_0_0[1775:1768]};
      top_0[2] = {1'b0,layer_1_0[1783:1776]} - {1'b0, layer_0_0[1783:1776]};
      top_1[0] = {1'b0,layer_1_1[1767:1760]} - {1'b0, layer_0_1[1767:1760]};
      top_1[1] = {1'b0,layer_1_1[1775:1768]} - {1'b0, layer_0_1[1775:1768]};
      top_1[2] = {1'b0,layer_1_1[1783:1776]} - {1'b0, layer_0_1[1783:1776]};
      top_2[0] = {1'b0,layer_1_2[1767:1760]} - {1'b0, layer_0_2[1767:1760]};
      top_2[1] = {1'b0,layer_1_2[1775:1768]} - {1'b0, layer_0_2[1775:1768]};
      top_2[2] = {1'b0,layer_1_2[1783:1776]} - {1'b0, layer_0_2[1783:1776]};
      mid_0[0] = {1'b0,layer_2_0[1767:1760]} - {1'b0, layer_1_0[1767:1760]};
      mid_0[1] = {1'b0,layer_2_0[1775:1768]} - {1'b0, layer_1_0[1775:1768]};
      mid_0[2] = {1'b0,layer_2_0[1783:1776]} - {1'b0, layer_1_0[1783:1776]};
      mid_1[0] = {1'b0,layer_2_1[1767:1760]} - {1'b0, layer_1_1[1767:1760]};
      mid_1[1] = {1'b0,layer_2_1[1775:1768]} - {1'b0, layer_1_1[1775:1768]};
      mid_1[2] = {1'b0,layer_2_1[1783:1776]} - {1'b0, layer_1_1[1783:1776]};
      mid_2[0] = {1'b0,layer_2_2[1767:1760]} - {1'b0, layer_1_2[1767:1760]};
      mid_2[1] = {1'b0,layer_2_2[1775:1768]} - {1'b0, layer_1_2[1775:1768]};
      mid_2[2] = {1'b0,layer_2_2[1783:1776]} - {1'b0, layer_1_2[1783:1776]};
      btm_0[0] = {1'b0,layer_3_0[1767:1760]} - {1'b0, layer_2_0[1767:1760]};
      btm_0[1] = {1'b0,layer_3_0[1775:1768]} - {1'b0, layer_2_0[1775:1768]};
      btm_0[2] = {1'b0,layer_3_0[1783:1776]} - {1'b0, layer_2_0[1783:1776]};
      btm_1[0] = {1'b0,layer_3_1[1767:1760]} - {1'b0, layer_2_1[1767:1760]};
      btm_1[1] = {1'b0,layer_3_1[1775:1768]} - {1'b0, layer_2_1[1775:1768]};
      btm_1[2] = {1'b0,layer_3_1[1783:1776]} - {1'b0, layer_2_1[1783:1776]};
      btm_2[0] = {1'b0,layer_3_2[1767:1760]} - {1'b0, layer_2_2[1767:1760]};
      btm_2[1] = {1'b0,layer_3_2[1775:1768]} - {1'b0, layer_2_2[1775:1768]};
      btm_2[2] = {1'b0,layer_3_2[1783:1776]} - {1'b0, layer_2_2[1783:1776]};
    end
    'd222: begin
      top_0[0] = {1'b0,layer_1_0[1775:1768]} - {1'b0, layer_0_0[1775:1768]};
      top_0[1] = {1'b0,layer_1_0[1783:1776]} - {1'b0, layer_0_0[1783:1776]};
      top_0[2] = {1'b0,layer_1_0[1791:1784]} - {1'b0, layer_0_0[1791:1784]};
      top_1[0] = {1'b0,layer_1_1[1775:1768]} - {1'b0, layer_0_1[1775:1768]};
      top_1[1] = {1'b0,layer_1_1[1783:1776]} - {1'b0, layer_0_1[1783:1776]};
      top_1[2] = {1'b0,layer_1_1[1791:1784]} - {1'b0, layer_0_1[1791:1784]};
      top_2[0] = {1'b0,layer_1_2[1775:1768]} - {1'b0, layer_0_2[1775:1768]};
      top_2[1] = {1'b0,layer_1_2[1783:1776]} - {1'b0, layer_0_2[1783:1776]};
      top_2[2] = {1'b0,layer_1_2[1791:1784]} - {1'b0, layer_0_2[1791:1784]};
      mid_0[0] = {1'b0,layer_2_0[1775:1768]} - {1'b0, layer_1_0[1775:1768]};
      mid_0[1] = {1'b0,layer_2_0[1783:1776]} - {1'b0, layer_1_0[1783:1776]};
      mid_0[2] = {1'b0,layer_2_0[1791:1784]} - {1'b0, layer_1_0[1791:1784]};
      mid_1[0] = {1'b0,layer_2_1[1775:1768]} - {1'b0, layer_1_1[1775:1768]};
      mid_1[1] = {1'b0,layer_2_1[1783:1776]} - {1'b0, layer_1_1[1783:1776]};
      mid_1[2] = {1'b0,layer_2_1[1791:1784]} - {1'b0, layer_1_1[1791:1784]};
      mid_2[0] = {1'b0,layer_2_2[1775:1768]} - {1'b0, layer_1_2[1775:1768]};
      mid_2[1] = {1'b0,layer_2_2[1783:1776]} - {1'b0, layer_1_2[1783:1776]};
      mid_2[2] = {1'b0,layer_2_2[1791:1784]} - {1'b0, layer_1_2[1791:1784]};
      btm_0[0] = {1'b0,layer_3_0[1775:1768]} - {1'b0, layer_2_0[1775:1768]};
      btm_0[1] = {1'b0,layer_3_0[1783:1776]} - {1'b0, layer_2_0[1783:1776]};
      btm_0[2] = {1'b0,layer_3_0[1791:1784]} - {1'b0, layer_2_0[1791:1784]};
      btm_1[0] = {1'b0,layer_3_1[1775:1768]} - {1'b0, layer_2_1[1775:1768]};
      btm_1[1] = {1'b0,layer_3_1[1783:1776]} - {1'b0, layer_2_1[1783:1776]};
      btm_1[2] = {1'b0,layer_3_1[1791:1784]} - {1'b0, layer_2_1[1791:1784]};
      btm_2[0] = {1'b0,layer_3_2[1775:1768]} - {1'b0, layer_2_2[1775:1768]};
      btm_2[1] = {1'b0,layer_3_2[1783:1776]} - {1'b0, layer_2_2[1783:1776]};
      btm_2[2] = {1'b0,layer_3_2[1791:1784]} - {1'b0, layer_2_2[1791:1784]};
    end
    'd223: begin
      top_0[0] = {1'b0,layer_1_0[1783:1776]} - {1'b0, layer_0_0[1783:1776]};
      top_0[1] = {1'b0,layer_1_0[1791:1784]} - {1'b0, layer_0_0[1791:1784]};
      top_0[2] = {1'b0,layer_1_0[1799:1792]} - {1'b0, layer_0_0[1799:1792]};
      top_1[0] = {1'b0,layer_1_1[1783:1776]} - {1'b0, layer_0_1[1783:1776]};
      top_1[1] = {1'b0,layer_1_1[1791:1784]} - {1'b0, layer_0_1[1791:1784]};
      top_1[2] = {1'b0,layer_1_1[1799:1792]} - {1'b0, layer_0_1[1799:1792]};
      top_2[0] = {1'b0,layer_1_2[1783:1776]} - {1'b0, layer_0_2[1783:1776]};
      top_2[1] = {1'b0,layer_1_2[1791:1784]} - {1'b0, layer_0_2[1791:1784]};
      top_2[2] = {1'b0,layer_1_2[1799:1792]} - {1'b0, layer_0_2[1799:1792]};
      mid_0[0] = {1'b0,layer_2_0[1783:1776]} - {1'b0, layer_1_0[1783:1776]};
      mid_0[1] = {1'b0,layer_2_0[1791:1784]} - {1'b0, layer_1_0[1791:1784]};
      mid_0[2] = {1'b0,layer_2_0[1799:1792]} - {1'b0, layer_1_0[1799:1792]};
      mid_1[0] = {1'b0,layer_2_1[1783:1776]} - {1'b0, layer_1_1[1783:1776]};
      mid_1[1] = {1'b0,layer_2_1[1791:1784]} - {1'b0, layer_1_1[1791:1784]};
      mid_1[2] = {1'b0,layer_2_1[1799:1792]} - {1'b0, layer_1_1[1799:1792]};
      mid_2[0] = {1'b0,layer_2_2[1783:1776]} - {1'b0, layer_1_2[1783:1776]};
      mid_2[1] = {1'b0,layer_2_2[1791:1784]} - {1'b0, layer_1_2[1791:1784]};
      mid_2[2] = {1'b0,layer_2_2[1799:1792]} - {1'b0, layer_1_2[1799:1792]};
      btm_0[0] = {1'b0,layer_3_0[1783:1776]} - {1'b0, layer_2_0[1783:1776]};
      btm_0[1] = {1'b0,layer_3_0[1791:1784]} - {1'b0, layer_2_0[1791:1784]};
      btm_0[2] = {1'b0,layer_3_0[1799:1792]} - {1'b0, layer_2_0[1799:1792]};
      btm_1[0] = {1'b0,layer_3_1[1783:1776]} - {1'b0, layer_2_1[1783:1776]};
      btm_1[1] = {1'b0,layer_3_1[1791:1784]} - {1'b0, layer_2_1[1791:1784]};
      btm_1[2] = {1'b0,layer_3_1[1799:1792]} - {1'b0, layer_2_1[1799:1792]};
      btm_2[0] = {1'b0,layer_3_2[1783:1776]} - {1'b0, layer_2_2[1783:1776]};
      btm_2[1] = {1'b0,layer_3_2[1791:1784]} - {1'b0, layer_2_2[1791:1784]};
      btm_2[2] = {1'b0,layer_3_2[1799:1792]} - {1'b0, layer_2_2[1799:1792]};
    end
    'd224: begin
      top_0[0] = {1'b0,layer_1_0[1791:1784]} - {1'b0, layer_0_0[1791:1784]};
      top_0[1] = {1'b0,layer_1_0[1799:1792]} - {1'b0, layer_0_0[1799:1792]};
      top_0[2] = {1'b0,layer_1_0[1807:1800]} - {1'b0, layer_0_0[1807:1800]};
      top_1[0] = {1'b0,layer_1_1[1791:1784]} - {1'b0, layer_0_1[1791:1784]};
      top_1[1] = {1'b0,layer_1_1[1799:1792]} - {1'b0, layer_0_1[1799:1792]};
      top_1[2] = {1'b0,layer_1_1[1807:1800]} - {1'b0, layer_0_1[1807:1800]};
      top_2[0] = {1'b0,layer_1_2[1791:1784]} - {1'b0, layer_0_2[1791:1784]};
      top_2[1] = {1'b0,layer_1_2[1799:1792]} - {1'b0, layer_0_2[1799:1792]};
      top_2[2] = {1'b0,layer_1_2[1807:1800]} - {1'b0, layer_0_2[1807:1800]};
      mid_0[0] = {1'b0,layer_2_0[1791:1784]} - {1'b0, layer_1_0[1791:1784]};
      mid_0[1] = {1'b0,layer_2_0[1799:1792]} - {1'b0, layer_1_0[1799:1792]};
      mid_0[2] = {1'b0,layer_2_0[1807:1800]} - {1'b0, layer_1_0[1807:1800]};
      mid_1[0] = {1'b0,layer_2_1[1791:1784]} - {1'b0, layer_1_1[1791:1784]};
      mid_1[1] = {1'b0,layer_2_1[1799:1792]} - {1'b0, layer_1_1[1799:1792]};
      mid_1[2] = {1'b0,layer_2_1[1807:1800]} - {1'b0, layer_1_1[1807:1800]};
      mid_2[0] = {1'b0,layer_2_2[1791:1784]} - {1'b0, layer_1_2[1791:1784]};
      mid_2[1] = {1'b0,layer_2_2[1799:1792]} - {1'b0, layer_1_2[1799:1792]};
      mid_2[2] = {1'b0,layer_2_2[1807:1800]} - {1'b0, layer_1_2[1807:1800]};
      btm_0[0] = {1'b0,layer_3_0[1791:1784]} - {1'b0, layer_2_0[1791:1784]};
      btm_0[1] = {1'b0,layer_3_0[1799:1792]} - {1'b0, layer_2_0[1799:1792]};
      btm_0[2] = {1'b0,layer_3_0[1807:1800]} - {1'b0, layer_2_0[1807:1800]};
      btm_1[0] = {1'b0,layer_3_1[1791:1784]} - {1'b0, layer_2_1[1791:1784]};
      btm_1[1] = {1'b0,layer_3_1[1799:1792]} - {1'b0, layer_2_1[1799:1792]};
      btm_1[2] = {1'b0,layer_3_1[1807:1800]} - {1'b0, layer_2_1[1807:1800]};
      btm_2[0] = {1'b0,layer_3_2[1791:1784]} - {1'b0, layer_2_2[1791:1784]};
      btm_2[1] = {1'b0,layer_3_2[1799:1792]} - {1'b0, layer_2_2[1799:1792]};
      btm_2[2] = {1'b0,layer_3_2[1807:1800]} - {1'b0, layer_2_2[1807:1800]};
    end
    'd225: begin
      top_0[0] = {1'b0,layer_1_0[1799:1792]} - {1'b0, layer_0_0[1799:1792]};
      top_0[1] = {1'b0,layer_1_0[1807:1800]} - {1'b0, layer_0_0[1807:1800]};
      top_0[2] = {1'b0,layer_1_0[1815:1808]} - {1'b0, layer_0_0[1815:1808]};
      top_1[0] = {1'b0,layer_1_1[1799:1792]} - {1'b0, layer_0_1[1799:1792]};
      top_1[1] = {1'b0,layer_1_1[1807:1800]} - {1'b0, layer_0_1[1807:1800]};
      top_1[2] = {1'b0,layer_1_1[1815:1808]} - {1'b0, layer_0_1[1815:1808]};
      top_2[0] = {1'b0,layer_1_2[1799:1792]} - {1'b0, layer_0_2[1799:1792]};
      top_2[1] = {1'b0,layer_1_2[1807:1800]} - {1'b0, layer_0_2[1807:1800]};
      top_2[2] = {1'b0,layer_1_2[1815:1808]} - {1'b0, layer_0_2[1815:1808]};
      mid_0[0] = {1'b0,layer_2_0[1799:1792]} - {1'b0, layer_1_0[1799:1792]};
      mid_0[1] = {1'b0,layer_2_0[1807:1800]} - {1'b0, layer_1_0[1807:1800]};
      mid_0[2] = {1'b0,layer_2_0[1815:1808]} - {1'b0, layer_1_0[1815:1808]};
      mid_1[0] = {1'b0,layer_2_1[1799:1792]} - {1'b0, layer_1_1[1799:1792]};
      mid_1[1] = {1'b0,layer_2_1[1807:1800]} - {1'b0, layer_1_1[1807:1800]};
      mid_1[2] = {1'b0,layer_2_1[1815:1808]} - {1'b0, layer_1_1[1815:1808]};
      mid_2[0] = {1'b0,layer_2_2[1799:1792]} - {1'b0, layer_1_2[1799:1792]};
      mid_2[1] = {1'b0,layer_2_2[1807:1800]} - {1'b0, layer_1_2[1807:1800]};
      mid_2[2] = {1'b0,layer_2_2[1815:1808]} - {1'b0, layer_1_2[1815:1808]};
      btm_0[0] = {1'b0,layer_3_0[1799:1792]} - {1'b0, layer_2_0[1799:1792]};
      btm_0[1] = {1'b0,layer_3_0[1807:1800]} - {1'b0, layer_2_0[1807:1800]};
      btm_0[2] = {1'b0,layer_3_0[1815:1808]} - {1'b0, layer_2_0[1815:1808]};
      btm_1[0] = {1'b0,layer_3_1[1799:1792]} - {1'b0, layer_2_1[1799:1792]};
      btm_1[1] = {1'b0,layer_3_1[1807:1800]} - {1'b0, layer_2_1[1807:1800]};
      btm_1[2] = {1'b0,layer_3_1[1815:1808]} - {1'b0, layer_2_1[1815:1808]};
      btm_2[0] = {1'b0,layer_3_2[1799:1792]} - {1'b0, layer_2_2[1799:1792]};
      btm_2[1] = {1'b0,layer_3_2[1807:1800]} - {1'b0, layer_2_2[1807:1800]};
      btm_2[2] = {1'b0,layer_3_2[1815:1808]} - {1'b0, layer_2_2[1815:1808]};
    end
    'd226: begin
      top_0[0] = {1'b0,layer_1_0[1807:1800]} - {1'b0, layer_0_0[1807:1800]};
      top_0[1] = {1'b0,layer_1_0[1815:1808]} - {1'b0, layer_0_0[1815:1808]};
      top_0[2] = {1'b0,layer_1_0[1823:1816]} - {1'b0, layer_0_0[1823:1816]};
      top_1[0] = {1'b0,layer_1_1[1807:1800]} - {1'b0, layer_0_1[1807:1800]};
      top_1[1] = {1'b0,layer_1_1[1815:1808]} - {1'b0, layer_0_1[1815:1808]};
      top_1[2] = {1'b0,layer_1_1[1823:1816]} - {1'b0, layer_0_1[1823:1816]};
      top_2[0] = {1'b0,layer_1_2[1807:1800]} - {1'b0, layer_0_2[1807:1800]};
      top_2[1] = {1'b0,layer_1_2[1815:1808]} - {1'b0, layer_0_2[1815:1808]};
      top_2[2] = {1'b0,layer_1_2[1823:1816]} - {1'b0, layer_0_2[1823:1816]};
      mid_0[0] = {1'b0,layer_2_0[1807:1800]} - {1'b0, layer_1_0[1807:1800]};
      mid_0[1] = {1'b0,layer_2_0[1815:1808]} - {1'b0, layer_1_0[1815:1808]};
      mid_0[2] = {1'b0,layer_2_0[1823:1816]} - {1'b0, layer_1_0[1823:1816]};
      mid_1[0] = {1'b0,layer_2_1[1807:1800]} - {1'b0, layer_1_1[1807:1800]};
      mid_1[1] = {1'b0,layer_2_1[1815:1808]} - {1'b0, layer_1_1[1815:1808]};
      mid_1[2] = {1'b0,layer_2_1[1823:1816]} - {1'b0, layer_1_1[1823:1816]};
      mid_2[0] = {1'b0,layer_2_2[1807:1800]} - {1'b0, layer_1_2[1807:1800]};
      mid_2[1] = {1'b0,layer_2_2[1815:1808]} - {1'b0, layer_1_2[1815:1808]};
      mid_2[2] = {1'b0,layer_2_2[1823:1816]} - {1'b0, layer_1_2[1823:1816]};
      btm_0[0] = {1'b0,layer_3_0[1807:1800]} - {1'b0, layer_2_0[1807:1800]};
      btm_0[1] = {1'b0,layer_3_0[1815:1808]} - {1'b0, layer_2_0[1815:1808]};
      btm_0[2] = {1'b0,layer_3_0[1823:1816]} - {1'b0, layer_2_0[1823:1816]};
      btm_1[0] = {1'b0,layer_3_1[1807:1800]} - {1'b0, layer_2_1[1807:1800]};
      btm_1[1] = {1'b0,layer_3_1[1815:1808]} - {1'b0, layer_2_1[1815:1808]};
      btm_1[2] = {1'b0,layer_3_1[1823:1816]} - {1'b0, layer_2_1[1823:1816]};
      btm_2[0] = {1'b0,layer_3_2[1807:1800]} - {1'b0, layer_2_2[1807:1800]};
      btm_2[1] = {1'b0,layer_3_2[1815:1808]} - {1'b0, layer_2_2[1815:1808]};
      btm_2[2] = {1'b0,layer_3_2[1823:1816]} - {1'b0, layer_2_2[1823:1816]};
    end
    'd227: begin
      top_0[0] = {1'b0,layer_1_0[1815:1808]} - {1'b0, layer_0_0[1815:1808]};
      top_0[1] = {1'b0,layer_1_0[1823:1816]} - {1'b0, layer_0_0[1823:1816]};
      top_0[2] = {1'b0,layer_1_0[1831:1824]} - {1'b0, layer_0_0[1831:1824]};
      top_1[0] = {1'b0,layer_1_1[1815:1808]} - {1'b0, layer_0_1[1815:1808]};
      top_1[1] = {1'b0,layer_1_1[1823:1816]} - {1'b0, layer_0_1[1823:1816]};
      top_1[2] = {1'b0,layer_1_1[1831:1824]} - {1'b0, layer_0_1[1831:1824]};
      top_2[0] = {1'b0,layer_1_2[1815:1808]} - {1'b0, layer_0_2[1815:1808]};
      top_2[1] = {1'b0,layer_1_2[1823:1816]} - {1'b0, layer_0_2[1823:1816]};
      top_2[2] = {1'b0,layer_1_2[1831:1824]} - {1'b0, layer_0_2[1831:1824]};
      mid_0[0] = {1'b0,layer_2_0[1815:1808]} - {1'b0, layer_1_0[1815:1808]};
      mid_0[1] = {1'b0,layer_2_0[1823:1816]} - {1'b0, layer_1_0[1823:1816]};
      mid_0[2] = {1'b0,layer_2_0[1831:1824]} - {1'b0, layer_1_0[1831:1824]};
      mid_1[0] = {1'b0,layer_2_1[1815:1808]} - {1'b0, layer_1_1[1815:1808]};
      mid_1[1] = {1'b0,layer_2_1[1823:1816]} - {1'b0, layer_1_1[1823:1816]};
      mid_1[2] = {1'b0,layer_2_1[1831:1824]} - {1'b0, layer_1_1[1831:1824]};
      mid_2[0] = {1'b0,layer_2_2[1815:1808]} - {1'b0, layer_1_2[1815:1808]};
      mid_2[1] = {1'b0,layer_2_2[1823:1816]} - {1'b0, layer_1_2[1823:1816]};
      mid_2[2] = {1'b0,layer_2_2[1831:1824]} - {1'b0, layer_1_2[1831:1824]};
      btm_0[0] = {1'b0,layer_3_0[1815:1808]} - {1'b0, layer_2_0[1815:1808]};
      btm_0[1] = {1'b0,layer_3_0[1823:1816]} - {1'b0, layer_2_0[1823:1816]};
      btm_0[2] = {1'b0,layer_3_0[1831:1824]} - {1'b0, layer_2_0[1831:1824]};
      btm_1[0] = {1'b0,layer_3_1[1815:1808]} - {1'b0, layer_2_1[1815:1808]};
      btm_1[1] = {1'b0,layer_3_1[1823:1816]} - {1'b0, layer_2_1[1823:1816]};
      btm_1[2] = {1'b0,layer_3_1[1831:1824]} - {1'b0, layer_2_1[1831:1824]};
      btm_2[0] = {1'b0,layer_3_2[1815:1808]} - {1'b0, layer_2_2[1815:1808]};
      btm_2[1] = {1'b0,layer_3_2[1823:1816]} - {1'b0, layer_2_2[1823:1816]};
      btm_2[2] = {1'b0,layer_3_2[1831:1824]} - {1'b0, layer_2_2[1831:1824]};
    end
    'd228: begin
      top_0[0] = {1'b0,layer_1_0[1823:1816]} - {1'b0, layer_0_0[1823:1816]};
      top_0[1] = {1'b0,layer_1_0[1831:1824]} - {1'b0, layer_0_0[1831:1824]};
      top_0[2] = {1'b0,layer_1_0[1839:1832]} - {1'b0, layer_0_0[1839:1832]};
      top_1[0] = {1'b0,layer_1_1[1823:1816]} - {1'b0, layer_0_1[1823:1816]};
      top_1[1] = {1'b0,layer_1_1[1831:1824]} - {1'b0, layer_0_1[1831:1824]};
      top_1[2] = {1'b0,layer_1_1[1839:1832]} - {1'b0, layer_0_1[1839:1832]};
      top_2[0] = {1'b0,layer_1_2[1823:1816]} - {1'b0, layer_0_2[1823:1816]};
      top_2[1] = {1'b0,layer_1_2[1831:1824]} - {1'b0, layer_0_2[1831:1824]};
      top_2[2] = {1'b0,layer_1_2[1839:1832]} - {1'b0, layer_0_2[1839:1832]};
      mid_0[0] = {1'b0,layer_2_0[1823:1816]} - {1'b0, layer_1_0[1823:1816]};
      mid_0[1] = {1'b0,layer_2_0[1831:1824]} - {1'b0, layer_1_0[1831:1824]};
      mid_0[2] = {1'b0,layer_2_0[1839:1832]} - {1'b0, layer_1_0[1839:1832]};
      mid_1[0] = {1'b0,layer_2_1[1823:1816]} - {1'b0, layer_1_1[1823:1816]};
      mid_1[1] = {1'b0,layer_2_1[1831:1824]} - {1'b0, layer_1_1[1831:1824]};
      mid_1[2] = {1'b0,layer_2_1[1839:1832]} - {1'b0, layer_1_1[1839:1832]};
      mid_2[0] = {1'b0,layer_2_2[1823:1816]} - {1'b0, layer_1_2[1823:1816]};
      mid_2[1] = {1'b0,layer_2_2[1831:1824]} - {1'b0, layer_1_2[1831:1824]};
      mid_2[2] = {1'b0,layer_2_2[1839:1832]} - {1'b0, layer_1_2[1839:1832]};
      btm_0[0] = {1'b0,layer_3_0[1823:1816]} - {1'b0, layer_2_0[1823:1816]};
      btm_0[1] = {1'b0,layer_3_0[1831:1824]} - {1'b0, layer_2_0[1831:1824]};
      btm_0[2] = {1'b0,layer_3_0[1839:1832]} - {1'b0, layer_2_0[1839:1832]};
      btm_1[0] = {1'b0,layer_3_1[1823:1816]} - {1'b0, layer_2_1[1823:1816]};
      btm_1[1] = {1'b0,layer_3_1[1831:1824]} - {1'b0, layer_2_1[1831:1824]};
      btm_1[2] = {1'b0,layer_3_1[1839:1832]} - {1'b0, layer_2_1[1839:1832]};
      btm_2[0] = {1'b0,layer_3_2[1823:1816]} - {1'b0, layer_2_2[1823:1816]};
      btm_2[1] = {1'b0,layer_3_2[1831:1824]} - {1'b0, layer_2_2[1831:1824]};
      btm_2[2] = {1'b0,layer_3_2[1839:1832]} - {1'b0, layer_2_2[1839:1832]};
    end
    'd229: begin
      top_0[0] = {1'b0,layer_1_0[1831:1824]} - {1'b0, layer_0_0[1831:1824]};
      top_0[1] = {1'b0,layer_1_0[1839:1832]} - {1'b0, layer_0_0[1839:1832]};
      top_0[2] = {1'b0,layer_1_0[1847:1840]} - {1'b0, layer_0_0[1847:1840]};
      top_1[0] = {1'b0,layer_1_1[1831:1824]} - {1'b0, layer_0_1[1831:1824]};
      top_1[1] = {1'b0,layer_1_1[1839:1832]} - {1'b0, layer_0_1[1839:1832]};
      top_1[2] = {1'b0,layer_1_1[1847:1840]} - {1'b0, layer_0_1[1847:1840]};
      top_2[0] = {1'b0,layer_1_2[1831:1824]} - {1'b0, layer_0_2[1831:1824]};
      top_2[1] = {1'b0,layer_1_2[1839:1832]} - {1'b0, layer_0_2[1839:1832]};
      top_2[2] = {1'b0,layer_1_2[1847:1840]} - {1'b0, layer_0_2[1847:1840]};
      mid_0[0] = {1'b0,layer_2_0[1831:1824]} - {1'b0, layer_1_0[1831:1824]};
      mid_0[1] = {1'b0,layer_2_0[1839:1832]} - {1'b0, layer_1_0[1839:1832]};
      mid_0[2] = {1'b0,layer_2_0[1847:1840]} - {1'b0, layer_1_0[1847:1840]};
      mid_1[0] = {1'b0,layer_2_1[1831:1824]} - {1'b0, layer_1_1[1831:1824]};
      mid_1[1] = {1'b0,layer_2_1[1839:1832]} - {1'b0, layer_1_1[1839:1832]};
      mid_1[2] = {1'b0,layer_2_1[1847:1840]} - {1'b0, layer_1_1[1847:1840]};
      mid_2[0] = {1'b0,layer_2_2[1831:1824]} - {1'b0, layer_1_2[1831:1824]};
      mid_2[1] = {1'b0,layer_2_2[1839:1832]} - {1'b0, layer_1_2[1839:1832]};
      mid_2[2] = {1'b0,layer_2_2[1847:1840]} - {1'b0, layer_1_2[1847:1840]};
      btm_0[0] = {1'b0,layer_3_0[1831:1824]} - {1'b0, layer_2_0[1831:1824]};
      btm_0[1] = {1'b0,layer_3_0[1839:1832]} - {1'b0, layer_2_0[1839:1832]};
      btm_0[2] = {1'b0,layer_3_0[1847:1840]} - {1'b0, layer_2_0[1847:1840]};
      btm_1[0] = {1'b0,layer_3_1[1831:1824]} - {1'b0, layer_2_1[1831:1824]};
      btm_1[1] = {1'b0,layer_3_1[1839:1832]} - {1'b0, layer_2_1[1839:1832]};
      btm_1[2] = {1'b0,layer_3_1[1847:1840]} - {1'b0, layer_2_1[1847:1840]};
      btm_2[0] = {1'b0,layer_3_2[1831:1824]} - {1'b0, layer_2_2[1831:1824]};
      btm_2[1] = {1'b0,layer_3_2[1839:1832]} - {1'b0, layer_2_2[1839:1832]};
      btm_2[2] = {1'b0,layer_3_2[1847:1840]} - {1'b0, layer_2_2[1847:1840]};
    end
    'd230: begin
      top_0[0] = {1'b0,layer_1_0[1839:1832]} - {1'b0, layer_0_0[1839:1832]};
      top_0[1] = {1'b0,layer_1_0[1847:1840]} - {1'b0, layer_0_0[1847:1840]};
      top_0[2] = {1'b0,layer_1_0[1855:1848]} - {1'b0, layer_0_0[1855:1848]};
      top_1[0] = {1'b0,layer_1_1[1839:1832]} - {1'b0, layer_0_1[1839:1832]};
      top_1[1] = {1'b0,layer_1_1[1847:1840]} - {1'b0, layer_0_1[1847:1840]};
      top_1[2] = {1'b0,layer_1_1[1855:1848]} - {1'b0, layer_0_1[1855:1848]};
      top_2[0] = {1'b0,layer_1_2[1839:1832]} - {1'b0, layer_0_2[1839:1832]};
      top_2[1] = {1'b0,layer_1_2[1847:1840]} - {1'b0, layer_0_2[1847:1840]};
      top_2[2] = {1'b0,layer_1_2[1855:1848]} - {1'b0, layer_0_2[1855:1848]};
      mid_0[0] = {1'b0,layer_2_0[1839:1832]} - {1'b0, layer_1_0[1839:1832]};
      mid_0[1] = {1'b0,layer_2_0[1847:1840]} - {1'b0, layer_1_0[1847:1840]};
      mid_0[2] = {1'b0,layer_2_0[1855:1848]} - {1'b0, layer_1_0[1855:1848]};
      mid_1[0] = {1'b0,layer_2_1[1839:1832]} - {1'b0, layer_1_1[1839:1832]};
      mid_1[1] = {1'b0,layer_2_1[1847:1840]} - {1'b0, layer_1_1[1847:1840]};
      mid_1[2] = {1'b0,layer_2_1[1855:1848]} - {1'b0, layer_1_1[1855:1848]};
      mid_2[0] = {1'b0,layer_2_2[1839:1832]} - {1'b0, layer_1_2[1839:1832]};
      mid_2[1] = {1'b0,layer_2_2[1847:1840]} - {1'b0, layer_1_2[1847:1840]};
      mid_2[2] = {1'b0,layer_2_2[1855:1848]} - {1'b0, layer_1_2[1855:1848]};
      btm_0[0] = {1'b0,layer_3_0[1839:1832]} - {1'b0, layer_2_0[1839:1832]};
      btm_0[1] = {1'b0,layer_3_0[1847:1840]} - {1'b0, layer_2_0[1847:1840]};
      btm_0[2] = {1'b0,layer_3_0[1855:1848]} - {1'b0, layer_2_0[1855:1848]};
      btm_1[0] = {1'b0,layer_3_1[1839:1832]} - {1'b0, layer_2_1[1839:1832]};
      btm_1[1] = {1'b0,layer_3_1[1847:1840]} - {1'b0, layer_2_1[1847:1840]};
      btm_1[2] = {1'b0,layer_3_1[1855:1848]} - {1'b0, layer_2_1[1855:1848]};
      btm_2[0] = {1'b0,layer_3_2[1839:1832]} - {1'b0, layer_2_2[1839:1832]};
      btm_2[1] = {1'b0,layer_3_2[1847:1840]} - {1'b0, layer_2_2[1847:1840]};
      btm_2[2] = {1'b0,layer_3_2[1855:1848]} - {1'b0, layer_2_2[1855:1848]};
    end
    'd231: begin
      top_0[0] = {1'b0,layer_1_0[1847:1840]} - {1'b0, layer_0_0[1847:1840]};
      top_0[1] = {1'b0,layer_1_0[1855:1848]} - {1'b0, layer_0_0[1855:1848]};
      top_0[2] = {1'b0,layer_1_0[1863:1856]} - {1'b0, layer_0_0[1863:1856]};
      top_1[0] = {1'b0,layer_1_1[1847:1840]} - {1'b0, layer_0_1[1847:1840]};
      top_1[1] = {1'b0,layer_1_1[1855:1848]} - {1'b0, layer_0_1[1855:1848]};
      top_1[2] = {1'b0,layer_1_1[1863:1856]} - {1'b0, layer_0_1[1863:1856]};
      top_2[0] = {1'b0,layer_1_2[1847:1840]} - {1'b0, layer_0_2[1847:1840]};
      top_2[1] = {1'b0,layer_1_2[1855:1848]} - {1'b0, layer_0_2[1855:1848]};
      top_2[2] = {1'b0,layer_1_2[1863:1856]} - {1'b0, layer_0_2[1863:1856]};
      mid_0[0] = {1'b0,layer_2_0[1847:1840]} - {1'b0, layer_1_0[1847:1840]};
      mid_0[1] = {1'b0,layer_2_0[1855:1848]} - {1'b0, layer_1_0[1855:1848]};
      mid_0[2] = {1'b0,layer_2_0[1863:1856]} - {1'b0, layer_1_0[1863:1856]};
      mid_1[0] = {1'b0,layer_2_1[1847:1840]} - {1'b0, layer_1_1[1847:1840]};
      mid_1[1] = {1'b0,layer_2_1[1855:1848]} - {1'b0, layer_1_1[1855:1848]};
      mid_1[2] = {1'b0,layer_2_1[1863:1856]} - {1'b0, layer_1_1[1863:1856]};
      mid_2[0] = {1'b0,layer_2_2[1847:1840]} - {1'b0, layer_1_2[1847:1840]};
      mid_2[1] = {1'b0,layer_2_2[1855:1848]} - {1'b0, layer_1_2[1855:1848]};
      mid_2[2] = {1'b0,layer_2_2[1863:1856]} - {1'b0, layer_1_2[1863:1856]};
      btm_0[0] = {1'b0,layer_3_0[1847:1840]} - {1'b0, layer_2_0[1847:1840]};
      btm_0[1] = {1'b0,layer_3_0[1855:1848]} - {1'b0, layer_2_0[1855:1848]};
      btm_0[2] = {1'b0,layer_3_0[1863:1856]} - {1'b0, layer_2_0[1863:1856]};
      btm_1[0] = {1'b0,layer_3_1[1847:1840]} - {1'b0, layer_2_1[1847:1840]};
      btm_1[1] = {1'b0,layer_3_1[1855:1848]} - {1'b0, layer_2_1[1855:1848]};
      btm_1[2] = {1'b0,layer_3_1[1863:1856]} - {1'b0, layer_2_1[1863:1856]};
      btm_2[0] = {1'b0,layer_3_2[1847:1840]} - {1'b0, layer_2_2[1847:1840]};
      btm_2[1] = {1'b0,layer_3_2[1855:1848]} - {1'b0, layer_2_2[1855:1848]};
      btm_2[2] = {1'b0,layer_3_2[1863:1856]} - {1'b0, layer_2_2[1863:1856]};
    end
    'd232: begin
      top_0[0] = {1'b0,layer_1_0[1855:1848]} - {1'b0, layer_0_0[1855:1848]};
      top_0[1] = {1'b0,layer_1_0[1863:1856]} - {1'b0, layer_0_0[1863:1856]};
      top_0[2] = {1'b0,layer_1_0[1871:1864]} - {1'b0, layer_0_0[1871:1864]};
      top_1[0] = {1'b0,layer_1_1[1855:1848]} - {1'b0, layer_0_1[1855:1848]};
      top_1[1] = {1'b0,layer_1_1[1863:1856]} - {1'b0, layer_0_1[1863:1856]};
      top_1[2] = {1'b0,layer_1_1[1871:1864]} - {1'b0, layer_0_1[1871:1864]};
      top_2[0] = {1'b0,layer_1_2[1855:1848]} - {1'b0, layer_0_2[1855:1848]};
      top_2[1] = {1'b0,layer_1_2[1863:1856]} - {1'b0, layer_0_2[1863:1856]};
      top_2[2] = {1'b0,layer_1_2[1871:1864]} - {1'b0, layer_0_2[1871:1864]};
      mid_0[0] = {1'b0,layer_2_0[1855:1848]} - {1'b0, layer_1_0[1855:1848]};
      mid_0[1] = {1'b0,layer_2_0[1863:1856]} - {1'b0, layer_1_0[1863:1856]};
      mid_0[2] = {1'b0,layer_2_0[1871:1864]} - {1'b0, layer_1_0[1871:1864]};
      mid_1[0] = {1'b0,layer_2_1[1855:1848]} - {1'b0, layer_1_1[1855:1848]};
      mid_1[1] = {1'b0,layer_2_1[1863:1856]} - {1'b0, layer_1_1[1863:1856]};
      mid_1[2] = {1'b0,layer_2_1[1871:1864]} - {1'b0, layer_1_1[1871:1864]};
      mid_2[0] = {1'b0,layer_2_2[1855:1848]} - {1'b0, layer_1_2[1855:1848]};
      mid_2[1] = {1'b0,layer_2_2[1863:1856]} - {1'b0, layer_1_2[1863:1856]};
      mid_2[2] = {1'b0,layer_2_2[1871:1864]} - {1'b0, layer_1_2[1871:1864]};
      btm_0[0] = {1'b0,layer_3_0[1855:1848]} - {1'b0, layer_2_0[1855:1848]};
      btm_0[1] = {1'b0,layer_3_0[1863:1856]} - {1'b0, layer_2_0[1863:1856]};
      btm_0[2] = {1'b0,layer_3_0[1871:1864]} - {1'b0, layer_2_0[1871:1864]};
      btm_1[0] = {1'b0,layer_3_1[1855:1848]} - {1'b0, layer_2_1[1855:1848]};
      btm_1[1] = {1'b0,layer_3_1[1863:1856]} - {1'b0, layer_2_1[1863:1856]};
      btm_1[2] = {1'b0,layer_3_1[1871:1864]} - {1'b0, layer_2_1[1871:1864]};
      btm_2[0] = {1'b0,layer_3_2[1855:1848]} - {1'b0, layer_2_2[1855:1848]};
      btm_2[1] = {1'b0,layer_3_2[1863:1856]} - {1'b0, layer_2_2[1863:1856]};
      btm_2[2] = {1'b0,layer_3_2[1871:1864]} - {1'b0, layer_2_2[1871:1864]};
    end
    'd233: begin
      top_0[0] = {1'b0,layer_1_0[1863:1856]} - {1'b0, layer_0_0[1863:1856]};
      top_0[1] = {1'b0,layer_1_0[1871:1864]} - {1'b0, layer_0_0[1871:1864]};
      top_0[2] = {1'b0,layer_1_0[1879:1872]} - {1'b0, layer_0_0[1879:1872]};
      top_1[0] = {1'b0,layer_1_1[1863:1856]} - {1'b0, layer_0_1[1863:1856]};
      top_1[1] = {1'b0,layer_1_1[1871:1864]} - {1'b0, layer_0_1[1871:1864]};
      top_1[2] = {1'b0,layer_1_1[1879:1872]} - {1'b0, layer_0_1[1879:1872]};
      top_2[0] = {1'b0,layer_1_2[1863:1856]} - {1'b0, layer_0_2[1863:1856]};
      top_2[1] = {1'b0,layer_1_2[1871:1864]} - {1'b0, layer_0_2[1871:1864]};
      top_2[2] = {1'b0,layer_1_2[1879:1872]} - {1'b0, layer_0_2[1879:1872]};
      mid_0[0] = {1'b0,layer_2_0[1863:1856]} - {1'b0, layer_1_0[1863:1856]};
      mid_0[1] = {1'b0,layer_2_0[1871:1864]} - {1'b0, layer_1_0[1871:1864]};
      mid_0[2] = {1'b0,layer_2_0[1879:1872]} - {1'b0, layer_1_0[1879:1872]};
      mid_1[0] = {1'b0,layer_2_1[1863:1856]} - {1'b0, layer_1_1[1863:1856]};
      mid_1[1] = {1'b0,layer_2_1[1871:1864]} - {1'b0, layer_1_1[1871:1864]};
      mid_1[2] = {1'b0,layer_2_1[1879:1872]} - {1'b0, layer_1_1[1879:1872]};
      mid_2[0] = {1'b0,layer_2_2[1863:1856]} - {1'b0, layer_1_2[1863:1856]};
      mid_2[1] = {1'b0,layer_2_2[1871:1864]} - {1'b0, layer_1_2[1871:1864]};
      mid_2[2] = {1'b0,layer_2_2[1879:1872]} - {1'b0, layer_1_2[1879:1872]};
      btm_0[0] = {1'b0,layer_3_0[1863:1856]} - {1'b0, layer_2_0[1863:1856]};
      btm_0[1] = {1'b0,layer_3_0[1871:1864]} - {1'b0, layer_2_0[1871:1864]};
      btm_0[2] = {1'b0,layer_3_0[1879:1872]} - {1'b0, layer_2_0[1879:1872]};
      btm_1[0] = {1'b0,layer_3_1[1863:1856]} - {1'b0, layer_2_1[1863:1856]};
      btm_1[1] = {1'b0,layer_3_1[1871:1864]} - {1'b0, layer_2_1[1871:1864]};
      btm_1[2] = {1'b0,layer_3_1[1879:1872]} - {1'b0, layer_2_1[1879:1872]};
      btm_2[0] = {1'b0,layer_3_2[1863:1856]} - {1'b0, layer_2_2[1863:1856]};
      btm_2[1] = {1'b0,layer_3_2[1871:1864]} - {1'b0, layer_2_2[1871:1864]};
      btm_2[2] = {1'b0,layer_3_2[1879:1872]} - {1'b0, layer_2_2[1879:1872]};
    end
    'd234: begin
      top_0[0] = {1'b0,layer_1_0[1871:1864]} - {1'b0, layer_0_0[1871:1864]};
      top_0[1] = {1'b0,layer_1_0[1879:1872]} - {1'b0, layer_0_0[1879:1872]};
      top_0[2] = {1'b0,layer_1_0[1887:1880]} - {1'b0, layer_0_0[1887:1880]};
      top_1[0] = {1'b0,layer_1_1[1871:1864]} - {1'b0, layer_0_1[1871:1864]};
      top_1[1] = {1'b0,layer_1_1[1879:1872]} - {1'b0, layer_0_1[1879:1872]};
      top_1[2] = {1'b0,layer_1_1[1887:1880]} - {1'b0, layer_0_1[1887:1880]};
      top_2[0] = {1'b0,layer_1_2[1871:1864]} - {1'b0, layer_0_2[1871:1864]};
      top_2[1] = {1'b0,layer_1_2[1879:1872]} - {1'b0, layer_0_2[1879:1872]};
      top_2[2] = {1'b0,layer_1_2[1887:1880]} - {1'b0, layer_0_2[1887:1880]};
      mid_0[0] = {1'b0,layer_2_0[1871:1864]} - {1'b0, layer_1_0[1871:1864]};
      mid_0[1] = {1'b0,layer_2_0[1879:1872]} - {1'b0, layer_1_0[1879:1872]};
      mid_0[2] = {1'b0,layer_2_0[1887:1880]} - {1'b0, layer_1_0[1887:1880]};
      mid_1[0] = {1'b0,layer_2_1[1871:1864]} - {1'b0, layer_1_1[1871:1864]};
      mid_1[1] = {1'b0,layer_2_1[1879:1872]} - {1'b0, layer_1_1[1879:1872]};
      mid_1[2] = {1'b0,layer_2_1[1887:1880]} - {1'b0, layer_1_1[1887:1880]};
      mid_2[0] = {1'b0,layer_2_2[1871:1864]} - {1'b0, layer_1_2[1871:1864]};
      mid_2[1] = {1'b0,layer_2_2[1879:1872]} - {1'b0, layer_1_2[1879:1872]};
      mid_2[2] = {1'b0,layer_2_2[1887:1880]} - {1'b0, layer_1_2[1887:1880]};
      btm_0[0] = {1'b0,layer_3_0[1871:1864]} - {1'b0, layer_2_0[1871:1864]};
      btm_0[1] = {1'b0,layer_3_0[1879:1872]} - {1'b0, layer_2_0[1879:1872]};
      btm_0[2] = {1'b0,layer_3_0[1887:1880]} - {1'b0, layer_2_0[1887:1880]};
      btm_1[0] = {1'b0,layer_3_1[1871:1864]} - {1'b0, layer_2_1[1871:1864]};
      btm_1[1] = {1'b0,layer_3_1[1879:1872]} - {1'b0, layer_2_1[1879:1872]};
      btm_1[2] = {1'b0,layer_3_1[1887:1880]} - {1'b0, layer_2_1[1887:1880]};
      btm_2[0] = {1'b0,layer_3_2[1871:1864]} - {1'b0, layer_2_2[1871:1864]};
      btm_2[1] = {1'b0,layer_3_2[1879:1872]} - {1'b0, layer_2_2[1879:1872]};
      btm_2[2] = {1'b0,layer_3_2[1887:1880]} - {1'b0, layer_2_2[1887:1880]};
    end
    'd235: begin
      top_0[0] = {1'b0,layer_1_0[1879:1872]} - {1'b0, layer_0_0[1879:1872]};
      top_0[1] = {1'b0,layer_1_0[1887:1880]} - {1'b0, layer_0_0[1887:1880]};
      top_0[2] = {1'b0,layer_1_0[1895:1888]} - {1'b0, layer_0_0[1895:1888]};
      top_1[0] = {1'b0,layer_1_1[1879:1872]} - {1'b0, layer_0_1[1879:1872]};
      top_1[1] = {1'b0,layer_1_1[1887:1880]} - {1'b0, layer_0_1[1887:1880]};
      top_1[2] = {1'b0,layer_1_1[1895:1888]} - {1'b0, layer_0_1[1895:1888]};
      top_2[0] = {1'b0,layer_1_2[1879:1872]} - {1'b0, layer_0_2[1879:1872]};
      top_2[1] = {1'b0,layer_1_2[1887:1880]} - {1'b0, layer_0_2[1887:1880]};
      top_2[2] = {1'b0,layer_1_2[1895:1888]} - {1'b0, layer_0_2[1895:1888]};
      mid_0[0] = {1'b0,layer_2_0[1879:1872]} - {1'b0, layer_1_0[1879:1872]};
      mid_0[1] = {1'b0,layer_2_0[1887:1880]} - {1'b0, layer_1_0[1887:1880]};
      mid_0[2] = {1'b0,layer_2_0[1895:1888]} - {1'b0, layer_1_0[1895:1888]};
      mid_1[0] = {1'b0,layer_2_1[1879:1872]} - {1'b0, layer_1_1[1879:1872]};
      mid_1[1] = {1'b0,layer_2_1[1887:1880]} - {1'b0, layer_1_1[1887:1880]};
      mid_1[2] = {1'b0,layer_2_1[1895:1888]} - {1'b0, layer_1_1[1895:1888]};
      mid_2[0] = {1'b0,layer_2_2[1879:1872]} - {1'b0, layer_1_2[1879:1872]};
      mid_2[1] = {1'b0,layer_2_2[1887:1880]} - {1'b0, layer_1_2[1887:1880]};
      mid_2[2] = {1'b0,layer_2_2[1895:1888]} - {1'b0, layer_1_2[1895:1888]};
      btm_0[0] = {1'b0,layer_3_0[1879:1872]} - {1'b0, layer_2_0[1879:1872]};
      btm_0[1] = {1'b0,layer_3_0[1887:1880]} - {1'b0, layer_2_0[1887:1880]};
      btm_0[2] = {1'b0,layer_3_0[1895:1888]} - {1'b0, layer_2_0[1895:1888]};
      btm_1[0] = {1'b0,layer_3_1[1879:1872]} - {1'b0, layer_2_1[1879:1872]};
      btm_1[1] = {1'b0,layer_3_1[1887:1880]} - {1'b0, layer_2_1[1887:1880]};
      btm_1[2] = {1'b0,layer_3_1[1895:1888]} - {1'b0, layer_2_1[1895:1888]};
      btm_2[0] = {1'b0,layer_3_2[1879:1872]} - {1'b0, layer_2_2[1879:1872]};
      btm_2[1] = {1'b0,layer_3_2[1887:1880]} - {1'b0, layer_2_2[1887:1880]};
      btm_2[2] = {1'b0,layer_3_2[1895:1888]} - {1'b0, layer_2_2[1895:1888]};
    end
    'd236: begin
      top_0[0] = {1'b0,layer_1_0[1887:1880]} - {1'b0, layer_0_0[1887:1880]};
      top_0[1] = {1'b0,layer_1_0[1895:1888]} - {1'b0, layer_0_0[1895:1888]};
      top_0[2] = {1'b0,layer_1_0[1903:1896]} - {1'b0, layer_0_0[1903:1896]};
      top_1[0] = {1'b0,layer_1_1[1887:1880]} - {1'b0, layer_0_1[1887:1880]};
      top_1[1] = {1'b0,layer_1_1[1895:1888]} - {1'b0, layer_0_1[1895:1888]};
      top_1[2] = {1'b0,layer_1_1[1903:1896]} - {1'b0, layer_0_1[1903:1896]};
      top_2[0] = {1'b0,layer_1_2[1887:1880]} - {1'b0, layer_0_2[1887:1880]};
      top_2[1] = {1'b0,layer_1_2[1895:1888]} - {1'b0, layer_0_2[1895:1888]};
      top_2[2] = {1'b0,layer_1_2[1903:1896]} - {1'b0, layer_0_2[1903:1896]};
      mid_0[0] = {1'b0,layer_2_0[1887:1880]} - {1'b0, layer_1_0[1887:1880]};
      mid_0[1] = {1'b0,layer_2_0[1895:1888]} - {1'b0, layer_1_0[1895:1888]};
      mid_0[2] = {1'b0,layer_2_0[1903:1896]} - {1'b0, layer_1_0[1903:1896]};
      mid_1[0] = {1'b0,layer_2_1[1887:1880]} - {1'b0, layer_1_1[1887:1880]};
      mid_1[1] = {1'b0,layer_2_1[1895:1888]} - {1'b0, layer_1_1[1895:1888]};
      mid_1[2] = {1'b0,layer_2_1[1903:1896]} - {1'b0, layer_1_1[1903:1896]};
      mid_2[0] = {1'b0,layer_2_2[1887:1880]} - {1'b0, layer_1_2[1887:1880]};
      mid_2[1] = {1'b0,layer_2_2[1895:1888]} - {1'b0, layer_1_2[1895:1888]};
      mid_2[2] = {1'b0,layer_2_2[1903:1896]} - {1'b0, layer_1_2[1903:1896]};
      btm_0[0] = {1'b0,layer_3_0[1887:1880]} - {1'b0, layer_2_0[1887:1880]};
      btm_0[1] = {1'b0,layer_3_0[1895:1888]} - {1'b0, layer_2_0[1895:1888]};
      btm_0[2] = {1'b0,layer_3_0[1903:1896]} - {1'b0, layer_2_0[1903:1896]};
      btm_1[0] = {1'b0,layer_3_1[1887:1880]} - {1'b0, layer_2_1[1887:1880]};
      btm_1[1] = {1'b0,layer_3_1[1895:1888]} - {1'b0, layer_2_1[1895:1888]};
      btm_1[2] = {1'b0,layer_3_1[1903:1896]} - {1'b0, layer_2_1[1903:1896]};
      btm_2[0] = {1'b0,layer_3_2[1887:1880]} - {1'b0, layer_2_2[1887:1880]};
      btm_2[1] = {1'b0,layer_3_2[1895:1888]} - {1'b0, layer_2_2[1895:1888]};
      btm_2[2] = {1'b0,layer_3_2[1903:1896]} - {1'b0, layer_2_2[1903:1896]};
    end
    'd237: begin
      top_0[0] = {1'b0,layer_1_0[1895:1888]} - {1'b0, layer_0_0[1895:1888]};
      top_0[1] = {1'b0,layer_1_0[1903:1896]} - {1'b0, layer_0_0[1903:1896]};
      top_0[2] = {1'b0,layer_1_0[1911:1904]} - {1'b0, layer_0_0[1911:1904]};
      top_1[0] = {1'b0,layer_1_1[1895:1888]} - {1'b0, layer_0_1[1895:1888]};
      top_1[1] = {1'b0,layer_1_1[1903:1896]} - {1'b0, layer_0_1[1903:1896]};
      top_1[2] = {1'b0,layer_1_1[1911:1904]} - {1'b0, layer_0_1[1911:1904]};
      top_2[0] = {1'b0,layer_1_2[1895:1888]} - {1'b0, layer_0_2[1895:1888]};
      top_2[1] = {1'b0,layer_1_2[1903:1896]} - {1'b0, layer_0_2[1903:1896]};
      top_2[2] = {1'b0,layer_1_2[1911:1904]} - {1'b0, layer_0_2[1911:1904]};
      mid_0[0] = {1'b0,layer_2_0[1895:1888]} - {1'b0, layer_1_0[1895:1888]};
      mid_0[1] = {1'b0,layer_2_0[1903:1896]} - {1'b0, layer_1_0[1903:1896]};
      mid_0[2] = {1'b0,layer_2_0[1911:1904]} - {1'b0, layer_1_0[1911:1904]};
      mid_1[0] = {1'b0,layer_2_1[1895:1888]} - {1'b0, layer_1_1[1895:1888]};
      mid_1[1] = {1'b0,layer_2_1[1903:1896]} - {1'b0, layer_1_1[1903:1896]};
      mid_1[2] = {1'b0,layer_2_1[1911:1904]} - {1'b0, layer_1_1[1911:1904]};
      mid_2[0] = {1'b0,layer_2_2[1895:1888]} - {1'b0, layer_1_2[1895:1888]};
      mid_2[1] = {1'b0,layer_2_2[1903:1896]} - {1'b0, layer_1_2[1903:1896]};
      mid_2[2] = {1'b0,layer_2_2[1911:1904]} - {1'b0, layer_1_2[1911:1904]};
      btm_0[0] = {1'b0,layer_3_0[1895:1888]} - {1'b0, layer_2_0[1895:1888]};
      btm_0[1] = {1'b0,layer_3_0[1903:1896]} - {1'b0, layer_2_0[1903:1896]};
      btm_0[2] = {1'b0,layer_3_0[1911:1904]} - {1'b0, layer_2_0[1911:1904]};
      btm_1[0] = {1'b0,layer_3_1[1895:1888]} - {1'b0, layer_2_1[1895:1888]};
      btm_1[1] = {1'b0,layer_3_1[1903:1896]} - {1'b0, layer_2_1[1903:1896]};
      btm_1[2] = {1'b0,layer_3_1[1911:1904]} - {1'b0, layer_2_1[1911:1904]};
      btm_2[0] = {1'b0,layer_3_2[1895:1888]} - {1'b0, layer_2_2[1895:1888]};
      btm_2[1] = {1'b0,layer_3_2[1903:1896]} - {1'b0, layer_2_2[1903:1896]};
      btm_2[2] = {1'b0,layer_3_2[1911:1904]} - {1'b0, layer_2_2[1911:1904]};
    end
    'd238: begin
      top_0[0] = {1'b0,layer_1_0[1903:1896]} - {1'b0, layer_0_0[1903:1896]};
      top_0[1] = {1'b0,layer_1_0[1911:1904]} - {1'b0, layer_0_0[1911:1904]};
      top_0[2] = {1'b0,layer_1_0[1919:1912]} - {1'b0, layer_0_0[1919:1912]};
      top_1[0] = {1'b0,layer_1_1[1903:1896]} - {1'b0, layer_0_1[1903:1896]};
      top_1[1] = {1'b0,layer_1_1[1911:1904]} - {1'b0, layer_0_1[1911:1904]};
      top_1[2] = {1'b0,layer_1_1[1919:1912]} - {1'b0, layer_0_1[1919:1912]};
      top_2[0] = {1'b0,layer_1_2[1903:1896]} - {1'b0, layer_0_2[1903:1896]};
      top_2[1] = {1'b0,layer_1_2[1911:1904]} - {1'b0, layer_0_2[1911:1904]};
      top_2[2] = {1'b0,layer_1_2[1919:1912]} - {1'b0, layer_0_2[1919:1912]};
      mid_0[0] = {1'b0,layer_2_0[1903:1896]} - {1'b0, layer_1_0[1903:1896]};
      mid_0[1] = {1'b0,layer_2_0[1911:1904]} - {1'b0, layer_1_0[1911:1904]};
      mid_0[2] = {1'b0,layer_2_0[1919:1912]} - {1'b0, layer_1_0[1919:1912]};
      mid_1[0] = {1'b0,layer_2_1[1903:1896]} - {1'b0, layer_1_1[1903:1896]};
      mid_1[1] = {1'b0,layer_2_1[1911:1904]} - {1'b0, layer_1_1[1911:1904]};
      mid_1[2] = {1'b0,layer_2_1[1919:1912]} - {1'b0, layer_1_1[1919:1912]};
      mid_2[0] = {1'b0,layer_2_2[1903:1896]} - {1'b0, layer_1_2[1903:1896]};
      mid_2[1] = {1'b0,layer_2_2[1911:1904]} - {1'b0, layer_1_2[1911:1904]};
      mid_2[2] = {1'b0,layer_2_2[1919:1912]} - {1'b0, layer_1_2[1919:1912]};
      btm_0[0] = {1'b0,layer_3_0[1903:1896]} - {1'b0, layer_2_0[1903:1896]};
      btm_0[1] = {1'b0,layer_3_0[1911:1904]} - {1'b0, layer_2_0[1911:1904]};
      btm_0[2] = {1'b0,layer_3_0[1919:1912]} - {1'b0, layer_2_0[1919:1912]};
      btm_1[0] = {1'b0,layer_3_1[1903:1896]} - {1'b0, layer_2_1[1903:1896]};
      btm_1[1] = {1'b0,layer_3_1[1911:1904]} - {1'b0, layer_2_1[1911:1904]};
      btm_1[2] = {1'b0,layer_3_1[1919:1912]} - {1'b0, layer_2_1[1919:1912]};
      btm_2[0] = {1'b0,layer_3_2[1903:1896]} - {1'b0, layer_2_2[1903:1896]};
      btm_2[1] = {1'b0,layer_3_2[1911:1904]} - {1'b0, layer_2_2[1911:1904]};
      btm_2[2] = {1'b0,layer_3_2[1919:1912]} - {1'b0, layer_2_2[1919:1912]};
    end
    'd239: begin
      top_0[0] = {1'b0,layer_1_0[1911:1904]} - {1'b0, layer_0_0[1911:1904]};
      top_0[1] = {1'b0,layer_1_0[1919:1912]} - {1'b0, layer_0_0[1919:1912]};
      top_0[2] = {1'b0,layer_1_0[1927:1920]} - {1'b0, layer_0_0[1927:1920]};
      top_1[0] = {1'b0,layer_1_1[1911:1904]} - {1'b0, layer_0_1[1911:1904]};
      top_1[1] = {1'b0,layer_1_1[1919:1912]} - {1'b0, layer_0_1[1919:1912]};
      top_1[2] = {1'b0,layer_1_1[1927:1920]} - {1'b0, layer_0_1[1927:1920]};
      top_2[0] = {1'b0,layer_1_2[1911:1904]} - {1'b0, layer_0_2[1911:1904]};
      top_2[1] = {1'b0,layer_1_2[1919:1912]} - {1'b0, layer_0_2[1919:1912]};
      top_2[2] = {1'b0,layer_1_2[1927:1920]} - {1'b0, layer_0_2[1927:1920]};
      mid_0[0] = {1'b0,layer_2_0[1911:1904]} - {1'b0, layer_1_0[1911:1904]};
      mid_0[1] = {1'b0,layer_2_0[1919:1912]} - {1'b0, layer_1_0[1919:1912]};
      mid_0[2] = {1'b0,layer_2_0[1927:1920]} - {1'b0, layer_1_0[1927:1920]};
      mid_1[0] = {1'b0,layer_2_1[1911:1904]} - {1'b0, layer_1_1[1911:1904]};
      mid_1[1] = {1'b0,layer_2_1[1919:1912]} - {1'b0, layer_1_1[1919:1912]};
      mid_1[2] = {1'b0,layer_2_1[1927:1920]} - {1'b0, layer_1_1[1927:1920]};
      mid_2[0] = {1'b0,layer_2_2[1911:1904]} - {1'b0, layer_1_2[1911:1904]};
      mid_2[1] = {1'b0,layer_2_2[1919:1912]} - {1'b0, layer_1_2[1919:1912]};
      mid_2[2] = {1'b0,layer_2_2[1927:1920]} - {1'b0, layer_1_2[1927:1920]};
      btm_0[0] = {1'b0,layer_3_0[1911:1904]} - {1'b0, layer_2_0[1911:1904]};
      btm_0[1] = {1'b0,layer_3_0[1919:1912]} - {1'b0, layer_2_0[1919:1912]};
      btm_0[2] = {1'b0,layer_3_0[1927:1920]} - {1'b0, layer_2_0[1927:1920]};
      btm_1[0] = {1'b0,layer_3_1[1911:1904]} - {1'b0, layer_2_1[1911:1904]};
      btm_1[1] = {1'b0,layer_3_1[1919:1912]} - {1'b0, layer_2_1[1919:1912]};
      btm_1[2] = {1'b0,layer_3_1[1927:1920]} - {1'b0, layer_2_1[1927:1920]};
      btm_2[0] = {1'b0,layer_3_2[1911:1904]} - {1'b0, layer_2_2[1911:1904]};
      btm_2[1] = {1'b0,layer_3_2[1919:1912]} - {1'b0, layer_2_2[1919:1912]};
      btm_2[2] = {1'b0,layer_3_2[1927:1920]} - {1'b0, layer_2_2[1927:1920]};
    end
    'd240: begin
      top_0[0] = {1'b0,layer_1_0[1919:1912]} - {1'b0, layer_0_0[1919:1912]};
      top_0[1] = {1'b0,layer_1_0[1927:1920]} - {1'b0, layer_0_0[1927:1920]};
      top_0[2] = {1'b0,layer_1_0[1935:1928]} - {1'b0, layer_0_0[1935:1928]};
      top_1[0] = {1'b0,layer_1_1[1919:1912]} - {1'b0, layer_0_1[1919:1912]};
      top_1[1] = {1'b0,layer_1_1[1927:1920]} - {1'b0, layer_0_1[1927:1920]};
      top_1[2] = {1'b0,layer_1_1[1935:1928]} - {1'b0, layer_0_1[1935:1928]};
      top_2[0] = {1'b0,layer_1_2[1919:1912]} - {1'b0, layer_0_2[1919:1912]};
      top_2[1] = {1'b0,layer_1_2[1927:1920]} - {1'b0, layer_0_2[1927:1920]};
      top_2[2] = {1'b0,layer_1_2[1935:1928]} - {1'b0, layer_0_2[1935:1928]};
      mid_0[0] = {1'b0,layer_2_0[1919:1912]} - {1'b0, layer_1_0[1919:1912]};
      mid_0[1] = {1'b0,layer_2_0[1927:1920]} - {1'b0, layer_1_0[1927:1920]};
      mid_0[2] = {1'b0,layer_2_0[1935:1928]} - {1'b0, layer_1_0[1935:1928]};
      mid_1[0] = {1'b0,layer_2_1[1919:1912]} - {1'b0, layer_1_1[1919:1912]};
      mid_1[1] = {1'b0,layer_2_1[1927:1920]} - {1'b0, layer_1_1[1927:1920]};
      mid_1[2] = {1'b0,layer_2_1[1935:1928]} - {1'b0, layer_1_1[1935:1928]};
      mid_2[0] = {1'b0,layer_2_2[1919:1912]} - {1'b0, layer_1_2[1919:1912]};
      mid_2[1] = {1'b0,layer_2_2[1927:1920]} - {1'b0, layer_1_2[1927:1920]};
      mid_2[2] = {1'b0,layer_2_2[1935:1928]} - {1'b0, layer_1_2[1935:1928]};
      btm_0[0] = {1'b0,layer_3_0[1919:1912]} - {1'b0, layer_2_0[1919:1912]};
      btm_0[1] = {1'b0,layer_3_0[1927:1920]} - {1'b0, layer_2_0[1927:1920]};
      btm_0[2] = {1'b0,layer_3_0[1935:1928]} - {1'b0, layer_2_0[1935:1928]};
      btm_1[0] = {1'b0,layer_3_1[1919:1912]} - {1'b0, layer_2_1[1919:1912]};
      btm_1[1] = {1'b0,layer_3_1[1927:1920]} - {1'b0, layer_2_1[1927:1920]};
      btm_1[2] = {1'b0,layer_3_1[1935:1928]} - {1'b0, layer_2_1[1935:1928]};
      btm_2[0] = {1'b0,layer_3_2[1919:1912]} - {1'b0, layer_2_2[1919:1912]};
      btm_2[1] = {1'b0,layer_3_2[1927:1920]} - {1'b0, layer_2_2[1927:1920]};
      btm_2[2] = {1'b0,layer_3_2[1935:1928]} - {1'b0, layer_2_2[1935:1928]};
    end
    'd241: begin
      top_0[0] = {1'b0,layer_1_0[1927:1920]} - {1'b0, layer_0_0[1927:1920]};
      top_0[1] = {1'b0,layer_1_0[1935:1928]} - {1'b0, layer_0_0[1935:1928]};
      top_0[2] = {1'b0,layer_1_0[1943:1936]} - {1'b0, layer_0_0[1943:1936]};
      top_1[0] = {1'b0,layer_1_1[1927:1920]} - {1'b0, layer_0_1[1927:1920]};
      top_1[1] = {1'b0,layer_1_1[1935:1928]} - {1'b0, layer_0_1[1935:1928]};
      top_1[2] = {1'b0,layer_1_1[1943:1936]} - {1'b0, layer_0_1[1943:1936]};
      top_2[0] = {1'b0,layer_1_2[1927:1920]} - {1'b0, layer_0_2[1927:1920]};
      top_2[1] = {1'b0,layer_1_2[1935:1928]} - {1'b0, layer_0_2[1935:1928]};
      top_2[2] = {1'b0,layer_1_2[1943:1936]} - {1'b0, layer_0_2[1943:1936]};
      mid_0[0] = {1'b0,layer_2_0[1927:1920]} - {1'b0, layer_1_0[1927:1920]};
      mid_0[1] = {1'b0,layer_2_0[1935:1928]} - {1'b0, layer_1_0[1935:1928]};
      mid_0[2] = {1'b0,layer_2_0[1943:1936]} - {1'b0, layer_1_0[1943:1936]};
      mid_1[0] = {1'b0,layer_2_1[1927:1920]} - {1'b0, layer_1_1[1927:1920]};
      mid_1[1] = {1'b0,layer_2_1[1935:1928]} - {1'b0, layer_1_1[1935:1928]};
      mid_1[2] = {1'b0,layer_2_1[1943:1936]} - {1'b0, layer_1_1[1943:1936]};
      mid_2[0] = {1'b0,layer_2_2[1927:1920]} - {1'b0, layer_1_2[1927:1920]};
      mid_2[1] = {1'b0,layer_2_2[1935:1928]} - {1'b0, layer_1_2[1935:1928]};
      mid_2[2] = {1'b0,layer_2_2[1943:1936]} - {1'b0, layer_1_2[1943:1936]};
      btm_0[0] = {1'b0,layer_3_0[1927:1920]} - {1'b0, layer_2_0[1927:1920]};
      btm_0[1] = {1'b0,layer_3_0[1935:1928]} - {1'b0, layer_2_0[1935:1928]};
      btm_0[2] = {1'b0,layer_3_0[1943:1936]} - {1'b0, layer_2_0[1943:1936]};
      btm_1[0] = {1'b0,layer_3_1[1927:1920]} - {1'b0, layer_2_1[1927:1920]};
      btm_1[1] = {1'b0,layer_3_1[1935:1928]} - {1'b0, layer_2_1[1935:1928]};
      btm_1[2] = {1'b0,layer_3_1[1943:1936]} - {1'b0, layer_2_1[1943:1936]};
      btm_2[0] = {1'b0,layer_3_2[1927:1920]} - {1'b0, layer_2_2[1927:1920]};
      btm_2[1] = {1'b0,layer_3_2[1935:1928]} - {1'b0, layer_2_2[1935:1928]};
      btm_2[2] = {1'b0,layer_3_2[1943:1936]} - {1'b0, layer_2_2[1943:1936]};
    end
    'd242: begin
      top_0[0] = {1'b0,layer_1_0[1935:1928]} - {1'b0, layer_0_0[1935:1928]};
      top_0[1] = {1'b0,layer_1_0[1943:1936]} - {1'b0, layer_0_0[1943:1936]};
      top_0[2] = {1'b0,layer_1_0[1951:1944]} - {1'b0, layer_0_0[1951:1944]};
      top_1[0] = {1'b0,layer_1_1[1935:1928]} - {1'b0, layer_0_1[1935:1928]};
      top_1[1] = {1'b0,layer_1_1[1943:1936]} - {1'b0, layer_0_1[1943:1936]};
      top_1[2] = {1'b0,layer_1_1[1951:1944]} - {1'b0, layer_0_1[1951:1944]};
      top_2[0] = {1'b0,layer_1_2[1935:1928]} - {1'b0, layer_0_2[1935:1928]};
      top_2[1] = {1'b0,layer_1_2[1943:1936]} - {1'b0, layer_0_2[1943:1936]};
      top_2[2] = {1'b0,layer_1_2[1951:1944]} - {1'b0, layer_0_2[1951:1944]};
      mid_0[0] = {1'b0,layer_2_0[1935:1928]} - {1'b0, layer_1_0[1935:1928]};
      mid_0[1] = {1'b0,layer_2_0[1943:1936]} - {1'b0, layer_1_0[1943:1936]};
      mid_0[2] = {1'b0,layer_2_0[1951:1944]} - {1'b0, layer_1_0[1951:1944]};
      mid_1[0] = {1'b0,layer_2_1[1935:1928]} - {1'b0, layer_1_1[1935:1928]};
      mid_1[1] = {1'b0,layer_2_1[1943:1936]} - {1'b0, layer_1_1[1943:1936]};
      mid_1[2] = {1'b0,layer_2_1[1951:1944]} - {1'b0, layer_1_1[1951:1944]};
      mid_2[0] = {1'b0,layer_2_2[1935:1928]} - {1'b0, layer_1_2[1935:1928]};
      mid_2[1] = {1'b0,layer_2_2[1943:1936]} - {1'b0, layer_1_2[1943:1936]};
      mid_2[2] = {1'b0,layer_2_2[1951:1944]} - {1'b0, layer_1_2[1951:1944]};
      btm_0[0] = {1'b0,layer_3_0[1935:1928]} - {1'b0, layer_2_0[1935:1928]};
      btm_0[1] = {1'b0,layer_3_0[1943:1936]} - {1'b0, layer_2_0[1943:1936]};
      btm_0[2] = {1'b0,layer_3_0[1951:1944]} - {1'b0, layer_2_0[1951:1944]};
      btm_1[0] = {1'b0,layer_3_1[1935:1928]} - {1'b0, layer_2_1[1935:1928]};
      btm_1[1] = {1'b0,layer_3_1[1943:1936]} - {1'b0, layer_2_1[1943:1936]};
      btm_1[2] = {1'b0,layer_3_1[1951:1944]} - {1'b0, layer_2_1[1951:1944]};
      btm_2[0] = {1'b0,layer_3_2[1935:1928]} - {1'b0, layer_2_2[1935:1928]};
      btm_2[1] = {1'b0,layer_3_2[1943:1936]} - {1'b0, layer_2_2[1943:1936]};
      btm_2[2] = {1'b0,layer_3_2[1951:1944]} - {1'b0, layer_2_2[1951:1944]};
    end
    'd243: begin
      top_0[0] = {1'b0,layer_1_0[1943:1936]} - {1'b0, layer_0_0[1943:1936]};
      top_0[1] = {1'b0,layer_1_0[1951:1944]} - {1'b0, layer_0_0[1951:1944]};
      top_0[2] = {1'b0,layer_1_0[1959:1952]} - {1'b0, layer_0_0[1959:1952]};
      top_1[0] = {1'b0,layer_1_1[1943:1936]} - {1'b0, layer_0_1[1943:1936]};
      top_1[1] = {1'b0,layer_1_1[1951:1944]} - {1'b0, layer_0_1[1951:1944]};
      top_1[2] = {1'b0,layer_1_1[1959:1952]} - {1'b0, layer_0_1[1959:1952]};
      top_2[0] = {1'b0,layer_1_2[1943:1936]} - {1'b0, layer_0_2[1943:1936]};
      top_2[1] = {1'b0,layer_1_2[1951:1944]} - {1'b0, layer_0_2[1951:1944]};
      top_2[2] = {1'b0,layer_1_2[1959:1952]} - {1'b0, layer_0_2[1959:1952]};
      mid_0[0] = {1'b0,layer_2_0[1943:1936]} - {1'b0, layer_1_0[1943:1936]};
      mid_0[1] = {1'b0,layer_2_0[1951:1944]} - {1'b0, layer_1_0[1951:1944]};
      mid_0[2] = {1'b0,layer_2_0[1959:1952]} - {1'b0, layer_1_0[1959:1952]};
      mid_1[0] = {1'b0,layer_2_1[1943:1936]} - {1'b0, layer_1_1[1943:1936]};
      mid_1[1] = {1'b0,layer_2_1[1951:1944]} - {1'b0, layer_1_1[1951:1944]};
      mid_1[2] = {1'b0,layer_2_1[1959:1952]} - {1'b0, layer_1_1[1959:1952]};
      mid_2[0] = {1'b0,layer_2_2[1943:1936]} - {1'b0, layer_1_2[1943:1936]};
      mid_2[1] = {1'b0,layer_2_2[1951:1944]} - {1'b0, layer_1_2[1951:1944]};
      mid_2[2] = {1'b0,layer_2_2[1959:1952]} - {1'b0, layer_1_2[1959:1952]};
      btm_0[0] = {1'b0,layer_3_0[1943:1936]} - {1'b0, layer_2_0[1943:1936]};
      btm_0[1] = {1'b0,layer_3_0[1951:1944]} - {1'b0, layer_2_0[1951:1944]};
      btm_0[2] = {1'b0,layer_3_0[1959:1952]} - {1'b0, layer_2_0[1959:1952]};
      btm_1[0] = {1'b0,layer_3_1[1943:1936]} - {1'b0, layer_2_1[1943:1936]};
      btm_1[1] = {1'b0,layer_3_1[1951:1944]} - {1'b0, layer_2_1[1951:1944]};
      btm_1[2] = {1'b0,layer_3_1[1959:1952]} - {1'b0, layer_2_1[1959:1952]};
      btm_2[0] = {1'b0,layer_3_2[1943:1936]} - {1'b0, layer_2_2[1943:1936]};
      btm_2[1] = {1'b0,layer_3_2[1951:1944]} - {1'b0, layer_2_2[1951:1944]};
      btm_2[2] = {1'b0,layer_3_2[1959:1952]} - {1'b0, layer_2_2[1959:1952]};
    end
    'd244: begin
      top_0[0] = {1'b0,layer_1_0[1951:1944]} - {1'b0, layer_0_0[1951:1944]};
      top_0[1] = {1'b0,layer_1_0[1959:1952]} - {1'b0, layer_0_0[1959:1952]};
      top_0[2] = {1'b0,layer_1_0[1967:1960]} - {1'b0, layer_0_0[1967:1960]};
      top_1[0] = {1'b0,layer_1_1[1951:1944]} - {1'b0, layer_0_1[1951:1944]};
      top_1[1] = {1'b0,layer_1_1[1959:1952]} - {1'b0, layer_0_1[1959:1952]};
      top_1[2] = {1'b0,layer_1_1[1967:1960]} - {1'b0, layer_0_1[1967:1960]};
      top_2[0] = {1'b0,layer_1_2[1951:1944]} - {1'b0, layer_0_2[1951:1944]};
      top_2[1] = {1'b0,layer_1_2[1959:1952]} - {1'b0, layer_0_2[1959:1952]};
      top_2[2] = {1'b0,layer_1_2[1967:1960]} - {1'b0, layer_0_2[1967:1960]};
      mid_0[0] = {1'b0,layer_2_0[1951:1944]} - {1'b0, layer_1_0[1951:1944]};
      mid_0[1] = {1'b0,layer_2_0[1959:1952]} - {1'b0, layer_1_0[1959:1952]};
      mid_0[2] = {1'b0,layer_2_0[1967:1960]} - {1'b0, layer_1_0[1967:1960]};
      mid_1[0] = {1'b0,layer_2_1[1951:1944]} - {1'b0, layer_1_1[1951:1944]};
      mid_1[1] = {1'b0,layer_2_1[1959:1952]} - {1'b0, layer_1_1[1959:1952]};
      mid_1[2] = {1'b0,layer_2_1[1967:1960]} - {1'b0, layer_1_1[1967:1960]};
      mid_2[0] = {1'b0,layer_2_2[1951:1944]} - {1'b0, layer_1_2[1951:1944]};
      mid_2[1] = {1'b0,layer_2_2[1959:1952]} - {1'b0, layer_1_2[1959:1952]};
      mid_2[2] = {1'b0,layer_2_2[1967:1960]} - {1'b0, layer_1_2[1967:1960]};
      btm_0[0] = {1'b0,layer_3_0[1951:1944]} - {1'b0, layer_2_0[1951:1944]};
      btm_0[1] = {1'b0,layer_3_0[1959:1952]} - {1'b0, layer_2_0[1959:1952]};
      btm_0[2] = {1'b0,layer_3_0[1967:1960]} - {1'b0, layer_2_0[1967:1960]};
      btm_1[0] = {1'b0,layer_3_1[1951:1944]} - {1'b0, layer_2_1[1951:1944]};
      btm_1[1] = {1'b0,layer_3_1[1959:1952]} - {1'b0, layer_2_1[1959:1952]};
      btm_1[2] = {1'b0,layer_3_1[1967:1960]} - {1'b0, layer_2_1[1967:1960]};
      btm_2[0] = {1'b0,layer_3_2[1951:1944]} - {1'b0, layer_2_2[1951:1944]};
      btm_2[1] = {1'b0,layer_3_2[1959:1952]} - {1'b0, layer_2_2[1959:1952]};
      btm_2[2] = {1'b0,layer_3_2[1967:1960]} - {1'b0, layer_2_2[1967:1960]};
    end
    'd245: begin
      top_0[0] = {1'b0,layer_1_0[1959:1952]} - {1'b0, layer_0_0[1959:1952]};
      top_0[1] = {1'b0,layer_1_0[1967:1960]} - {1'b0, layer_0_0[1967:1960]};
      top_0[2] = {1'b0,layer_1_0[1975:1968]} - {1'b0, layer_0_0[1975:1968]};
      top_1[0] = {1'b0,layer_1_1[1959:1952]} - {1'b0, layer_0_1[1959:1952]};
      top_1[1] = {1'b0,layer_1_1[1967:1960]} - {1'b0, layer_0_1[1967:1960]};
      top_1[2] = {1'b0,layer_1_1[1975:1968]} - {1'b0, layer_0_1[1975:1968]};
      top_2[0] = {1'b0,layer_1_2[1959:1952]} - {1'b0, layer_0_2[1959:1952]};
      top_2[1] = {1'b0,layer_1_2[1967:1960]} - {1'b0, layer_0_2[1967:1960]};
      top_2[2] = {1'b0,layer_1_2[1975:1968]} - {1'b0, layer_0_2[1975:1968]};
      mid_0[0] = {1'b0,layer_2_0[1959:1952]} - {1'b0, layer_1_0[1959:1952]};
      mid_0[1] = {1'b0,layer_2_0[1967:1960]} - {1'b0, layer_1_0[1967:1960]};
      mid_0[2] = {1'b0,layer_2_0[1975:1968]} - {1'b0, layer_1_0[1975:1968]};
      mid_1[0] = {1'b0,layer_2_1[1959:1952]} - {1'b0, layer_1_1[1959:1952]};
      mid_1[1] = {1'b0,layer_2_1[1967:1960]} - {1'b0, layer_1_1[1967:1960]};
      mid_1[2] = {1'b0,layer_2_1[1975:1968]} - {1'b0, layer_1_1[1975:1968]};
      mid_2[0] = {1'b0,layer_2_2[1959:1952]} - {1'b0, layer_1_2[1959:1952]};
      mid_2[1] = {1'b0,layer_2_2[1967:1960]} - {1'b0, layer_1_2[1967:1960]};
      mid_2[2] = {1'b0,layer_2_2[1975:1968]} - {1'b0, layer_1_2[1975:1968]};
      btm_0[0] = {1'b0,layer_3_0[1959:1952]} - {1'b0, layer_2_0[1959:1952]};
      btm_0[1] = {1'b0,layer_3_0[1967:1960]} - {1'b0, layer_2_0[1967:1960]};
      btm_0[2] = {1'b0,layer_3_0[1975:1968]} - {1'b0, layer_2_0[1975:1968]};
      btm_1[0] = {1'b0,layer_3_1[1959:1952]} - {1'b0, layer_2_1[1959:1952]};
      btm_1[1] = {1'b0,layer_3_1[1967:1960]} - {1'b0, layer_2_1[1967:1960]};
      btm_1[2] = {1'b0,layer_3_1[1975:1968]} - {1'b0, layer_2_1[1975:1968]};
      btm_2[0] = {1'b0,layer_3_2[1959:1952]} - {1'b0, layer_2_2[1959:1952]};
      btm_2[1] = {1'b0,layer_3_2[1967:1960]} - {1'b0, layer_2_2[1967:1960]};
      btm_2[2] = {1'b0,layer_3_2[1975:1968]} - {1'b0, layer_2_2[1975:1968]};
    end
    'd246: begin
      top_0[0] = {1'b0,layer_1_0[1967:1960]} - {1'b0, layer_0_0[1967:1960]};
      top_0[1] = {1'b0,layer_1_0[1975:1968]} - {1'b0, layer_0_0[1975:1968]};
      top_0[2] = {1'b0,layer_1_0[1983:1976]} - {1'b0, layer_0_0[1983:1976]};
      top_1[0] = {1'b0,layer_1_1[1967:1960]} - {1'b0, layer_0_1[1967:1960]};
      top_1[1] = {1'b0,layer_1_1[1975:1968]} - {1'b0, layer_0_1[1975:1968]};
      top_1[2] = {1'b0,layer_1_1[1983:1976]} - {1'b0, layer_0_1[1983:1976]};
      top_2[0] = {1'b0,layer_1_2[1967:1960]} - {1'b0, layer_0_2[1967:1960]};
      top_2[1] = {1'b0,layer_1_2[1975:1968]} - {1'b0, layer_0_2[1975:1968]};
      top_2[2] = {1'b0,layer_1_2[1983:1976]} - {1'b0, layer_0_2[1983:1976]};
      mid_0[0] = {1'b0,layer_2_0[1967:1960]} - {1'b0, layer_1_0[1967:1960]};
      mid_0[1] = {1'b0,layer_2_0[1975:1968]} - {1'b0, layer_1_0[1975:1968]};
      mid_0[2] = {1'b0,layer_2_0[1983:1976]} - {1'b0, layer_1_0[1983:1976]};
      mid_1[0] = {1'b0,layer_2_1[1967:1960]} - {1'b0, layer_1_1[1967:1960]};
      mid_1[1] = {1'b0,layer_2_1[1975:1968]} - {1'b0, layer_1_1[1975:1968]};
      mid_1[2] = {1'b0,layer_2_1[1983:1976]} - {1'b0, layer_1_1[1983:1976]};
      mid_2[0] = {1'b0,layer_2_2[1967:1960]} - {1'b0, layer_1_2[1967:1960]};
      mid_2[1] = {1'b0,layer_2_2[1975:1968]} - {1'b0, layer_1_2[1975:1968]};
      mid_2[2] = {1'b0,layer_2_2[1983:1976]} - {1'b0, layer_1_2[1983:1976]};
      btm_0[0] = {1'b0,layer_3_0[1967:1960]} - {1'b0, layer_2_0[1967:1960]};
      btm_0[1] = {1'b0,layer_3_0[1975:1968]} - {1'b0, layer_2_0[1975:1968]};
      btm_0[2] = {1'b0,layer_3_0[1983:1976]} - {1'b0, layer_2_0[1983:1976]};
      btm_1[0] = {1'b0,layer_3_1[1967:1960]} - {1'b0, layer_2_1[1967:1960]};
      btm_1[1] = {1'b0,layer_3_1[1975:1968]} - {1'b0, layer_2_1[1975:1968]};
      btm_1[2] = {1'b0,layer_3_1[1983:1976]} - {1'b0, layer_2_1[1983:1976]};
      btm_2[0] = {1'b0,layer_3_2[1967:1960]} - {1'b0, layer_2_2[1967:1960]};
      btm_2[1] = {1'b0,layer_3_2[1975:1968]} - {1'b0, layer_2_2[1975:1968]};
      btm_2[2] = {1'b0,layer_3_2[1983:1976]} - {1'b0, layer_2_2[1983:1976]};
    end
    'd247: begin
      top_0[0] = {1'b0,layer_1_0[1975:1968]} - {1'b0, layer_0_0[1975:1968]};
      top_0[1] = {1'b0,layer_1_0[1983:1976]} - {1'b0, layer_0_0[1983:1976]};
      top_0[2] = {1'b0,layer_1_0[1991:1984]} - {1'b0, layer_0_0[1991:1984]};
      top_1[0] = {1'b0,layer_1_1[1975:1968]} - {1'b0, layer_0_1[1975:1968]};
      top_1[1] = {1'b0,layer_1_1[1983:1976]} - {1'b0, layer_0_1[1983:1976]};
      top_1[2] = {1'b0,layer_1_1[1991:1984]} - {1'b0, layer_0_1[1991:1984]};
      top_2[0] = {1'b0,layer_1_2[1975:1968]} - {1'b0, layer_0_2[1975:1968]};
      top_2[1] = {1'b0,layer_1_2[1983:1976]} - {1'b0, layer_0_2[1983:1976]};
      top_2[2] = {1'b0,layer_1_2[1991:1984]} - {1'b0, layer_0_2[1991:1984]};
      mid_0[0] = {1'b0,layer_2_0[1975:1968]} - {1'b0, layer_1_0[1975:1968]};
      mid_0[1] = {1'b0,layer_2_0[1983:1976]} - {1'b0, layer_1_0[1983:1976]};
      mid_0[2] = {1'b0,layer_2_0[1991:1984]} - {1'b0, layer_1_0[1991:1984]};
      mid_1[0] = {1'b0,layer_2_1[1975:1968]} - {1'b0, layer_1_1[1975:1968]};
      mid_1[1] = {1'b0,layer_2_1[1983:1976]} - {1'b0, layer_1_1[1983:1976]};
      mid_1[2] = {1'b0,layer_2_1[1991:1984]} - {1'b0, layer_1_1[1991:1984]};
      mid_2[0] = {1'b0,layer_2_2[1975:1968]} - {1'b0, layer_1_2[1975:1968]};
      mid_2[1] = {1'b0,layer_2_2[1983:1976]} - {1'b0, layer_1_2[1983:1976]};
      mid_2[2] = {1'b0,layer_2_2[1991:1984]} - {1'b0, layer_1_2[1991:1984]};
      btm_0[0] = {1'b0,layer_3_0[1975:1968]} - {1'b0, layer_2_0[1975:1968]};
      btm_0[1] = {1'b0,layer_3_0[1983:1976]} - {1'b0, layer_2_0[1983:1976]};
      btm_0[2] = {1'b0,layer_3_0[1991:1984]} - {1'b0, layer_2_0[1991:1984]};
      btm_1[0] = {1'b0,layer_3_1[1975:1968]} - {1'b0, layer_2_1[1975:1968]};
      btm_1[1] = {1'b0,layer_3_1[1983:1976]} - {1'b0, layer_2_1[1983:1976]};
      btm_1[2] = {1'b0,layer_3_1[1991:1984]} - {1'b0, layer_2_1[1991:1984]};
      btm_2[0] = {1'b0,layer_3_2[1975:1968]} - {1'b0, layer_2_2[1975:1968]};
      btm_2[1] = {1'b0,layer_3_2[1983:1976]} - {1'b0, layer_2_2[1983:1976]};
      btm_2[2] = {1'b0,layer_3_2[1991:1984]} - {1'b0, layer_2_2[1991:1984]};
    end
    'd248: begin
      top_0[0] = {1'b0,layer_1_0[1983:1976]} - {1'b0, layer_0_0[1983:1976]};
      top_0[1] = {1'b0,layer_1_0[1991:1984]} - {1'b0, layer_0_0[1991:1984]};
      top_0[2] = {1'b0,layer_1_0[1999:1992]} - {1'b0, layer_0_0[1999:1992]};
      top_1[0] = {1'b0,layer_1_1[1983:1976]} - {1'b0, layer_0_1[1983:1976]};
      top_1[1] = {1'b0,layer_1_1[1991:1984]} - {1'b0, layer_0_1[1991:1984]};
      top_1[2] = {1'b0,layer_1_1[1999:1992]} - {1'b0, layer_0_1[1999:1992]};
      top_2[0] = {1'b0,layer_1_2[1983:1976]} - {1'b0, layer_0_2[1983:1976]};
      top_2[1] = {1'b0,layer_1_2[1991:1984]} - {1'b0, layer_0_2[1991:1984]};
      top_2[2] = {1'b0,layer_1_2[1999:1992]} - {1'b0, layer_0_2[1999:1992]};
      mid_0[0] = {1'b0,layer_2_0[1983:1976]} - {1'b0, layer_1_0[1983:1976]};
      mid_0[1] = {1'b0,layer_2_0[1991:1984]} - {1'b0, layer_1_0[1991:1984]};
      mid_0[2] = {1'b0,layer_2_0[1999:1992]} - {1'b0, layer_1_0[1999:1992]};
      mid_1[0] = {1'b0,layer_2_1[1983:1976]} - {1'b0, layer_1_1[1983:1976]};
      mid_1[1] = {1'b0,layer_2_1[1991:1984]} - {1'b0, layer_1_1[1991:1984]};
      mid_1[2] = {1'b0,layer_2_1[1999:1992]} - {1'b0, layer_1_1[1999:1992]};
      mid_2[0] = {1'b0,layer_2_2[1983:1976]} - {1'b0, layer_1_2[1983:1976]};
      mid_2[1] = {1'b0,layer_2_2[1991:1984]} - {1'b0, layer_1_2[1991:1984]};
      mid_2[2] = {1'b0,layer_2_2[1999:1992]} - {1'b0, layer_1_2[1999:1992]};
      btm_0[0] = {1'b0,layer_3_0[1983:1976]} - {1'b0, layer_2_0[1983:1976]};
      btm_0[1] = {1'b0,layer_3_0[1991:1984]} - {1'b0, layer_2_0[1991:1984]};
      btm_0[2] = {1'b0,layer_3_0[1999:1992]} - {1'b0, layer_2_0[1999:1992]};
      btm_1[0] = {1'b0,layer_3_1[1983:1976]} - {1'b0, layer_2_1[1983:1976]};
      btm_1[1] = {1'b0,layer_3_1[1991:1984]} - {1'b0, layer_2_1[1991:1984]};
      btm_1[2] = {1'b0,layer_3_1[1999:1992]} - {1'b0, layer_2_1[1999:1992]};
      btm_2[0] = {1'b0,layer_3_2[1983:1976]} - {1'b0, layer_2_2[1983:1976]};
      btm_2[1] = {1'b0,layer_3_2[1991:1984]} - {1'b0, layer_2_2[1991:1984]};
      btm_2[2] = {1'b0,layer_3_2[1999:1992]} - {1'b0, layer_2_2[1999:1992]};
    end
    'd249: begin
      top_0[0] = {1'b0,layer_1_0[1991:1984]} - {1'b0, layer_0_0[1991:1984]};
      top_0[1] = {1'b0,layer_1_0[1999:1992]} - {1'b0, layer_0_0[1999:1992]};
      top_0[2] = {1'b0,layer_1_0[2007:2000]} - {1'b0, layer_0_0[2007:2000]};
      top_1[0] = {1'b0,layer_1_1[1991:1984]} - {1'b0, layer_0_1[1991:1984]};
      top_1[1] = {1'b0,layer_1_1[1999:1992]} - {1'b0, layer_0_1[1999:1992]};
      top_1[2] = {1'b0,layer_1_1[2007:2000]} - {1'b0, layer_0_1[2007:2000]};
      top_2[0] = {1'b0,layer_1_2[1991:1984]} - {1'b0, layer_0_2[1991:1984]};
      top_2[1] = {1'b0,layer_1_2[1999:1992]} - {1'b0, layer_0_2[1999:1992]};
      top_2[2] = {1'b0,layer_1_2[2007:2000]} - {1'b0, layer_0_2[2007:2000]};
      mid_0[0] = {1'b0,layer_2_0[1991:1984]} - {1'b0, layer_1_0[1991:1984]};
      mid_0[1] = {1'b0,layer_2_0[1999:1992]} - {1'b0, layer_1_0[1999:1992]};
      mid_0[2] = {1'b0,layer_2_0[2007:2000]} - {1'b0, layer_1_0[2007:2000]};
      mid_1[0] = {1'b0,layer_2_1[1991:1984]} - {1'b0, layer_1_1[1991:1984]};
      mid_1[1] = {1'b0,layer_2_1[1999:1992]} - {1'b0, layer_1_1[1999:1992]};
      mid_1[2] = {1'b0,layer_2_1[2007:2000]} - {1'b0, layer_1_1[2007:2000]};
      mid_2[0] = {1'b0,layer_2_2[1991:1984]} - {1'b0, layer_1_2[1991:1984]};
      mid_2[1] = {1'b0,layer_2_2[1999:1992]} - {1'b0, layer_1_2[1999:1992]};
      mid_2[2] = {1'b0,layer_2_2[2007:2000]} - {1'b0, layer_1_2[2007:2000]};
      btm_0[0] = {1'b0,layer_3_0[1991:1984]} - {1'b0, layer_2_0[1991:1984]};
      btm_0[1] = {1'b0,layer_3_0[1999:1992]} - {1'b0, layer_2_0[1999:1992]};
      btm_0[2] = {1'b0,layer_3_0[2007:2000]} - {1'b0, layer_2_0[2007:2000]};
      btm_1[0] = {1'b0,layer_3_1[1991:1984]} - {1'b0, layer_2_1[1991:1984]};
      btm_1[1] = {1'b0,layer_3_1[1999:1992]} - {1'b0, layer_2_1[1999:1992]};
      btm_1[2] = {1'b0,layer_3_1[2007:2000]} - {1'b0, layer_2_1[2007:2000]};
      btm_2[0] = {1'b0,layer_3_2[1991:1984]} - {1'b0, layer_2_2[1991:1984]};
      btm_2[1] = {1'b0,layer_3_2[1999:1992]} - {1'b0, layer_2_2[1999:1992]};
      btm_2[2] = {1'b0,layer_3_2[2007:2000]} - {1'b0, layer_2_2[2007:2000]};
    end
    'd250: begin
      top_0[0] = {1'b0,layer_1_0[1999:1992]} - {1'b0, layer_0_0[1999:1992]};
      top_0[1] = {1'b0,layer_1_0[2007:2000]} - {1'b0, layer_0_0[2007:2000]};
      top_0[2] = {1'b0,layer_1_0[2015:2008]} - {1'b0, layer_0_0[2015:2008]};
      top_1[0] = {1'b0,layer_1_1[1999:1992]} - {1'b0, layer_0_1[1999:1992]};
      top_1[1] = {1'b0,layer_1_1[2007:2000]} - {1'b0, layer_0_1[2007:2000]};
      top_1[2] = {1'b0,layer_1_1[2015:2008]} - {1'b0, layer_0_1[2015:2008]};
      top_2[0] = {1'b0,layer_1_2[1999:1992]} - {1'b0, layer_0_2[1999:1992]};
      top_2[1] = {1'b0,layer_1_2[2007:2000]} - {1'b0, layer_0_2[2007:2000]};
      top_2[2] = {1'b0,layer_1_2[2015:2008]} - {1'b0, layer_0_2[2015:2008]};
      mid_0[0] = {1'b0,layer_2_0[1999:1992]} - {1'b0, layer_1_0[1999:1992]};
      mid_0[1] = {1'b0,layer_2_0[2007:2000]} - {1'b0, layer_1_0[2007:2000]};
      mid_0[2] = {1'b0,layer_2_0[2015:2008]} - {1'b0, layer_1_0[2015:2008]};
      mid_1[0] = {1'b0,layer_2_1[1999:1992]} - {1'b0, layer_1_1[1999:1992]};
      mid_1[1] = {1'b0,layer_2_1[2007:2000]} - {1'b0, layer_1_1[2007:2000]};
      mid_1[2] = {1'b0,layer_2_1[2015:2008]} - {1'b0, layer_1_1[2015:2008]};
      mid_2[0] = {1'b0,layer_2_2[1999:1992]} - {1'b0, layer_1_2[1999:1992]};
      mid_2[1] = {1'b0,layer_2_2[2007:2000]} - {1'b0, layer_1_2[2007:2000]};
      mid_2[2] = {1'b0,layer_2_2[2015:2008]} - {1'b0, layer_1_2[2015:2008]};
      btm_0[0] = {1'b0,layer_3_0[1999:1992]} - {1'b0, layer_2_0[1999:1992]};
      btm_0[1] = {1'b0,layer_3_0[2007:2000]} - {1'b0, layer_2_0[2007:2000]};
      btm_0[2] = {1'b0,layer_3_0[2015:2008]} - {1'b0, layer_2_0[2015:2008]};
      btm_1[0] = {1'b0,layer_3_1[1999:1992]} - {1'b0, layer_2_1[1999:1992]};
      btm_1[1] = {1'b0,layer_3_1[2007:2000]} - {1'b0, layer_2_1[2007:2000]};
      btm_1[2] = {1'b0,layer_3_1[2015:2008]} - {1'b0, layer_2_1[2015:2008]};
      btm_2[0] = {1'b0,layer_3_2[1999:1992]} - {1'b0, layer_2_2[1999:1992]};
      btm_2[1] = {1'b0,layer_3_2[2007:2000]} - {1'b0, layer_2_2[2007:2000]};
      btm_2[2] = {1'b0,layer_3_2[2015:2008]} - {1'b0, layer_2_2[2015:2008]};
    end
    'd251: begin
      top_0[0] = {1'b0,layer_1_0[2007:2000]} - {1'b0, layer_0_0[2007:2000]};
      top_0[1] = {1'b0,layer_1_0[2015:2008]} - {1'b0, layer_0_0[2015:2008]};
      top_0[2] = {1'b0,layer_1_0[2023:2016]} - {1'b0, layer_0_0[2023:2016]};
      top_1[0] = {1'b0,layer_1_1[2007:2000]} - {1'b0, layer_0_1[2007:2000]};
      top_1[1] = {1'b0,layer_1_1[2015:2008]} - {1'b0, layer_0_1[2015:2008]};
      top_1[2] = {1'b0,layer_1_1[2023:2016]} - {1'b0, layer_0_1[2023:2016]};
      top_2[0] = {1'b0,layer_1_2[2007:2000]} - {1'b0, layer_0_2[2007:2000]};
      top_2[1] = {1'b0,layer_1_2[2015:2008]} - {1'b0, layer_0_2[2015:2008]};
      top_2[2] = {1'b0,layer_1_2[2023:2016]} - {1'b0, layer_0_2[2023:2016]};
      mid_0[0] = {1'b0,layer_2_0[2007:2000]} - {1'b0, layer_1_0[2007:2000]};
      mid_0[1] = {1'b0,layer_2_0[2015:2008]} - {1'b0, layer_1_0[2015:2008]};
      mid_0[2] = {1'b0,layer_2_0[2023:2016]} - {1'b0, layer_1_0[2023:2016]};
      mid_1[0] = {1'b0,layer_2_1[2007:2000]} - {1'b0, layer_1_1[2007:2000]};
      mid_1[1] = {1'b0,layer_2_1[2015:2008]} - {1'b0, layer_1_1[2015:2008]};
      mid_1[2] = {1'b0,layer_2_1[2023:2016]} - {1'b0, layer_1_1[2023:2016]};
      mid_2[0] = {1'b0,layer_2_2[2007:2000]} - {1'b0, layer_1_2[2007:2000]};
      mid_2[1] = {1'b0,layer_2_2[2015:2008]} - {1'b0, layer_1_2[2015:2008]};
      mid_2[2] = {1'b0,layer_2_2[2023:2016]} - {1'b0, layer_1_2[2023:2016]};
      btm_0[0] = {1'b0,layer_3_0[2007:2000]} - {1'b0, layer_2_0[2007:2000]};
      btm_0[1] = {1'b0,layer_3_0[2015:2008]} - {1'b0, layer_2_0[2015:2008]};
      btm_0[2] = {1'b0,layer_3_0[2023:2016]} - {1'b0, layer_2_0[2023:2016]};
      btm_1[0] = {1'b0,layer_3_1[2007:2000]} - {1'b0, layer_2_1[2007:2000]};
      btm_1[1] = {1'b0,layer_3_1[2015:2008]} - {1'b0, layer_2_1[2015:2008]};
      btm_1[2] = {1'b0,layer_3_1[2023:2016]} - {1'b0, layer_2_1[2023:2016]};
      btm_2[0] = {1'b0,layer_3_2[2007:2000]} - {1'b0, layer_2_2[2007:2000]};
      btm_2[1] = {1'b0,layer_3_2[2015:2008]} - {1'b0, layer_2_2[2015:2008]};
      btm_2[2] = {1'b0,layer_3_2[2023:2016]} - {1'b0, layer_2_2[2023:2016]};
    end
    'd252: begin
      top_0[0] = {1'b0,layer_1_0[2015:2008]} - {1'b0, layer_0_0[2015:2008]};
      top_0[1] = {1'b0,layer_1_0[2023:2016]} - {1'b0, layer_0_0[2023:2016]};
      top_0[2] = {1'b0,layer_1_0[2031:2024]} - {1'b0, layer_0_0[2031:2024]};
      top_1[0] = {1'b0,layer_1_1[2015:2008]} - {1'b0, layer_0_1[2015:2008]};
      top_1[1] = {1'b0,layer_1_1[2023:2016]} - {1'b0, layer_0_1[2023:2016]};
      top_1[2] = {1'b0,layer_1_1[2031:2024]} - {1'b0, layer_0_1[2031:2024]};
      top_2[0] = {1'b0,layer_1_2[2015:2008]} - {1'b0, layer_0_2[2015:2008]};
      top_2[1] = {1'b0,layer_1_2[2023:2016]} - {1'b0, layer_0_2[2023:2016]};
      top_2[2] = {1'b0,layer_1_2[2031:2024]} - {1'b0, layer_0_2[2031:2024]};
      mid_0[0] = {1'b0,layer_2_0[2015:2008]} - {1'b0, layer_1_0[2015:2008]};
      mid_0[1] = {1'b0,layer_2_0[2023:2016]} - {1'b0, layer_1_0[2023:2016]};
      mid_0[2] = {1'b0,layer_2_0[2031:2024]} - {1'b0, layer_1_0[2031:2024]};
      mid_1[0] = {1'b0,layer_2_1[2015:2008]} - {1'b0, layer_1_1[2015:2008]};
      mid_1[1] = {1'b0,layer_2_1[2023:2016]} - {1'b0, layer_1_1[2023:2016]};
      mid_1[2] = {1'b0,layer_2_1[2031:2024]} - {1'b0, layer_1_1[2031:2024]};
      mid_2[0] = {1'b0,layer_2_2[2015:2008]} - {1'b0, layer_1_2[2015:2008]};
      mid_2[1] = {1'b0,layer_2_2[2023:2016]} - {1'b0, layer_1_2[2023:2016]};
      mid_2[2] = {1'b0,layer_2_2[2031:2024]} - {1'b0, layer_1_2[2031:2024]};
      btm_0[0] = {1'b0,layer_3_0[2015:2008]} - {1'b0, layer_2_0[2015:2008]};
      btm_0[1] = {1'b0,layer_3_0[2023:2016]} - {1'b0, layer_2_0[2023:2016]};
      btm_0[2] = {1'b0,layer_3_0[2031:2024]} - {1'b0, layer_2_0[2031:2024]};
      btm_1[0] = {1'b0,layer_3_1[2015:2008]} - {1'b0, layer_2_1[2015:2008]};
      btm_1[1] = {1'b0,layer_3_1[2023:2016]} - {1'b0, layer_2_1[2023:2016]};
      btm_1[2] = {1'b0,layer_3_1[2031:2024]} - {1'b0, layer_2_1[2031:2024]};
      btm_2[0] = {1'b0,layer_3_2[2015:2008]} - {1'b0, layer_2_2[2015:2008]};
      btm_2[1] = {1'b0,layer_3_2[2023:2016]} - {1'b0, layer_2_2[2023:2016]};
      btm_2[2] = {1'b0,layer_3_2[2031:2024]} - {1'b0, layer_2_2[2031:2024]};
    end
    'd253: begin
      top_0[0] = {1'b0,layer_1_0[2023:2016]} - {1'b0, layer_0_0[2023:2016]};
      top_0[1] = {1'b0,layer_1_0[2031:2024]} - {1'b0, layer_0_0[2031:2024]};
      top_0[2] = {1'b0,layer_1_0[2039:2032]} - {1'b0, layer_0_0[2039:2032]};
      top_1[0] = {1'b0,layer_1_1[2023:2016]} - {1'b0, layer_0_1[2023:2016]};
      top_1[1] = {1'b0,layer_1_1[2031:2024]} - {1'b0, layer_0_1[2031:2024]};
      top_1[2] = {1'b0,layer_1_1[2039:2032]} - {1'b0, layer_0_1[2039:2032]};
      top_2[0] = {1'b0,layer_1_2[2023:2016]} - {1'b0, layer_0_2[2023:2016]};
      top_2[1] = {1'b0,layer_1_2[2031:2024]} - {1'b0, layer_0_2[2031:2024]};
      top_2[2] = {1'b0,layer_1_2[2039:2032]} - {1'b0, layer_0_2[2039:2032]};
      mid_0[0] = {1'b0,layer_2_0[2023:2016]} - {1'b0, layer_1_0[2023:2016]};
      mid_0[1] = {1'b0,layer_2_0[2031:2024]} - {1'b0, layer_1_0[2031:2024]};
      mid_0[2] = {1'b0,layer_2_0[2039:2032]} - {1'b0, layer_1_0[2039:2032]};
      mid_1[0] = {1'b0,layer_2_1[2023:2016]} - {1'b0, layer_1_1[2023:2016]};
      mid_1[1] = {1'b0,layer_2_1[2031:2024]} - {1'b0, layer_1_1[2031:2024]};
      mid_1[2] = {1'b0,layer_2_1[2039:2032]} - {1'b0, layer_1_1[2039:2032]};
      mid_2[0] = {1'b0,layer_2_2[2023:2016]} - {1'b0, layer_1_2[2023:2016]};
      mid_2[1] = {1'b0,layer_2_2[2031:2024]} - {1'b0, layer_1_2[2031:2024]};
      mid_2[2] = {1'b0,layer_2_2[2039:2032]} - {1'b0, layer_1_2[2039:2032]};
      btm_0[0] = {1'b0,layer_3_0[2023:2016]} - {1'b0, layer_2_0[2023:2016]};
      btm_0[1] = {1'b0,layer_3_0[2031:2024]} - {1'b0, layer_2_0[2031:2024]};
      btm_0[2] = {1'b0,layer_3_0[2039:2032]} - {1'b0, layer_2_0[2039:2032]};
      btm_1[0] = {1'b0,layer_3_1[2023:2016]} - {1'b0, layer_2_1[2023:2016]};
      btm_1[1] = {1'b0,layer_3_1[2031:2024]} - {1'b0, layer_2_1[2031:2024]};
      btm_1[2] = {1'b0,layer_3_1[2039:2032]} - {1'b0, layer_2_1[2039:2032]};
      btm_2[0] = {1'b0,layer_3_2[2023:2016]} - {1'b0, layer_2_2[2023:2016]};
      btm_2[1] = {1'b0,layer_3_2[2031:2024]} - {1'b0, layer_2_2[2031:2024]};
      btm_2[2] = {1'b0,layer_3_2[2039:2032]} - {1'b0, layer_2_2[2039:2032]};
    end
    'd254: begin
      top_0[0] = {1'b0,layer_1_0[2031:2024]} - {1'b0, layer_0_0[2031:2024]};
      top_0[1] = {1'b0,layer_1_0[2039:2032]} - {1'b0, layer_0_0[2039:2032]};
      top_0[2] = {1'b0,layer_1_0[2047:2040]} - {1'b0, layer_0_0[2047:2040]};
      top_1[0] = {1'b0,layer_1_1[2031:2024]} - {1'b0, layer_0_1[2031:2024]};
      top_1[1] = {1'b0,layer_1_1[2039:2032]} - {1'b0, layer_0_1[2039:2032]};
      top_1[2] = {1'b0,layer_1_1[2047:2040]} - {1'b0, layer_0_1[2047:2040]};
      top_2[0] = {1'b0,layer_1_2[2031:2024]} - {1'b0, layer_0_2[2031:2024]};
      top_2[1] = {1'b0,layer_1_2[2039:2032]} - {1'b0, layer_0_2[2039:2032]};
      top_2[2] = {1'b0,layer_1_2[2047:2040]} - {1'b0, layer_0_2[2047:2040]};
      mid_0[0] = {1'b0,layer_2_0[2031:2024]} - {1'b0, layer_1_0[2031:2024]};
      mid_0[1] = {1'b0,layer_2_0[2039:2032]} - {1'b0, layer_1_0[2039:2032]};
      mid_0[2] = {1'b0,layer_2_0[2047:2040]} - {1'b0, layer_1_0[2047:2040]};
      mid_1[0] = {1'b0,layer_2_1[2031:2024]} - {1'b0, layer_1_1[2031:2024]};
      mid_1[1] = {1'b0,layer_2_1[2039:2032]} - {1'b0, layer_1_1[2039:2032]};
      mid_1[2] = {1'b0,layer_2_1[2047:2040]} - {1'b0, layer_1_1[2047:2040]};
      mid_2[0] = {1'b0,layer_2_2[2031:2024]} - {1'b0, layer_1_2[2031:2024]};
      mid_2[1] = {1'b0,layer_2_2[2039:2032]} - {1'b0, layer_1_2[2039:2032]};
      mid_2[2] = {1'b0,layer_2_2[2047:2040]} - {1'b0, layer_1_2[2047:2040]};
      btm_0[0] = {1'b0,layer_3_0[2031:2024]} - {1'b0, layer_2_0[2031:2024]};
      btm_0[1] = {1'b0,layer_3_0[2039:2032]} - {1'b0, layer_2_0[2039:2032]};
      btm_0[2] = {1'b0,layer_3_0[2047:2040]} - {1'b0, layer_2_0[2047:2040]};
      btm_1[0] = {1'b0,layer_3_1[2031:2024]} - {1'b0, layer_2_1[2031:2024]};
      btm_1[1] = {1'b0,layer_3_1[2039:2032]} - {1'b0, layer_2_1[2039:2032]};
      btm_1[2] = {1'b0,layer_3_1[2047:2040]} - {1'b0, layer_2_1[2047:2040]};
      btm_2[0] = {1'b0,layer_3_2[2031:2024]} - {1'b0, layer_2_2[2031:2024]};
      btm_2[1] = {1'b0,layer_3_2[2039:2032]} - {1'b0, layer_2_2[2039:2032]};
      btm_2[2] = {1'b0,layer_3_2[2047:2040]} - {1'b0, layer_2_2[2047:2040]};
    end
    'd255: begin
      top_0[0] = {1'b0,layer_1_0[2039:2032]} - {1'b0, layer_0_0[2039:2032]};
      top_0[1] = {1'b0,layer_1_0[2047:2040]} - {1'b0, layer_0_0[2047:2040]};
      top_0[2] = {1'b0,layer_1_0[2055:2048]} - {1'b0, layer_0_0[2055:2048]};
      top_1[0] = {1'b0,layer_1_1[2039:2032]} - {1'b0, layer_0_1[2039:2032]};
      top_1[1] = {1'b0,layer_1_1[2047:2040]} - {1'b0, layer_0_1[2047:2040]};
      top_1[2] = {1'b0,layer_1_1[2055:2048]} - {1'b0, layer_0_1[2055:2048]};
      top_2[0] = {1'b0,layer_1_2[2039:2032]} - {1'b0, layer_0_2[2039:2032]};
      top_2[1] = {1'b0,layer_1_2[2047:2040]} - {1'b0, layer_0_2[2047:2040]};
      top_2[2] = {1'b0,layer_1_2[2055:2048]} - {1'b0, layer_0_2[2055:2048]};
      mid_0[0] = {1'b0,layer_2_0[2039:2032]} - {1'b0, layer_1_0[2039:2032]};
      mid_0[1] = {1'b0,layer_2_0[2047:2040]} - {1'b0, layer_1_0[2047:2040]};
      mid_0[2] = {1'b0,layer_2_0[2055:2048]} - {1'b0, layer_1_0[2055:2048]};
      mid_1[0] = {1'b0,layer_2_1[2039:2032]} - {1'b0, layer_1_1[2039:2032]};
      mid_1[1] = {1'b0,layer_2_1[2047:2040]} - {1'b0, layer_1_1[2047:2040]};
      mid_1[2] = {1'b0,layer_2_1[2055:2048]} - {1'b0, layer_1_1[2055:2048]};
      mid_2[0] = {1'b0,layer_2_2[2039:2032]} - {1'b0, layer_1_2[2039:2032]};
      mid_2[1] = {1'b0,layer_2_2[2047:2040]} - {1'b0, layer_1_2[2047:2040]};
      mid_2[2] = {1'b0,layer_2_2[2055:2048]} - {1'b0, layer_1_2[2055:2048]};
      btm_0[0] = {1'b0,layer_3_0[2039:2032]} - {1'b0, layer_2_0[2039:2032]};
      btm_0[1] = {1'b0,layer_3_0[2047:2040]} - {1'b0, layer_2_0[2047:2040]};
      btm_0[2] = {1'b0,layer_3_0[2055:2048]} - {1'b0, layer_2_0[2055:2048]};
      btm_1[0] = {1'b0,layer_3_1[2039:2032]} - {1'b0, layer_2_1[2039:2032]};
      btm_1[1] = {1'b0,layer_3_1[2047:2040]} - {1'b0, layer_2_1[2047:2040]};
      btm_1[2] = {1'b0,layer_3_1[2055:2048]} - {1'b0, layer_2_1[2055:2048]};
      btm_2[0] = {1'b0,layer_3_2[2039:2032]} - {1'b0, layer_2_2[2039:2032]};
      btm_2[1] = {1'b0,layer_3_2[2047:2040]} - {1'b0, layer_2_2[2047:2040]};
      btm_2[2] = {1'b0,layer_3_2[2055:2048]} - {1'b0, layer_2_2[2055:2048]};
    end
    'd256: begin
      top_0[0] = {1'b0,layer_1_0[2047:2040]} - {1'b0, layer_0_0[2047:2040]};
      top_0[1] = {1'b0,layer_1_0[2055:2048]} - {1'b0, layer_0_0[2055:2048]};
      top_0[2] = {1'b0,layer_1_0[2063:2056]} - {1'b0, layer_0_0[2063:2056]};
      top_1[0] = {1'b0,layer_1_1[2047:2040]} - {1'b0, layer_0_1[2047:2040]};
      top_1[1] = {1'b0,layer_1_1[2055:2048]} - {1'b0, layer_0_1[2055:2048]};
      top_1[2] = {1'b0,layer_1_1[2063:2056]} - {1'b0, layer_0_1[2063:2056]};
      top_2[0] = {1'b0,layer_1_2[2047:2040]} - {1'b0, layer_0_2[2047:2040]};
      top_2[1] = {1'b0,layer_1_2[2055:2048]} - {1'b0, layer_0_2[2055:2048]};
      top_2[2] = {1'b0,layer_1_2[2063:2056]} - {1'b0, layer_0_2[2063:2056]};
      mid_0[0] = {1'b0,layer_2_0[2047:2040]} - {1'b0, layer_1_0[2047:2040]};
      mid_0[1] = {1'b0,layer_2_0[2055:2048]} - {1'b0, layer_1_0[2055:2048]};
      mid_0[2] = {1'b0,layer_2_0[2063:2056]} - {1'b0, layer_1_0[2063:2056]};
      mid_1[0] = {1'b0,layer_2_1[2047:2040]} - {1'b0, layer_1_1[2047:2040]};
      mid_1[1] = {1'b0,layer_2_1[2055:2048]} - {1'b0, layer_1_1[2055:2048]};
      mid_1[2] = {1'b0,layer_2_1[2063:2056]} - {1'b0, layer_1_1[2063:2056]};
      mid_2[0] = {1'b0,layer_2_2[2047:2040]} - {1'b0, layer_1_2[2047:2040]};
      mid_2[1] = {1'b0,layer_2_2[2055:2048]} - {1'b0, layer_1_2[2055:2048]};
      mid_2[2] = {1'b0,layer_2_2[2063:2056]} - {1'b0, layer_1_2[2063:2056]};
      btm_0[0] = {1'b0,layer_3_0[2047:2040]} - {1'b0, layer_2_0[2047:2040]};
      btm_0[1] = {1'b0,layer_3_0[2055:2048]} - {1'b0, layer_2_0[2055:2048]};
      btm_0[2] = {1'b0,layer_3_0[2063:2056]} - {1'b0, layer_2_0[2063:2056]};
      btm_1[0] = {1'b0,layer_3_1[2047:2040]} - {1'b0, layer_2_1[2047:2040]};
      btm_1[1] = {1'b0,layer_3_1[2055:2048]} - {1'b0, layer_2_1[2055:2048]};
      btm_1[2] = {1'b0,layer_3_1[2063:2056]} - {1'b0, layer_2_1[2063:2056]};
      btm_2[0] = {1'b0,layer_3_2[2047:2040]} - {1'b0, layer_2_2[2047:2040]};
      btm_2[1] = {1'b0,layer_3_2[2055:2048]} - {1'b0, layer_2_2[2055:2048]};
      btm_2[2] = {1'b0,layer_3_2[2063:2056]} - {1'b0, layer_2_2[2063:2056]};
    end
    'd257: begin
      top_0[0] = {1'b0,layer_1_0[2055:2048]} - {1'b0, layer_0_0[2055:2048]};
      top_0[1] = {1'b0,layer_1_0[2063:2056]} - {1'b0, layer_0_0[2063:2056]};
      top_0[2] = {1'b0,layer_1_0[2071:2064]} - {1'b0, layer_0_0[2071:2064]};
      top_1[0] = {1'b0,layer_1_1[2055:2048]} - {1'b0, layer_0_1[2055:2048]};
      top_1[1] = {1'b0,layer_1_1[2063:2056]} - {1'b0, layer_0_1[2063:2056]};
      top_1[2] = {1'b0,layer_1_1[2071:2064]} - {1'b0, layer_0_1[2071:2064]};
      top_2[0] = {1'b0,layer_1_2[2055:2048]} - {1'b0, layer_0_2[2055:2048]};
      top_2[1] = {1'b0,layer_1_2[2063:2056]} - {1'b0, layer_0_2[2063:2056]};
      top_2[2] = {1'b0,layer_1_2[2071:2064]} - {1'b0, layer_0_2[2071:2064]};
      mid_0[0] = {1'b0,layer_2_0[2055:2048]} - {1'b0, layer_1_0[2055:2048]};
      mid_0[1] = {1'b0,layer_2_0[2063:2056]} - {1'b0, layer_1_0[2063:2056]};
      mid_0[2] = {1'b0,layer_2_0[2071:2064]} - {1'b0, layer_1_0[2071:2064]};
      mid_1[0] = {1'b0,layer_2_1[2055:2048]} - {1'b0, layer_1_1[2055:2048]};
      mid_1[1] = {1'b0,layer_2_1[2063:2056]} - {1'b0, layer_1_1[2063:2056]};
      mid_1[2] = {1'b0,layer_2_1[2071:2064]} - {1'b0, layer_1_1[2071:2064]};
      mid_2[0] = {1'b0,layer_2_2[2055:2048]} - {1'b0, layer_1_2[2055:2048]};
      mid_2[1] = {1'b0,layer_2_2[2063:2056]} - {1'b0, layer_1_2[2063:2056]};
      mid_2[2] = {1'b0,layer_2_2[2071:2064]} - {1'b0, layer_1_2[2071:2064]};
      btm_0[0] = {1'b0,layer_3_0[2055:2048]} - {1'b0, layer_2_0[2055:2048]};
      btm_0[1] = {1'b0,layer_3_0[2063:2056]} - {1'b0, layer_2_0[2063:2056]};
      btm_0[2] = {1'b0,layer_3_0[2071:2064]} - {1'b0, layer_2_0[2071:2064]};
      btm_1[0] = {1'b0,layer_3_1[2055:2048]} - {1'b0, layer_2_1[2055:2048]};
      btm_1[1] = {1'b0,layer_3_1[2063:2056]} - {1'b0, layer_2_1[2063:2056]};
      btm_1[2] = {1'b0,layer_3_1[2071:2064]} - {1'b0, layer_2_1[2071:2064]};
      btm_2[0] = {1'b0,layer_3_2[2055:2048]} - {1'b0, layer_2_2[2055:2048]};
      btm_2[1] = {1'b0,layer_3_2[2063:2056]} - {1'b0, layer_2_2[2063:2056]};
      btm_2[2] = {1'b0,layer_3_2[2071:2064]} - {1'b0, layer_2_2[2071:2064]};
    end
    'd258: begin
      top_0[0] = {1'b0,layer_1_0[2063:2056]} - {1'b0, layer_0_0[2063:2056]};
      top_0[1] = {1'b0,layer_1_0[2071:2064]} - {1'b0, layer_0_0[2071:2064]};
      top_0[2] = {1'b0,layer_1_0[2079:2072]} - {1'b0, layer_0_0[2079:2072]};
      top_1[0] = {1'b0,layer_1_1[2063:2056]} - {1'b0, layer_0_1[2063:2056]};
      top_1[1] = {1'b0,layer_1_1[2071:2064]} - {1'b0, layer_0_1[2071:2064]};
      top_1[2] = {1'b0,layer_1_1[2079:2072]} - {1'b0, layer_0_1[2079:2072]};
      top_2[0] = {1'b0,layer_1_2[2063:2056]} - {1'b0, layer_0_2[2063:2056]};
      top_2[1] = {1'b0,layer_1_2[2071:2064]} - {1'b0, layer_0_2[2071:2064]};
      top_2[2] = {1'b0,layer_1_2[2079:2072]} - {1'b0, layer_0_2[2079:2072]};
      mid_0[0] = {1'b0,layer_2_0[2063:2056]} - {1'b0, layer_1_0[2063:2056]};
      mid_0[1] = {1'b0,layer_2_0[2071:2064]} - {1'b0, layer_1_0[2071:2064]};
      mid_0[2] = {1'b0,layer_2_0[2079:2072]} - {1'b0, layer_1_0[2079:2072]};
      mid_1[0] = {1'b0,layer_2_1[2063:2056]} - {1'b0, layer_1_1[2063:2056]};
      mid_1[1] = {1'b0,layer_2_1[2071:2064]} - {1'b0, layer_1_1[2071:2064]};
      mid_1[2] = {1'b0,layer_2_1[2079:2072]} - {1'b0, layer_1_1[2079:2072]};
      mid_2[0] = {1'b0,layer_2_2[2063:2056]} - {1'b0, layer_1_2[2063:2056]};
      mid_2[1] = {1'b0,layer_2_2[2071:2064]} - {1'b0, layer_1_2[2071:2064]};
      mid_2[2] = {1'b0,layer_2_2[2079:2072]} - {1'b0, layer_1_2[2079:2072]};
      btm_0[0] = {1'b0,layer_3_0[2063:2056]} - {1'b0, layer_2_0[2063:2056]};
      btm_0[1] = {1'b0,layer_3_0[2071:2064]} - {1'b0, layer_2_0[2071:2064]};
      btm_0[2] = {1'b0,layer_3_0[2079:2072]} - {1'b0, layer_2_0[2079:2072]};
      btm_1[0] = {1'b0,layer_3_1[2063:2056]} - {1'b0, layer_2_1[2063:2056]};
      btm_1[1] = {1'b0,layer_3_1[2071:2064]} - {1'b0, layer_2_1[2071:2064]};
      btm_1[2] = {1'b0,layer_3_1[2079:2072]} - {1'b0, layer_2_1[2079:2072]};
      btm_2[0] = {1'b0,layer_3_2[2063:2056]} - {1'b0, layer_2_2[2063:2056]};
      btm_2[1] = {1'b0,layer_3_2[2071:2064]} - {1'b0, layer_2_2[2071:2064]};
      btm_2[2] = {1'b0,layer_3_2[2079:2072]} - {1'b0, layer_2_2[2079:2072]};
    end
    'd259: begin
      top_0[0] = {1'b0,layer_1_0[2071:2064]} - {1'b0, layer_0_0[2071:2064]};
      top_0[1] = {1'b0,layer_1_0[2079:2072]} - {1'b0, layer_0_0[2079:2072]};
      top_0[2] = {1'b0,layer_1_0[2087:2080]} - {1'b0, layer_0_0[2087:2080]};
      top_1[0] = {1'b0,layer_1_1[2071:2064]} - {1'b0, layer_0_1[2071:2064]};
      top_1[1] = {1'b0,layer_1_1[2079:2072]} - {1'b0, layer_0_1[2079:2072]};
      top_1[2] = {1'b0,layer_1_1[2087:2080]} - {1'b0, layer_0_1[2087:2080]};
      top_2[0] = {1'b0,layer_1_2[2071:2064]} - {1'b0, layer_0_2[2071:2064]};
      top_2[1] = {1'b0,layer_1_2[2079:2072]} - {1'b0, layer_0_2[2079:2072]};
      top_2[2] = {1'b0,layer_1_2[2087:2080]} - {1'b0, layer_0_2[2087:2080]};
      mid_0[0] = {1'b0,layer_2_0[2071:2064]} - {1'b0, layer_1_0[2071:2064]};
      mid_0[1] = {1'b0,layer_2_0[2079:2072]} - {1'b0, layer_1_0[2079:2072]};
      mid_0[2] = {1'b0,layer_2_0[2087:2080]} - {1'b0, layer_1_0[2087:2080]};
      mid_1[0] = {1'b0,layer_2_1[2071:2064]} - {1'b0, layer_1_1[2071:2064]};
      mid_1[1] = {1'b0,layer_2_1[2079:2072]} - {1'b0, layer_1_1[2079:2072]};
      mid_1[2] = {1'b0,layer_2_1[2087:2080]} - {1'b0, layer_1_1[2087:2080]};
      mid_2[0] = {1'b0,layer_2_2[2071:2064]} - {1'b0, layer_1_2[2071:2064]};
      mid_2[1] = {1'b0,layer_2_2[2079:2072]} - {1'b0, layer_1_2[2079:2072]};
      mid_2[2] = {1'b0,layer_2_2[2087:2080]} - {1'b0, layer_1_2[2087:2080]};
      btm_0[0] = {1'b0,layer_3_0[2071:2064]} - {1'b0, layer_2_0[2071:2064]};
      btm_0[1] = {1'b0,layer_3_0[2079:2072]} - {1'b0, layer_2_0[2079:2072]};
      btm_0[2] = {1'b0,layer_3_0[2087:2080]} - {1'b0, layer_2_0[2087:2080]};
      btm_1[0] = {1'b0,layer_3_1[2071:2064]} - {1'b0, layer_2_1[2071:2064]};
      btm_1[1] = {1'b0,layer_3_1[2079:2072]} - {1'b0, layer_2_1[2079:2072]};
      btm_1[2] = {1'b0,layer_3_1[2087:2080]} - {1'b0, layer_2_1[2087:2080]};
      btm_2[0] = {1'b0,layer_3_2[2071:2064]} - {1'b0, layer_2_2[2071:2064]};
      btm_2[1] = {1'b0,layer_3_2[2079:2072]} - {1'b0, layer_2_2[2079:2072]};
      btm_2[2] = {1'b0,layer_3_2[2087:2080]} - {1'b0, layer_2_2[2087:2080]};
    end
    'd260: begin
      top_0[0] = {1'b0,layer_1_0[2079:2072]} - {1'b0, layer_0_0[2079:2072]};
      top_0[1] = {1'b0,layer_1_0[2087:2080]} - {1'b0, layer_0_0[2087:2080]};
      top_0[2] = {1'b0,layer_1_0[2095:2088]} - {1'b0, layer_0_0[2095:2088]};
      top_1[0] = {1'b0,layer_1_1[2079:2072]} - {1'b0, layer_0_1[2079:2072]};
      top_1[1] = {1'b0,layer_1_1[2087:2080]} - {1'b0, layer_0_1[2087:2080]};
      top_1[2] = {1'b0,layer_1_1[2095:2088]} - {1'b0, layer_0_1[2095:2088]};
      top_2[0] = {1'b0,layer_1_2[2079:2072]} - {1'b0, layer_0_2[2079:2072]};
      top_2[1] = {1'b0,layer_1_2[2087:2080]} - {1'b0, layer_0_2[2087:2080]};
      top_2[2] = {1'b0,layer_1_2[2095:2088]} - {1'b0, layer_0_2[2095:2088]};
      mid_0[0] = {1'b0,layer_2_0[2079:2072]} - {1'b0, layer_1_0[2079:2072]};
      mid_0[1] = {1'b0,layer_2_0[2087:2080]} - {1'b0, layer_1_0[2087:2080]};
      mid_0[2] = {1'b0,layer_2_0[2095:2088]} - {1'b0, layer_1_0[2095:2088]};
      mid_1[0] = {1'b0,layer_2_1[2079:2072]} - {1'b0, layer_1_1[2079:2072]};
      mid_1[1] = {1'b0,layer_2_1[2087:2080]} - {1'b0, layer_1_1[2087:2080]};
      mid_1[2] = {1'b0,layer_2_1[2095:2088]} - {1'b0, layer_1_1[2095:2088]};
      mid_2[0] = {1'b0,layer_2_2[2079:2072]} - {1'b0, layer_1_2[2079:2072]};
      mid_2[1] = {1'b0,layer_2_2[2087:2080]} - {1'b0, layer_1_2[2087:2080]};
      mid_2[2] = {1'b0,layer_2_2[2095:2088]} - {1'b0, layer_1_2[2095:2088]};
      btm_0[0] = {1'b0,layer_3_0[2079:2072]} - {1'b0, layer_2_0[2079:2072]};
      btm_0[1] = {1'b0,layer_3_0[2087:2080]} - {1'b0, layer_2_0[2087:2080]};
      btm_0[2] = {1'b0,layer_3_0[2095:2088]} - {1'b0, layer_2_0[2095:2088]};
      btm_1[0] = {1'b0,layer_3_1[2079:2072]} - {1'b0, layer_2_1[2079:2072]};
      btm_1[1] = {1'b0,layer_3_1[2087:2080]} - {1'b0, layer_2_1[2087:2080]};
      btm_1[2] = {1'b0,layer_3_1[2095:2088]} - {1'b0, layer_2_1[2095:2088]};
      btm_2[0] = {1'b0,layer_3_2[2079:2072]} - {1'b0, layer_2_2[2079:2072]};
      btm_2[1] = {1'b0,layer_3_2[2087:2080]} - {1'b0, layer_2_2[2087:2080]};
      btm_2[2] = {1'b0,layer_3_2[2095:2088]} - {1'b0, layer_2_2[2095:2088]};
    end
    'd261: begin
      top_0[0] = {1'b0,layer_1_0[2087:2080]} - {1'b0, layer_0_0[2087:2080]};
      top_0[1] = {1'b0,layer_1_0[2095:2088]} - {1'b0, layer_0_0[2095:2088]};
      top_0[2] = {1'b0,layer_1_0[2103:2096]} - {1'b0, layer_0_0[2103:2096]};
      top_1[0] = {1'b0,layer_1_1[2087:2080]} - {1'b0, layer_0_1[2087:2080]};
      top_1[1] = {1'b0,layer_1_1[2095:2088]} - {1'b0, layer_0_1[2095:2088]};
      top_1[2] = {1'b0,layer_1_1[2103:2096]} - {1'b0, layer_0_1[2103:2096]};
      top_2[0] = {1'b0,layer_1_2[2087:2080]} - {1'b0, layer_0_2[2087:2080]};
      top_2[1] = {1'b0,layer_1_2[2095:2088]} - {1'b0, layer_0_2[2095:2088]};
      top_2[2] = {1'b0,layer_1_2[2103:2096]} - {1'b0, layer_0_2[2103:2096]};
      mid_0[0] = {1'b0,layer_2_0[2087:2080]} - {1'b0, layer_1_0[2087:2080]};
      mid_0[1] = {1'b0,layer_2_0[2095:2088]} - {1'b0, layer_1_0[2095:2088]};
      mid_0[2] = {1'b0,layer_2_0[2103:2096]} - {1'b0, layer_1_0[2103:2096]};
      mid_1[0] = {1'b0,layer_2_1[2087:2080]} - {1'b0, layer_1_1[2087:2080]};
      mid_1[1] = {1'b0,layer_2_1[2095:2088]} - {1'b0, layer_1_1[2095:2088]};
      mid_1[2] = {1'b0,layer_2_1[2103:2096]} - {1'b0, layer_1_1[2103:2096]};
      mid_2[0] = {1'b0,layer_2_2[2087:2080]} - {1'b0, layer_1_2[2087:2080]};
      mid_2[1] = {1'b0,layer_2_2[2095:2088]} - {1'b0, layer_1_2[2095:2088]};
      mid_2[2] = {1'b0,layer_2_2[2103:2096]} - {1'b0, layer_1_2[2103:2096]};
      btm_0[0] = {1'b0,layer_3_0[2087:2080]} - {1'b0, layer_2_0[2087:2080]};
      btm_0[1] = {1'b0,layer_3_0[2095:2088]} - {1'b0, layer_2_0[2095:2088]};
      btm_0[2] = {1'b0,layer_3_0[2103:2096]} - {1'b0, layer_2_0[2103:2096]};
      btm_1[0] = {1'b0,layer_3_1[2087:2080]} - {1'b0, layer_2_1[2087:2080]};
      btm_1[1] = {1'b0,layer_3_1[2095:2088]} - {1'b0, layer_2_1[2095:2088]};
      btm_1[2] = {1'b0,layer_3_1[2103:2096]} - {1'b0, layer_2_1[2103:2096]};
      btm_2[0] = {1'b0,layer_3_2[2087:2080]} - {1'b0, layer_2_2[2087:2080]};
      btm_2[1] = {1'b0,layer_3_2[2095:2088]} - {1'b0, layer_2_2[2095:2088]};
      btm_2[2] = {1'b0,layer_3_2[2103:2096]} - {1'b0, layer_2_2[2103:2096]};
    end
    'd262: begin
      top_0[0] = {1'b0,layer_1_0[2095:2088]} - {1'b0, layer_0_0[2095:2088]};
      top_0[1] = {1'b0,layer_1_0[2103:2096]} - {1'b0, layer_0_0[2103:2096]};
      top_0[2] = {1'b0,layer_1_0[2111:2104]} - {1'b0, layer_0_0[2111:2104]};
      top_1[0] = {1'b0,layer_1_1[2095:2088]} - {1'b0, layer_0_1[2095:2088]};
      top_1[1] = {1'b0,layer_1_1[2103:2096]} - {1'b0, layer_0_1[2103:2096]};
      top_1[2] = {1'b0,layer_1_1[2111:2104]} - {1'b0, layer_0_1[2111:2104]};
      top_2[0] = {1'b0,layer_1_2[2095:2088]} - {1'b0, layer_0_2[2095:2088]};
      top_2[1] = {1'b0,layer_1_2[2103:2096]} - {1'b0, layer_0_2[2103:2096]};
      top_2[2] = {1'b0,layer_1_2[2111:2104]} - {1'b0, layer_0_2[2111:2104]};
      mid_0[0] = {1'b0,layer_2_0[2095:2088]} - {1'b0, layer_1_0[2095:2088]};
      mid_0[1] = {1'b0,layer_2_0[2103:2096]} - {1'b0, layer_1_0[2103:2096]};
      mid_0[2] = {1'b0,layer_2_0[2111:2104]} - {1'b0, layer_1_0[2111:2104]};
      mid_1[0] = {1'b0,layer_2_1[2095:2088]} - {1'b0, layer_1_1[2095:2088]};
      mid_1[1] = {1'b0,layer_2_1[2103:2096]} - {1'b0, layer_1_1[2103:2096]};
      mid_1[2] = {1'b0,layer_2_1[2111:2104]} - {1'b0, layer_1_1[2111:2104]};
      mid_2[0] = {1'b0,layer_2_2[2095:2088]} - {1'b0, layer_1_2[2095:2088]};
      mid_2[1] = {1'b0,layer_2_2[2103:2096]} - {1'b0, layer_1_2[2103:2096]};
      mid_2[2] = {1'b0,layer_2_2[2111:2104]} - {1'b0, layer_1_2[2111:2104]};
      btm_0[0] = {1'b0,layer_3_0[2095:2088]} - {1'b0, layer_2_0[2095:2088]};
      btm_0[1] = {1'b0,layer_3_0[2103:2096]} - {1'b0, layer_2_0[2103:2096]};
      btm_0[2] = {1'b0,layer_3_0[2111:2104]} - {1'b0, layer_2_0[2111:2104]};
      btm_1[0] = {1'b0,layer_3_1[2095:2088]} - {1'b0, layer_2_1[2095:2088]};
      btm_1[1] = {1'b0,layer_3_1[2103:2096]} - {1'b0, layer_2_1[2103:2096]};
      btm_1[2] = {1'b0,layer_3_1[2111:2104]} - {1'b0, layer_2_1[2111:2104]};
      btm_2[0] = {1'b0,layer_3_2[2095:2088]} - {1'b0, layer_2_2[2095:2088]};
      btm_2[1] = {1'b0,layer_3_2[2103:2096]} - {1'b0, layer_2_2[2103:2096]};
      btm_2[2] = {1'b0,layer_3_2[2111:2104]} - {1'b0, layer_2_2[2111:2104]};
    end
    'd263: begin
      top_0[0] = {1'b0,layer_1_0[2103:2096]} - {1'b0, layer_0_0[2103:2096]};
      top_0[1] = {1'b0,layer_1_0[2111:2104]} - {1'b0, layer_0_0[2111:2104]};
      top_0[2] = {1'b0,layer_1_0[2119:2112]} - {1'b0, layer_0_0[2119:2112]};
      top_1[0] = {1'b0,layer_1_1[2103:2096]} - {1'b0, layer_0_1[2103:2096]};
      top_1[1] = {1'b0,layer_1_1[2111:2104]} - {1'b0, layer_0_1[2111:2104]};
      top_1[2] = {1'b0,layer_1_1[2119:2112]} - {1'b0, layer_0_1[2119:2112]};
      top_2[0] = {1'b0,layer_1_2[2103:2096]} - {1'b0, layer_0_2[2103:2096]};
      top_2[1] = {1'b0,layer_1_2[2111:2104]} - {1'b0, layer_0_2[2111:2104]};
      top_2[2] = {1'b0,layer_1_2[2119:2112]} - {1'b0, layer_0_2[2119:2112]};
      mid_0[0] = {1'b0,layer_2_0[2103:2096]} - {1'b0, layer_1_0[2103:2096]};
      mid_0[1] = {1'b0,layer_2_0[2111:2104]} - {1'b0, layer_1_0[2111:2104]};
      mid_0[2] = {1'b0,layer_2_0[2119:2112]} - {1'b0, layer_1_0[2119:2112]};
      mid_1[0] = {1'b0,layer_2_1[2103:2096]} - {1'b0, layer_1_1[2103:2096]};
      mid_1[1] = {1'b0,layer_2_1[2111:2104]} - {1'b0, layer_1_1[2111:2104]};
      mid_1[2] = {1'b0,layer_2_1[2119:2112]} - {1'b0, layer_1_1[2119:2112]};
      mid_2[0] = {1'b0,layer_2_2[2103:2096]} - {1'b0, layer_1_2[2103:2096]};
      mid_2[1] = {1'b0,layer_2_2[2111:2104]} - {1'b0, layer_1_2[2111:2104]};
      mid_2[2] = {1'b0,layer_2_2[2119:2112]} - {1'b0, layer_1_2[2119:2112]};
      btm_0[0] = {1'b0,layer_3_0[2103:2096]} - {1'b0, layer_2_0[2103:2096]};
      btm_0[1] = {1'b0,layer_3_0[2111:2104]} - {1'b0, layer_2_0[2111:2104]};
      btm_0[2] = {1'b0,layer_3_0[2119:2112]} - {1'b0, layer_2_0[2119:2112]};
      btm_1[0] = {1'b0,layer_3_1[2103:2096]} - {1'b0, layer_2_1[2103:2096]};
      btm_1[1] = {1'b0,layer_3_1[2111:2104]} - {1'b0, layer_2_1[2111:2104]};
      btm_1[2] = {1'b0,layer_3_1[2119:2112]} - {1'b0, layer_2_1[2119:2112]};
      btm_2[0] = {1'b0,layer_3_2[2103:2096]} - {1'b0, layer_2_2[2103:2096]};
      btm_2[1] = {1'b0,layer_3_2[2111:2104]} - {1'b0, layer_2_2[2111:2104]};
      btm_2[2] = {1'b0,layer_3_2[2119:2112]} - {1'b0, layer_2_2[2119:2112]};
    end
    'd264: begin
      top_0[0] = {1'b0,layer_1_0[2111:2104]} - {1'b0, layer_0_0[2111:2104]};
      top_0[1] = {1'b0,layer_1_0[2119:2112]} - {1'b0, layer_0_0[2119:2112]};
      top_0[2] = {1'b0,layer_1_0[2127:2120]} - {1'b0, layer_0_0[2127:2120]};
      top_1[0] = {1'b0,layer_1_1[2111:2104]} - {1'b0, layer_0_1[2111:2104]};
      top_1[1] = {1'b0,layer_1_1[2119:2112]} - {1'b0, layer_0_1[2119:2112]};
      top_1[2] = {1'b0,layer_1_1[2127:2120]} - {1'b0, layer_0_1[2127:2120]};
      top_2[0] = {1'b0,layer_1_2[2111:2104]} - {1'b0, layer_0_2[2111:2104]};
      top_2[1] = {1'b0,layer_1_2[2119:2112]} - {1'b0, layer_0_2[2119:2112]};
      top_2[2] = {1'b0,layer_1_2[2127:2120]} - {1'b0, layer_0_2[2127:2120]};
      mid_0[0] = {1'b0,layer_2_0[2111:2104]} - {1'b0, layer_1_0[2111:2104]};
      mid_0[1] = {1'b0,layer_2_0[2119:2112]} - {1'b0, layer_1_0[2119:2112]};
      mid_0[2] = {1'b0,layer_2_0[2127:2120]} - {1'b0, layer_1_0[2127:2120]};
      mid_1[0] = {1'b0,layer_2_1[2111:2104]} - {1'b0, layer_1_1[2111:2104]};
      mid_1[1] = {1'b0,layer_2_1[2119:2112]} - {1'b0, layer_1_1[2119:2112]};
      mid_1[2] = {1'b0,layer_2_1[2127:2120]} - {1'b0, layer_1_1[2127:2120]};
      mid_2[0] = {1'b0,layer_2_2[2111:2104]} - {1'b0, layer_1_2[2111:2104]};
      mid_2[1] = {1'b0,layer_2_2[2119:2112]} - {1'b0, layer_1_2[2119:2112]};
      mid_2[2] = {1'b0,layer_2_2[2127:2120]} - {1'b0, layer_1_2[2127:2120]};
      btm_0[0] = {1'b0,layer_3_0[2111:2104]} - {1'b0, layer_2_0[2111:2104]};
      btm_0[1] = {1'b0,layer_3_0[2119:2112]} - {1'b0, layer_2_0[2119:2112]};
      btm_0[2] = {1'b0,layer_3_0[2127:2120]} - {1'b0, layer_2_0[2127:2120]};
      btm_1[0] = {1'b0,layer_3_1[2111:2104]} - {1'b0, layer_2_1[2111:2104]};
      btm_1[1] = {1'b0,layer_3_1[2119:2112]} - {1'b0, layer_2_1[2119:2112]};
      btm_1[2] = {1'b0,layer_3_1[2127:2120]} - {1'b0, layer_2_1[2127:2120]};
      btm_2[0] = {1'b0,layer_3_2[2111:2104]} - {1'b0, layer_2_2[2111:2104]};
      btm_2[1] = {1'b0,layer_3_2[2119:2112]} - {1'b0, layer_2_2[2119:2112]};
      btm_2[2] = {1'b0,layer_3_2[2127:2120]} - {1'b0, layer_2_2[2127:2120]};
    end
    'd265: begin
      top_0[0] = {1'b0,layer_1_0[2119:2112]} - {1'b0, layer_0_0[2119:2112]};
      top_0[1] = {1'b0,layer_1_0[2127:2120]} - {1'b0, layer_0_0[2127:2120]};
      top_0[2] = {1'b0,layer_1_0[2135:2128]} - {1'b0, layer_0_0[2135:2128]};
      top_1[0] = {1'b0,layer_1_1[2119:2112]} - {1'b0, layer_0_1[2119:2112]};
      top_1[1] = {1'b0,layer_1_1[2127:2120]} - {1'b0, layer_0_1[2127:2120]};
      top_1[2] = {1'b0,layer_1_1[2135:2128]} - {1'b0, layer_0_1[2135:2128]};
      top_2[0] = {1'b0,layer_1_2[2119:2112]} - {1'b0, layer_0_2[2119:2112]};
      top_2[1] = {1'b0,layer_1_2[2127:2120]} - {1'b0, layer_0_2[2127:2120]};
      top_2[2] = {1'b0,layer_1_2[2135:2128]} - {1'b0, layer_0_2[2135:2128]};
      mid_0[0] = {1'b0,layer_2_0[2119:2112]} - {1'b0, layer_1_0[2119:2112]};
      mid_0[1] = {1'b0,layer_2_0[2127:2120]} - {1'b0, layer_1_0[2127:2120]};
      mid_0[2] = {1'b0,layer_2_0[2135:2128]} - {1'b0, layer_1_0[2135:2128]};
      mid_1[0] = {1'b0,layer_2_1[2119:2112]} - {1'b0, layer_1_1[2119:2112]};
      mid_1[1] = {1'b0,layer_2_1[2127:2120]} - {1'b0, layer_1_1[2127:2120]};
      mid_1[2] = {1'b0,layer_2_1[2135:2128]} - {1'b0, layer_1_1[2135:2128]};
      mid_2[0] = {1'b0,layer_2_2[2119:2112]} - {1'b0, layer_1_2[2119:2112]};
      mid_2[1] = {1'b0,layer_2_2[2127:2120]} - {1'b0, layer_1_2[2127:2120]};
      mid_2[2] = {1'b0,layer_2_2[2135:2128]} - {1'b0, layer_1_2[2135:2128]};
      btm_0[0] = {1'b0,layer_3_0[2119:2112]} - {1'b0, layer_2_0[2119:2112]};
      btm_0[1] = {1'b0,layer_3_0[2127:2120]} - {1'b0, layer_2_0[2127:2120]};
      btm_0[2] = {1'b0,layer_3_0[2135:2128]} - {1'b0, layer_2_0[2135:2128]};
      btm_1[0] = {1'b0,layer_3_1[2119:2112]} - {1'b0, layer_2_1[2119:2112]};
      btm_1[1] = {1'b0,layer_3_1[2127:2120]} - {1'b0, layer_2_1[2127:2120]};
      btm_1[2] = {1'b0,layer_3_1[2135:2128]} - {1'b0, layer_2_1[2135:2128]};
      btm_2[0] = {1'b0,layer_3_2[2119:2112]} - {1'b0, layer_2_2[2119:2112]};
      btm_2[1] = {1'b0,layer_3_2[2127:2120]} - {1'b0, layer_2_2[2127:2120]};
      btm_2[2] = {1'b0,layer_3_2[2135:2128]} - {1'b0, layer_2_2[2135:2128]};
    end
    'd266: begin
      top_0[0] = {1'b0,layer_1_0[2127:2120]} - {1'b0, layer_0_0[2127:2120]};
      top_0[1] = {1'b0,layer_1_0[2135:2128]} - {1'b0, layer_0_0[2135:2128]};
      top_0[2] = {1'b0,layer_1_0[2143:2136]} - {1'b0, layer_0_0[2143:2136]};
      top_1[0] = {1'b0,layer_1_1[2127:2120]} - {1'b0, layer_0_1[2127:2120]};
      top_1[1] = {1'b0,layer_1_1[2135:2128]} - {1'b0, layer_0_1[2135:2128]};
      top_1[2] = {1'b0,layer_1_1[2143:2136]} - {1'b0, layer_0_1[2143:2136]};
      top_2[0] = {1'b0,layer_1_2[2127:2120]} - {1'b0, layer_0_2[2127:2120]};
      top_2[1] = {1'b0,layer_1_2[2135:2128]} - {1'b0, layer_0_2[2135:2128]};
      top_2[2] = {1'b0,layer_1_2[2143:2136]} - {1'b0, layer_0_2[2143:2136]};
      mid_0[0] = {1'b0,layer_2_0[2127:2120]} - {1'b0, layer_1_0[2127:2120]};
      mid_0[1] = {1'b0,layer_2_0[2135:2128]} - {1'b0, layer_1_0[2135:2128]};
      mid_0[2] = {1'b0,layer_2_0[2143:2136]} - {1'b0, layer_1_0[2143:2136]};
      mid_1[0] = {1'b0,layer_2_1[2127:2120]} - {1'b0, layer_1_1[2127:2120]};
      mid_1[1] = {1'b0,layer_2_1[2135:2128]} - {1'b0, layer_1_1[2135:2128]};
      mid_1[2] = {1'b0,layer_2_1[2143:2136]} - {1'b0, layer_1_1[2143:2136]};
      mid_2[0] = {1'b0,layer_2_2[2127:2120]} - {1'b0, layer_1_2[2127:2120]};
      mid_2[1] = {1'b0,layer_2_2[2135:2128]} - {1'b0, layer_1_2[2135:2128]};
      mid_2[2] = {1'b0,layer_2_2[2143:2136]} - {1'b0, layer_1_2[2143:2136]};
      btm_0[0] = {1'b0,layer_3_0[2127:2120]} - {1'b0, layer_2_0[2127:2120]};
      btm_0[1] = {1'b0,layer_3_0[2135:2128]} - {1'b0, layer_2_0[2135:2128]};
      btm_0[2] = {1'b0,layer_3_0[2143:2136]} - {1'b0, layer_2_0[2143:2136]};
      btm_1[0] = {1'b0,layer_3_1[2127:2120]} - {1'b0, layer_2_1[2127:2120]};
      btm_1[1] = {1'b0,layer_3_1[2135:2128]} - {1'b0, layer_2_1[2135:2128]};
      btm_1[2] = {1'b0,layer_3_1[2143:2136]} - {1'b0, layer_2_1[2143:2136]};
      btm_2[0] = {1'b0,layer_3_2[2127:2120]} - {1'b0, layer_2_2[2127:2120]};
      btm_2[1] = {1'b0,layer_3_2[2135:2128]} - {1'b0, layer_2_2[2135:2128]};
      btm_2[2] = {1'b0,layer_3_2[2143:2136]} - {1'b0, layer_2_2[2143:2136]};
    end
    'd267: begin
      top_0[0] = {1'b0,layer_1_0[2135:2128]} - {1'b0, layer_0_0[2135:2128]};
      top_0[1] = {1'b0,layer_1_0[2143:2136]} - {1'b0, layer_0_0[2143:2136]};
      top_0[2] = {1'b0,layer_1_0[2151:2144]} - {1'b0, layer_0_0[2151:2144]};
      top_1[0] = {1'b0,layer_1_1[2135:2128]} - {1'b0, layer_0_1[2135:2128]};
      top_1[1] = {1'b0,layer_1_1[2143:2136]} - {1'b0, layer_0_1[2143:2136]};
      top_1[2] = {1'b0,layer_1_1[2151:2144]} - {1'b0, layer_0_1[2151:2144]};
      top_2[0] = {1'b0,layer_1_2[2135:2128]} - {1'b0, layer_0_2[2135:2128]};
      top_2[1] = {1'b0,layer_1_2[2143:2136]} - {1'b0, layer_0_2[2143:2136]};
      top_2[2] = {1'b0,layer_1_2[2151:2144]} - {1'b0, layer_0_2[2151:2144]};
      mid_0[0] = {1'b0,layer_2_0[2135:2128]} - {1'b0, layer_1_0[2135:2128]};
      mid_0[1] = {1'b0,layer_2_0[2143:2136]} - {1'b0, layer_1_0[2143:2136]};
      mid_0[2] = {1'b0,layer_2_0[2151:2144]} - {1'b0, layer_1_0[2151:2144]};
      mid_1[0] = {1'b0,layer_2_1[2135:2128]} - {1'b0, layer_1_1[2135:2128]};
      mid_1[1] = {1'b0,layer_2_1[2143:2136]} - {1'b0, layer_1_1[2143:2136]};
      mid_1[2] = {1'b0,layer_2_1[2151:2144]} - {1'b0, layer_1_1[2151:2144]};
      mid_2[0] = {1'b0,layer_2_2[2135:2128]} - {1'b0, layer_1_2[2135:2128]};
      mid_2[1] = {1'b0,layer_2_2[2143:2136]} - {1'b0, layer_1_2[2143:2136]};
      mid_2[2] = {1'b0,layer_2_2[2151:2144]} - {1'b0, layer_1_2[2151:2144]};
      btm_0[0] = {1'b0,layer_3_0[2135:2128]} - {1'b0, layer_2_0[2135:2128]};
      btm_0[1] = {1'b0,layer_3_0[2143:2136]} - {1'b0, layer_2_0[2143:2136]};
      btm_0[2] = {1'b0,layer_3_0[2151:2144]} - {1'b0, layer_2_0[2151:2144]};
      btm_1[0] = {1'b0,layer_3_1[2135:2128]} - {1'b0, layer_2_1[2135:2128]};
      btm_1[1] = {1'b0,layer_3_1[2143:2136]} - {1'b0, layer_2_1[2143:2136]};
      btm_1[2] = {1'b0,layer_3_1[2151:2144]} - {1'b0, layer_2_1[2151:2144]};
      btm_2[0] = {1'b0,layer_3_2[2135:2128]} - {1'b0, layer_2_2[2135:2128]};
      btm_2[1] = {1'b0,layer_3_2[2143:2136]} - {1'b0, layer_2_2[2143:2136]};
      btm_2[2] = {1'b0,layer_3_2[2151:2144]} - {1'b0, layer_2_2[2151:2144]};
    end
    'd268: begin
      top_0[0] = {1'b0,layer_1_0[2143:2136]} - {1'b0, layer_0_0[2143:2136]};
      top_0[1] = {1'b0,layer_1_0[2151:2144]} - {1'b0, layer_0_0[2151:2144]};
      top_0[2] = {1'b0,layer_1_0[2159:2152]} - {1'b0, layer_0_0[2159:2152]};
      top_1[0] = {1'b0,layer_1_1[2143:2136]} - {1'b0, layer_0_1[2143:2136]};
      top_1[1] = {1'b0,layer_1_1[2151:2144]} - {1'b0, layer_0_1[2151:2144]};
      top_1[2] = {1'b0,layer_1_1[2159:2152]} - {1'b0, layer_0_1[2159:2152]};
      top_2[0] = {1'b0,layer_1_2[2143:2136]} - {1'b0, layer_0_2[2143:2136]};
      top_2[1] = {1'b0,layer_1_2[2151:2144]} - {1'b0, layer_0_2[2151:2144]};
      top_2[2] = {1'b0,layer_1_2[2159:2152]} - {1'b0, layer_0_2[2159:2152]};
      mid_0[0] = {1'b0,layer_2_0[2143:2136]} - {1'b0, layer_1_0[2143:2136]};
      mid_0[1] = {1'b0,layer_2_0[2151:2144]} - {1'b0, layer_1_0[2151:2144]};
      mid_0[2] = {1'b0,layer_2_0[2159:2152]} - {1'b0, layer_1_0[2159:2152]};
      mid_1[0] = {1'b0,layer_2_1[2143:2136]} - {1'b0, layer_1_1[2143:2136]};
      mid_1[1] = {1'b0,layer_2_1[2151:2144]} - {1'b0, layer_1_1[2151:2144]};
      mid_1[2] = {1'b0,layer_2_1[2159:2152]} - {1'b0, layer_1_1[2159:2152]};
      mid_2[0] = {1'b0,layer_2_2[2143:2136]} - {1'b0, layer_1_2[2143:2136]};
      mid_2[1] = {1'b0,layer_2_2[2151:2144]} - {1'b0, layer_1_2[2151:2144]};
      mid_2[2] = {1'b0,layer_2_2[2159:2152]} - {1'b0, layer_1_2[2159:2152]};
      btm_0[0] = {1'b0,layer_3_0[2143:2136]} - {1'b0, layer_2_0[2143:2136]};
      btm_0[1] = {1'b0,layer_3_0[2151:2144]} - {1'b0, layer_2_0[2151:2144]};
      btm_0[2] = {1'b0,layer_3_0[2159:2152]} - {1'b0, layer_2_0[2159:2152]};
      btm_1[0] = {1'b0,layer_3_1[2143:2136]} - {1'b0, layer_2_1[2143:2136]};
      btm_1[1] = {1'b0,layer_3_1[2151:2144]} - {1'b0, layer_2_1[2151:2144]};
      btm_1[2] = {1'b0,layer_3_1[2159:2152]} - {1'b0, layer_2_1[2159:2152]};
      btm_2[0] = {1'b0,layer_3_2[2143:2136]} - {1'b0, layer_2_2[2143:2136]};
      btm_2[1] = {1'b0,layer_3_2[2151:2144]} - {1'b0, layer_2_2[2151:2144]};
      btm_2[2] = {1'b0,layer_3_2[2159:2152]} - {1'b0, layer_2_2[2159:2152]};
    end
    'd269: begin
      top_0[0] = {1'b0,layer_1_0[2151:2144]} - {1'b0, layer_0_0[2151:2144]};
      top_0[1] = {1'b0,layer_1_0[2159:2152]} - {1'b0, layer_0_0[2159:2152]};
      top_0[2] = {1'b0,layer_1_0[2167:2160]} - {1'b0, layer_0_0[2167:2160]};
      top_1[0] = {1'b0,layer_1_1[2151:2144]} - {1'b0, layer_0_1[2151:2144]};
      top_1[1] = {1'b0,layer_1_1[2159:2152]} - {1'b0, layer_0_1[2159:2152]};
      top_1[2] = {1'b0,layer_1_1[2167:2160]} - {1'b0, layer_0_1[2167:2160]};
      top_2[0] = {1'b0,layer_1_2[2151:2144]} - {1'b0, layer_0_2[2151:2144]};
      top_2[1] = {1'b0,layer_1_2[2159:2152]} - {1'b0, layer_0_2[2159:2152]};
      top_2[2] = {1'b0,layer_1_2[2167:2160]} - {1'b0, layer_0_2[2167:2160]};
      mid_0[0] = {1'b0,layer_2_0[2151:2144]} - {1'b0, layer_1_0[2151:2144]};
      mid_0[1] = {1'b0,layer_2_0[2159:2152]} - {1'b0, layer_1_0[2159:2152]};
      mid_0[2] = {1'b0,layer_2_0[2167:2160]} - {1'b0, layer_1_0[2167:2160]};
      mid_1[0] = {1'b0,layer_2_1[2151:2144]} - {1'b0, layer_1_1[2151:2144]};
      mid_1[1] = {1'b0,layer_2_1[2159:2152]} - {1'b0, layer_1_1[2159:2152]};
      mid_1[2] = {1'b0,layer_2_1[2167:2160]} - {1'b0, layer_1_1[2167:2160]};
      mid_2[0] = {1'b0,layer_2_2[2151:2144]} - {1'b0, layer_1_2[2151:2144]};
      mid_2[1] = {1'b0,layer_2_2[2159:2152]} - {1'b0, layer_1_2[2159:2152]};
      mid_2[2] = {1'b0,layer_2_2[2167:2160]} - {1'b0, layer_1_2[2167:2160]};
      btm_0[0] = {1'b0,layer_3_0[2151:2144]} - {1'b0, layer_2_0[2151:2144]};
      btm_0[1] = {1'b0,layer_3_0[2159:2152]} - {1'b0, layer_2_0[2159:2152]};
      btm_0[2] = {1'b0,layer_3_0[2167:2160]} - {1'b0, layer_2_0[2167:2160]};
      btm_1[0] = {1'b0,layer_3_1[2151:2144]} - {1'b0, layer_2_1[2151:2144]};
      btm_1[1] = {1'b0,layer_3_1[2159:2152]} - {1'b0, layer_2_1[2159:2152]};
      btm_1[2] = {1'b0,layer_3_1[2167:2160]} - {1'b0, layer_2_1[2167:2160]};
      btm_2[0] = {1'b0,layer_3_2[2151:2144]} - {1'b0, layer_2_2[2151:2144]};
      btm_2[1] = {1'b0,layer_3_2[2159:2152]} - {1'b0, layer_2_2[2159:2152]};
      btm_2[2] = {1'b0,layer_3_2[2167:2160]} - {1'b0, layer_2_2[2167:2160]};
    end
    'd270: begin
      top_0[0] = {1'b0,layer_1_0[2159:2152]} - {1'b0, layer_0_0[2159:2152]};
      top_0[1] = {1'b0,layer_1_0[2167:2160]} - {1'b0, layer_0_0[2167:2160]};
      top_0[2] = {1'b0,layer_1_0[2175:2168]} - {1'b0, layer_0_0[2175:2168]};
      top_1[0] = {1'b0,layer_1_1[2159:2152]} - {1'b0, layer_0_1[2159:2152]};
      top_1[1] = {1'b0,layer_1_1[2167:2160]} - {1'b0, layer_0_1[2167:2160]};
      top_1[2] = {1'b0,layer_1_1[2175:2168]} - {1'b0, layer_0_1[2175:2168]};
      top_2[0] = {1'b0,layer_1_2[2159:2152]} - {1'b0, layer_0_2[2159:2152]};
      top_2[1] = {1'b0,layer_1_2[2167:2160]} - {1'b0, layer_0_2[2167:2160]};
      top_2[2] = {1'b0,layer_1_2[2175:2168]} - {1'b0, layer_0_2[2175:2168]};
      mid_0[0] = {1'b0,layer_2_0[2159:2152]} - {1'b0, layer_1_0[2159:2152]};
      mid_0[1] = {1'b0,layer_2_0[2167:2160]} - {1'b0, layer_1_0[2167:2160]};
      mid_0[2] = {1'b0,layer_2_0[2175:2168]} - {1'b0, layer_1_0[2175:2168]};
      mid_1[0] = {1'b0,layer_2_1[2159:2152]} - {1'b0, layer_1_1[2159:2152]};
      mid_1[1] = {1'b0,layer_2_1[2167:2160]} - {1'b0, layer_1_1[2167:2160]};
      mid_1[2] = {1'b0,layer_2_1[2175:2168]} - {1'b0, layer_1_1[2175:2168]};
      mid_2[0] = {1'b0,layer_2_2[2159:2152]} - {1'b0, layer_1_2[2159:2152]};
      mid_2[1] = {1'b0,layer_2_2[2167:2160]} - {1'b0, layer_1_2[2167:2160]};
      mid_2[2] = {1'b0,layer_2_2[2175:2168]} - {1'b0, layer_1_2[2175:2168]};
      btm_0[0] = {1'b0,layer_3_0[2159:2152]} - {1'b0, layer_2_0[2159:2152]};
      btm_0[1] = {1'b0,layer_3_0[2167:2160]} - {1'b0, layer_2_0[2167:2160]};
      btm_0[2] = {1'b0,layer_3_0[2175:2168]} - {1'b0, layer_2_0[2175:2168]};
      btm_1[0] = {1'b0,layer_3_1[2159:2152]} - {1'b0, layer_2_1[2159:2152]};
      btm_1[1] = {1'b0,layer_3_1[2167:2160]} - {1'b0, layer_2_1[2167:2160]};
      btm_1[2] = {1'b0,layer_3_1[2175:2168]} - {1'b0, layer_2_1[2175:2168]};
      btm_2[0] = {1'b0,layer_3_2[2159:2152]} - {1'b0, layer_2_2[2159:2152]};
      btm_2[1] = {1'b0,layer_3_2[2167:2160]} - {1'b0, layer_2_2[2167:2160]};
      btm_2[2] = {1'b0,layer_3_2[2175:2168]} - {1'b0, layer_2_2[2175:2168]};
    end
    'd271: begin
      top_0[0] = {1'b0,layer_1_0[2167:2160]} - {1'b0, layer_0_0[2167:2160]};
      top_0[1] = {1'b0,layer_1_0[2175:2168]} - {1'b0, layer_0_0[2175:2168]};
      top_0[2] = {1'b0,layer_1_0[2183:2176]} - {1'b0, layer_0_0[2183:2176]};
      top_1[0] = {1'b0,layer_1_1[2167:2160]} - {1'b0, layer_0_1[2167:2160]};
      top_1[1] = {1'b0,layer_1_1[2175:2168]} - {1'b0, layer_0_1[2175:2168]};
      top_1[2] = {1'b0,layer_1_1[2183:2176]} - {1'b0, layer_0_1[2183:2176]};
      top_2[0] = {1'b0,layer_1_2[2167:2160]} - {1'b0, layer_0_2[2167:2160]};
      top_2[1] = {1'b0,layer_1_2[2175:2168]} - {1'b0, layer_0_2[2175:2168]};
      top_2[2] = {1'b0,layer_1_2[2183:2176]} - {1'b0, layer_0_2[2183:2176]};
      mid_0[0] = {1'b0,layer_2_0[2167:2160]} - {1'b0, layer_1_0[2167:2160]};
      mid_0[1] = {1'b0,layer_2_0[2175:2168]} - {1'b0, layer_1_0[2175:2168]};
      mid_0[2] = {1'b0,layer_2_0[2183:2176]} - {1'b0, layer_1_0[2183:2176]};
      mid_1[0] = {1'b0,layer_2_1[2167:2160]} - {1'b0, layer_1_1[2167:2160]};
      mid_1[1] = {1'b0,layer_2_1[2175:2168]} - {1'b0, layer_1_1[2175:2168]};
      mid_1[2] = {1'b0,layer_2_1[2183:2176]} - {1'b0, layer_1_1[2183:2176]};
      mid_2[0] = {1'b0,layer_2_2[2167:2160]} - {1'b0, layer_1_2[2167:2160]};
      mid_2[1] = {1'b0,layer_2_2[2175:2168]} - {1'b0, layer_1_2[2175:2168]};
      mid_2[2] = {1'b0,layer_2_2[2183:2176]} - {1'b0, layer_1_2[2183:2176]};
      btm_0[0] = {1'b0,layer_3_0[2167:2160]} - {1'b0, layer_2_0[2167:2160]};
      btm_0[1] = {1'b0,layer_3_0[2175:2168]} - {1'b0, layer_2_0[2175:2168]};
      btm_0[2] = {1'b0,layer_3_0[2183:2176]} - {1'b0, layer_2_0[2183:2176]};
      btm_1[0] = {1'b0,layer_3_1[2167:2160]} - {1'b0, layer_2_1[2167:2160]};
      btm_1[1] = {1'b0,layer_3_1[2175:2168]} - {1'b0, layer_2_1[2175:2168]};
      btm_1[2] = {1'b0,layer_3_1[2183:2176]} - {1'b0, layer_2_1[2183:2176]};
      btm_2[0] = {1'b0,layer_3_2[2167:2160]} - {1'b0, layer_2_2[2167:2160]};
      btm_2[1] = {1'b0,layer_3_2[2175:2168]} - {1'b0, layer_2_2[2175:2168]};
      btm_2[2] = {1'b0,layer_3_2[2183:2176]} - {1'b0, layer_2_2[2183:2176]};
    end
    'd272: begin
      top_0[0] = {1'b0,layer_1_0[2175:2168]} - {1'b0, layer_0_0[2175:2168]};
      top_0[1] = {1'b0,layer_1_0[2183:2176]} - {1'b0, layer_0_0[2183:2176]};
      top_0[2] = {1'b0,layer_1_0[2191:2184]} - {1'b0, layer_0_0[2191:2184]};
      top_1[0] = {1'b0,layer_1_1[2175:2168]} - {1'b0, layer_0_1[2175:2168]};
      top_1[1] = {1'b0,layer_1_1[2183:2176]} - {1'b0, layer_0_1[2183:2176]};
      top_1[2] = {1'b0,layer_1_1[2191:2184]} - {1'b0, layer_0_1[2191:2184]};
      top_2[0] = {1'b0,layer_1_2[2175:2168]} - {1'b0, layer_0_2[2175:2168]};
      top_2[1] = {1'b0,layer_1_2[2183:2176]} - {1'b0, layer_0_2[2183:2176]};
      top_2[2] = {1'b0,layer_1_2[2191:2184]} - {1'b0, layer_0_2[2191:2184]};
      mid_0[0] = {1'b0,layer_2_0[2175:2168]} - {1'b0, layer_1_0[2175:2168]};
      mid_0[1] = {1'b0,layer_2_0[2183:2176]} - {1'b0, layer_1_0[2183:2176]};
      mid_0[2] = {1'b0,layer_2_0[2191:2184]} - {1'b0, layer_1_0[2191:2184]};
      mid_1[0] = {1'b0,layer_2_1[2175:2168]} - {1'b0, layer_1_1[2175:2168]};
      mid_1[1] = {1'b0,layer_2_1[2183:2176]} - {1'b0, layer_1_1[2183:2176]};
      mid_1[2] = {1'b0,layer_2_1[2191:2184]} - {1'b0, layer_1_1[2191:2184]};
      mid_2[0] = {1'b0,layer_2_2[2175:2168]} - {1'b0, layer_1_2[2175:2168]};
      mid_2[1] = {1'b0,layer_2_2[2183:2176]} - {1'b0, layer_1_2[2183:2176]};
      mid_2[2] = {1'b0,layer_2_2[2191:2184]} - {1'b0, layer_1_2[2191:2184]};
      btm_0[0] = {1'b0,layer_3_0[2175:2168]} - {1'b0, layer_2_0[2175:2168]};
      btm_0[1] = {1'b0,layer_3_0[2183:2176]} - {1'b0, layer_2_0[2183:2176]};
      btm_0[2] = {1'b0,layer_3_0[2191:2184]} - {1'b0, layer_2_0[2191:2184]};
      btm_1[0] = {1'b0,layer_3_1[2175:2168]} - {1'b0, layer_2_1[2175:2168]};
      btm_1[1] = {1'b0,layer_3_1[2183:2176]} - {1'b0, layer_2_1[2183:2176]};
      btm_1[2] = {1'b0,layer_3_1[2191:2184]} - {1'b0, layer_2_1[2191:2184]};
      btm_2[0] = {1'b0,layer_3_2[2175:2168]} - {1'b0, layer_2_2[2175:2168]};
      btm_2[1] = {1'b0,layer_3_2[2183:2176]} - {1'b0, layer_2_2[2183:2176]};
      btm_2[2] = {1'b0,layer_3_2[2191:2184]} - {1'b0, layer_2_2[2191:2184]};
    end
    'd273: begin
      top_0[0] = {1'b0,layer_1_0[2183:2176]} - {1'b0, layer_0_0[2183:2176]};
      top_0[1] = {1'b0,layer_1_0[2191:2184]} - {1'b0, layer_0_0[2191:2184]};
      top_0[2] = {1'b0,layer_1_0[2199:2192]} - {1'b0, layer_0_0[2199:2192]};
      top_1[0] = {1'b0,layer_1_1[2183:2176]} - {1'b0, layer_0_1[2183:2176]};
      top_1[1] = {1'b0,layer_1_1[2191:2184]} - {1'b0, layer_0_1[2191:2184]};
      top_1[2] = {1'b0,layer_1_1[2199:2192]} - {1'b0, layer_0_1[2199:2192]};
      top_2[0] = {1'b0,layer_1_2[2183:2176]} - {1'b0, layer_0_2[2183:2176]};
      top_2[1] = {1'b0,layer_1_2[2191:2184]} - {1'b0, layer_0_2[2191:2184]};
      top_2[2] = {1'b0,layer_1_2[2199:2192]} - {1'b0, layer_0_2[2199:2192]};
      mid_0[0] = {1'b0,layer_2_0[2183:2176]} - {1'b0, layer_1_0[2183:2176]};
      mid_0[1] = {1'b0,layer_2_0[2191:2184]} - {1'b0, layer_1_0[2191:2184]};
      mid_0[2] = {1'b0,layer_2_0[2199:2192]} - {1'b0, layer_1_0[2199:2192]};
      mid_1[0] = {1'b0,layer_2_1[2183:2176]} - {1'b0, layer_1_1[2183:2176]};
      mid_1[1] = {1'b0,layer_2_1[2191:2184]} - {1'b0, layer_1_1[2191:2184]};
      mid_1[2] = {1'b0,layer_2_1[2199:2192]} - {1'b0, layer_1_1[2199:2192]};
      mid_2[0] = {1'b0,layer_2_2[2183:2176]} - {1'b0, layer_1_2[2183:2176]};
      mid_2[1] = {1'b0,layer_2_2[2191:2184]} - {1'b0, layer_1_2[2191:2184]};
      mid_2[2] = {1'b0,layer_2_2[2199:2192]} - {1'b0, layer_1_2[2199:2192]};
      btm_0[0] = {1'b0,layer_3_0[2183:2176]} - {1'b0, layer_2_0[2183:2176]};
      btm_0[1] = {1'b0,layer_3_0[2191:2184]} - {1'b0, layer_2_0[2191:2184]};
      btm_0[2] = {1'b0,layer_3_0[2199:2192]} - {1'b0, layer_2_0[2199:2192]};
      btm_1[0] = {1'b0,layer_3_1[2183:2176]} - {1'b0, layer_2_1[2183:2176]};
      btm_1[1] = {1'b0,layer_3_1[2191:2184]} - {1'b0, layer_2_1[2191:2184]};
      btm_1[2] = {1'b0,layer_3_1[2199:2192]} - {1'b0, layer_2_1[2199:2192]};
      btm_2[0] = {1'b0,layer_3_2[2183:2176]} - {1'b0, layer_2_2[2183:2176]};
      btm_2[1] = {1'b0,layer_3_2[2191:2184]} - {1'b0, layer_2_2[2191:2184]};
      btm_2[2] = {1'b0,layer_3_2[2199:2192]} - {1'b0, layer_2_2[2199:2192]};
    end
    'd274: begin
      top_0[0] = {1'b0,layer_1_0[2191:2184]} - {1'b0, layer_0_0[2191:2184]};
      top_0[1] = {1'b0,layer_1_0[2199:2192]} - {1'b0, layer_0_0[2199:2192]};
      top_0[2] = {1'b0,layer_1_0[2207:2200]} - {1'b0, layer_0_0[2207:2200]};
      top_1[0] = {1'b0,layer_1_1[2191:2184]} - {1'b0, layer_0_1[2191:2184]};
      top_1[1] = {1'b0,layer_1_1[2199:2192]} - {1'b0, layer_0_1[2199:2192]};
      top_1[2] = {1'b0,layer_1_1[2207:2200]} - {1'b0, layer_0_1[2207:2200]};
      top_2[0] = {1'b0,layer_1_2[2191:2184]} - {1'b0, layer_0_2[2191:2184]};
      top_2[1] = {1'b0,layer_1_2[2199:2192]} - {1'b0, layer_0_2[2199:2192]};
      top_2[2] = {1'b0,layer_1_2[2207:2200]} - {1'b0, layer_0_2[2207:2200]};
      mid_0[0] = {1'b0,layer_2_0[2191:2184]} - {1'b0, layer_1_0[2191:2184]};
      mid_0[1] = {1'b0,layer_2_0[2199:2192]} - {1'b0, layer_1_0[2199:2192]};
      mid_0[2] = {1'b0,layer_2_0[2207:2200]} - {1'b0, layer_1_0[2207:2200]};
      mid_1[0] = {1'b0,layer_2_1[2191:2184]} - {1'b0, layer_1_1[2191:2184]};
      mid_1[1] = {1'b0,layer_2_1[2199:2192]} - {1'b0, layer_1_1[2199:2192]};
      mid_1[2] = {1'b0,layer_2_1[2207:2200]} - {1'b0, layer_1_1[2207:2200]};
      mid_2[0] = {1'b0,layer_2_2[2191:2184]} - {1'b0, layer_1_2[2191:2184]};
      mid_2[1] = {1'b0,layer_2_2[2199:2192]} - {1'b0, layer_1_2[2199:2192]};
      mid_2[2] = {1'b0,layer_2_2[2207:2200]} - {1'b0, layer_1_2[2207:2200]};
      btm_0[0] = {1'b0,layer_3_0[2191:2184]} - {1'b0, layer_2_0[2191:2184]};
      btm_0[1] = {1'b0,layer_3_0[2199:2192]} - {1'b0, layer_2_0[2199:2192]};
      btm_0[2] = {1'b0,layer_3_0[2207:2200]} - {1'b0, layer_2_0[2207:2200]};
      btm_1[0] = {1'b0,layer_3_1[2191:2184]} - {1'b0, layer_2_1[2191:2184]};
      btm_1[1] = {1'b0,layer_3_1[2199:2192]} - {1'b0, layer_2_1[2199:2192]};
      btm_1[2] = {1'b0,layer_3_1[2207:2200]} - {1'b0, layer_2_1[2207:2200]};
      btm_2[0] = {1'b0,layer_3_2[2191:2184]} - {1'b0, layer_2_2[2191:2184]};
      btm_2[1] = {1'b0,layer_3_2[2199:2192]} - {1'b0, layer_2_2[2199:2192]};
      btm_2[2] = {1'b0,layer_3_2[2207:2200]} - {1'b0, layer_2_2[2207:2200]};
    end
    'd275: begin
      top_0[0] = {1'b0,layer_1_0[2199:2192]} - {1'b0, layer_0_0[2199:2192]};
      top_0[1] = {1'b0,layer_1_0[2207:2200]} - {1'b0, layer_0_0[2207:2200]};
      top_0[2] = {1'b0,layer_1_0[2215:2208]} - {1'b0, layer_0_0[2215:2208]};
      top_1[0] = {1'b0,layer_1_1[2199:2192]} - {1'b0, layer_0_1[2199:2192]};
      top_1[1] = {1'b0,layer_1_1[2207:2200]} - {1'b0, layer_0_1[2207:2200]};
      top_1[2] = {1'b0,layer_1_1[2215:2208]} - {1'b0, layer_0_1[2215:2208]};
      top_2[0] = {1'b0,layer_1_2[2199:2192]} - {1'b0, layer_0_2[2199:2192]};
      top_2[1] = {1'b0,layer_1_2[2207:2200]} - {1'b0, layer_0_2[2207:2200]};
      top_2[2] = {1'b0,layer_1_2[2215:2208]} - {1'b0, layer_0_2[2215:2208]};
      mid_0[0] = {1'b0,layer_2_0[2199:2192]} - {1'b0, layer_1_0[2199:2192]};
      mid_0[1] = {1'b0,layer_2_0[2207:2200]} - {1'b0, layer_1_0[2207:2200]};
      mid_0[2] = {1'b0,layer_2_0[2215:2208]} - {1'b0, layer_1_0[2215:2208]};
      mid_1[0] = {1'b0,layer_2_1[2199:2192]} - {1'b0, layer_1_1[2199:2192]};
      mid_1[1] = {1'b0,layer_2_1[2207:2200]} - {1'b0, layer_1_1[2207:2200]};
      mid_1[2] = {1'b0,layer_2_1[2215:2208]} - {1'b0, layer_1_1[2215:2208]};
      mid_2[0] = {1'b0,layer_2_2[2199:2192]} - {1'b0, layer_1_2[2199:2192]};
      mid_2[1] = {1'b0,layer_2_2[2207:2200]} - {1'b0, layer_1_2[2207:2200]};
      mid_2[2] = {1'b0,layer_2_2[2215:2208]} - {1'b0, layer_1_2[2215:2208]};
      btm_0[0] = {1'b0,layer_3_0[2199:2192]} - {1'b0, layer_2_0[2199:2192]};
      btm_0[1] = {1'b0,layer_3_0[2207:2200]} - {1'b0, layer_2_0[2207:2200]};
      btm_0[2] = {1'b0,layer_3_0[2215:2208]} - {1'b0, layer_2_0[2215:2208]};
      btm_1[0] = {1'b0,layer_3_1[2199:2192]} - {1'b0, layer_2_1[2199:2192]};
      btm_1[1] = {1'b0,layer_3_1[2207:2200]} - {1'b0, layer_2_1[2207:2200]};
      btm_1[2] = {1'b0,layer_3_1[2215:2208]} - {1'b0, layer_2_1[2215:2208]};
      btm_2[0] = {1'b0,layer_3_2[2199:2192]} - {1'b0, layer_2_2[2199:2192]};
      btm_2[1] = {1'b0,layer_3_2[2207:2200]} - {1'b0, layer_2_2[2207:2200]};
      btm_2[2] = {1'b0,layer_3_2[2215:2208]} - {1'b0, layer_2_2[2215:2208]};
    end
    'd276: begin
      top_0[0] = {1'b0,layer_1_0[2207:2200]} - {1'b0, layer_0_0[2207:2200]};
      top_0[1] = {1'b0,layer_1_0[2215:2208]} - {1'b0, layer_0_0[2215:2208]};
      top_0[2] = {1'b0,layer_1_0[2223:2216]} - {1'b0, layer_0_0[2223:2216]};
      top_1[0] = {1'b0,layer_1_1[2207:2200]} - {1'b0, layer_0_1[2207:2200]};
      top_1[1] = {1'b0,layer_1_1[2215:2208]} - {1'b0, layer_0_1[2215:2208]};
      top_1[2] = {1'b0,layer_1_1[2223:2216]} - {1'b0, layer_0_1[2223:2216]};
      top_2[0] = {1'b0,layer_1_2[2207:2200]} - {1'b0, layer_0_2[2207:2200]};
      top_2[1] = {1'b0,layer_1_2[2215:2208]} - {1'b0, layer_0_2[2215:2208]};
      top_2[2] = {1'b0,layer_1_2[2223:2216]} - {1'b0, layer_0_2[2223:2216]};
      mid_0[0] = {1'b0,layer_2_0[2207:2200]} - {1'b0, layer_1_0[2207:2200]};
      mid_0[1] = {1'b0,layer_2_0[2215:2208]} - {1'b0, layer_1_0[2215:2208]};
      mid_0[2] = {1'b0,layer_2_0[2223:2216]} - {1'b0, layer_1_0[2223:2216]};
      mid_1[0] = {1'b0,layer_2_1[2207:2200]} - {1'b0, layer_1_1[2207:2200]};
      mid_1[1] = {1'b0,layer_2_1[2215:2208]} - {1'b0, layer_1_1[2215:2208]};
      mid_1[2] = {1'b0,layer_2_1[2223:2216]} - {1'b0, layer_1_1[2223:2216]};
      mid_2[0] = {1'b0,layer_2_2[2207:2200]} - {1'b0, layer_1_2[2207:2200]};
      mid_2[1] = {1'b0,layer_2_2[2215:2208]} - {1'b0, layer_1_2[2215:2208]};
      mid_2[2] = {1'b0,layer_2_2[2223:2216]} - {1'b0, layer_1_2[2223:2216]};
      btm_0[0] = {1'b0,layer_3_0[2207:2200]} - {1'b0, layer_2_0[2207:2200]};
      btm_0[1] = {1'b0,layer_3_0[2215:2208]} - {1'b0, layer_2_0[2215:2208]};
      btm_0[2] = {1'b0,layer_3_0[2223:2216]} - {1'b0, layer_2_0[2223:2216]};
      btm_1[0] = {1'b0,layer_3_1[2207:2200]} - {1'b0, layer_2_1[2207:2200]};
      btm_1[1] = {1'b0,layer_3_1[2215:2208]} - {1'b0, layer_2_1[2215:2208]};
      btm_1[2] = {1'b0,layer_3_1[2223:2216]} - {1'b0, layer_2_1[2223:2216]};
      btm_2[0] = {1'b0,layer_3_2[2207:2200]} - {1'b0, layer_2_2[2207:2200]};
      btm_2[1] = {1'b0,layer_3_2[2215:2208]} - {1'b0, layer_2_2[2215:2208]};
      btm_2[2] = {1'b0,layer_3_2[2223:2216]} - {1'b0, layer_2_2[2223:2216]};
    end
    'd277: begin
      top_0[0] = {1'b0,layer_1_0[2215:2208]} - {1'b0, layer_0_0[2215:2208]};
      top_0[1] = {1'b0,layer_1_0[2223:2216]} - {1'b0, layer_0_0[2223:2216]};
      top_0[2] = {1'b0,layer_1_0[2231:2224]} - {1'b0, layer_0_0[2231:2224]};
      top_1[0] = {1'b0,layer_1_1[2215:2208]} - {1'b0, layer_0_1[2215:2208]};
      top_1[1] = {1'b0,layer_1_1[2223:2216]} - {1'b0, layer_0_1[2223:2216]};
      top_1[2] = {1'b0,layer_1_1[2231:2224]} - {1'b0, layer_0_1[2231:2224]};
      top_2[0] = {1'b0,layer_1_2[2215:2208]} - {1'b0, layer_0_2[2215:2208]};
      top_2[1] = {1'b0,layer_1_2[2223:2216]} - {1'b0, layer_0_2[2223:2216]};
      top_2[2] = {1'b0,layer_1_2[2231:2224]} - {1'b0, layer_0_2[2231:2224]};
      mid_0[0] = {1'b0,layer_2_0[2215:2208]} - {1'b0, layer_1_0[2215:2208]};
      mid_0[1] = {1'b0,layer_2_0[2223:2216]} - {1'b0, layer_1_0[2223:2216]};
      mid_0[2] = {1'b0,layer_2_0[2231:2224]} - {1'b0, layer_1_0[2231:2224]};
      mid_1[0] = {1'b0,layer_2_1[2215:2208]} - {1'b0, layer_1_1[2215:2208]};
      mid_1[1] = {1'b0,layer_2_1[2223:2216]} - {1'b0, layer_1_1[2223:2216]};
      mid_1[2] = {1'b0,layer_2_1[2231:2224]} - {1'b0, layer_1_1[2231:2224]};
      mid_2[0] = {1'b0,layer_2_2[2215:2208]} - {1'b0, layer_1_2[2215:2208]};
      mid_2[1] = {1'b0,layer_2_2[2223:2216]} - {1'b0, layer_1_2[2223:2216]};
      mid_2[2] = {1'b0,layer_2_2[2231:2224]} - {1'b0, layer_1_2[2231:2224]};
      btm_0[0] = {1'b0,layer_3_0[2215:2208]} - {1'b0, layer_2_0[2215:2208]};
      btm_0[1] = {1'b0,layer_3_0[2223:2216]} - {1'b0, layer_2_0[2223:2216]};
      btm_0[2] = {1'b0,layer_3_0[2231:2224]} - {1'b0, layer_2_0[2231:2224]};
      btm_1[0] = {1'b0,layer_3_1[2215:2208]} - {1'b0, layer_2_1[2215:2208]};
      btm_1[1] = {1'b0,layer_3_1[2223:2216]} - {1'b0, layer_2_1[2223:2216]};
      btm_1[2] = {1'b0,layer_3_1[2231:2224]} - {1'b0, layer_2_1[2231:2224]};
      btm_2[0] = {1'b0,layer_3_2[2215:2208]} - {1'b0, layer_2_2[2215:2208]};
      btm_2[1] = {1'b0,layer_3_2[2223:2216]} - {1'b0, layer_2_2[2223:2216]};
      btm_2[2] = {1'b0,layer_3_2[2231:2224]} - {1'b0, layer_2_2[2231:2224]};
    end
    'd278: begin
      top_0[0] = {1'b0,layer_1_0[2223:2216]} - {1'b0, layer_0_0[2223:2216]};
      top_0[1] = {1'b0,layer_1_0[2231:2224]} - {1'b0, layer_0_0[2231:2224]};
      top_0[2] = {1'b0,layer_1_0[2239:2232]} - {1'b0, layer_0_0[2239:2232]};
      top_1[0] = {1'b0,layer_1_1[2223:2216]} - {1'b0, layer_0_1[2223:2216]};
      top_1[1] = {1'b0,layer_1_1[2231:2224]} - {1'b0, layer_0_1[2231:2224]};
      top_1[2] = {1'b0,layer_1_1[2239:2232]} - {1'b0, layer_0_1[2239:2232]};
      top_2[0] = {1'b0,layer_1_2[2223:2216]} - {1'b0, layer_0_2[2223:2216]};
      top_2[1] = {1'b0,layer_1_2[2231:2224]} - {1'b0, layer_0_2[2231:2224]};
      top_2[2] = {1'b0,layer_1_2[2239:2232]} - {1'b0, layer_0_2[2239:2232]};
      mid_0[0] = {1'b0,layer_2_0[2223:2216]} - {1'b0, layer_1_0[2223:2216]};
      mid_0[1] = {1'b0,layer_2_0[2231:2224]} - {1'b0, layer_1_0[2231:2224]};
      mid_0[2] = {1'b0,layer_2_0[2239:2232]} - {1'b0, layer_1_0[2239:2232]};
      mid_1[0] = {1'b0,layer_2_1[2223:2216]} - {1'b0, layer_1_1[2223:2216]};
      mid_1[1] = {1'b0,layer_2_1[2231:2224]} - {1'b0, layer_1_1[2231:2224]};
      mid_1[2] = {1'b0,layer_2_1[2239:2232]} - {1'b0, layer_1_1[2239:2232]};
      mid_2[0] = {1'b0,layer_2_2[2223:2216]} - {1'b0, layer_1_2[2223:2216]};
      mid_2[1] = {1'b0,layer_2_2[2231:2224]} - {1'b0, layer_1_2[2231:2224]};
      mid_2[2] = {1'b0,layer_2_2[2239:2232]} - {1'b0, layer_1_2[2239:2232]};
      btm_0[0] = {1'b0,layer_3_0[2223:2216]} - {1'b0, layer_2_0[2223:2216]};
      btm_0[1] = {1'b0,layer_3_0[2231:2224]} - {1'b0, layer_2_0[2231:2224]};
      btm_0[2] = {1'b0,layer_3_0[2239:2232]} - {1'b0, layer_2_0[2239:2232]};
      btm_1[0] = {1'b0,layer_3_1[2223:2216]} - {1'b0, layer_2_1[2223:2216]};
      btm_1[1] = {1'b0,layer_3_1[2231:2224]} - {1'b0, layer_2_1[2231:2224]};
      btm_1[2] = {1'b0,layer_3_1[2239:2232]} - {1'b0, layer_2_1[2239:2232]};
      btm_2[0] = {1'b0,layer_3_2[2223:2216]} - {1'b0, layer_2_2[2223:2216]};
      btm_2[1] = {1'b0,layer_3_2[2231:2224]} - {1'b0, layer_2_2[2231:2224]};
      btm_2[2] = {1'b0,layer_3_2[2239:2232]} - {1'b0, layer_2_2[2239:2232]};
    end
    'd279: begin
      top_0[0] = {1'b0,layer_1_0[2231:2224]} - {1'b0, layer_0_0[2231:2224]};
      top_0[1] = {1'b0,layer_1_0[2239:2232]} - {1'b0, layer_0_0[2239:2232]};
      top_0[2] = {1'b0,layer_1_0[2247:2240]} - {1'b0, layer_0_0[2247:2240]};
      top_1[0] = {1'b0,layer_1_1[2231:2224]} - {1'b0, layer_0_1[2231:2224]};
      top_1[1] = {1'b0,layer_1_1[2239:2232]} - {1'b0, layer_0_1[2239:2232]};
      top_1[2] = {1'b0,layer_1_1[2247:2240]} - {1'b0, layer_0_1[2247:2240]};
      top_2[0] = {1'b0,layer_1_2[2231:2224]} - {1'b0, layer_0_2[2231:2224]};
      top_2[1] = {1'b0,layer_1_2[2239:2232]} - {1'b0, layer_0_2[2239:2232]};
      top_2[2] = {1'b0,layer_1_2[2247:2240]} - {1'b0, layer_0_2[2247:2240]};
      mid_0[0] = {1'b0,layer_2_0[2231:2224]} - {1'b0, layer_1_0[2231:2224]};
      mid_0[1] = {1'b0,layer_2_0[2239:2232]} - {1'b0, layer_1_0[2239:2232]};
      mid_0[2] = {1'b0,layer_2_0[2247:2240]} - {1'b0, layer_1_0[2247:2240]};
      mid_1[0] = {1'b0,layer_2_1[2231:2224]} - {1'b0, layer_1_1[2231:2224]};
      mid_1[1] = {1'b0,layer_2_1[2239:2232]} - {1'b0, layer_1_1[2239:2232]};
      mid_1[2] = {1'b0,layer_2_1[2247:2240]} - {1'b0, layer_1_1[2247:2240]};
      mid_2[0] = {1'b0,layer_2_2[2231:2224]} - {1'b0, layer_1_2[2231:2224]};
      mid_2[1] = {1'b0,layer_2_2[2239:2232]} - {1'b0, layer_1_2[2239:2232]};
      mid_2[2] = {1'b0,layer_2_2[2247:2240]} - {1'b0, layer_1_2[2247:2240]};
      btm_0[0] = {1'b0,layer_3_0[2231:2224]} - {1'b0, layer_2_0[2231:2224]};
      btm_0[1] = {1'b0,layer_3_0[2239:2232]} - {1'b0, layer_2_0[2239:2232]};
      btm_0[2] = {1'b0,layer_3_0[2247:2240]} - {1'b0, layer_2_0[2247:2240]};
      btm_1[0] = {1'b0,layer_3_1[2231:2224]} - {1'b0, layer_2_1[2231:2224]};
      btm_1[1] = {1'b0,layer_3_1[2239:2232]} - {1'b0, layer_2_1[2239:2232]};
      btm_1[2] = {1'b0,layer_3_1[2247:2240]} - {1'b0, layer_2_1[2247:2240]};
      btm_2[0] = {1'b0,layer_3_2[2231:2224]} - {1'b0, layer_2_2[2231:2224]};
      btm_2[1] = {1'b0,layer_3_2[2239:2232]} - {1'b0, layer_2_2[2239:2232]};
      btm_2[2] = {1'b0,layer_3_2[2247:2240]} - {1'b0, layer_2_2[2247:2240]};
    end
    'd280: begin
      top_0[0] = {1'b0,layer_1_0[2239:2232]} - {1'b0, layer_0_0[2239:2232]};
      top_0[1] = {1'b0,layer_1_0[2247:2240]} - {1'b0, layer_0_0[2247:2240]};
      top_0[2] = {1'b0,layer_1_0[2255:2248]} - {1'b0, layer_0_0[2255:2248]};
      top_1[0] = {1'b0,layer_1_1[2239:2232]} - {1'b0, layer_0_1[2239:2232]};
      top_1[1] = {1'b0,layer_1_1[2247:2240]} - {1'b0, layer_0_1[2247:2240]};
      top_1[2] = {1'b0,layer_1_1[2255:2248]} - {1'b0, layer_0_1[2255:2248]};
      top_2[0] = {1'b0,layer_1_2[2239:2232]} - {1'b0, layer_0_2[2239:2232]};
      top_2[1] = {1'b0,layer_1_2[2247:2240]} - {1'b0, layer_0_2[2247:2240]};
      top_2[2] = {1'b0,layer_1_2[2255:2248]} - {1'b0, layer_0_2[2255:2248]};
      mid_0[0] = {1'b0,layer_2_0[2239:2232]} - {1'b0, layer_1_0[2239:2232]};
      mid_0[1] = {1'b0,layer_2_0[2247:2240]} - {1'b0, layer_1_0[2247:2240]};
      mid_0[2] = {1'b0,layer_2_0[2255:2248]} - {1'b0, layer_1_0[2255:2248]};
      mid_1[0] = {1'b0,layer_2_1[2239:2232]} - {1'b0, layer_1_1[2239:2232]};
      mid_1[1] = {1'b0,layer_2_1[2247:2240]} - {1'b0, layer_1_1[2247:2240]};
      mid_1[2] = {1'b0,layer_2_1[2255:2248]} - {1'b0, layer_1_1[2255:2248]};
      mid_2[0] = {1'b0,layer_2_2[2239:2232]} - {1'b0, layer_1_2[2239:2232]};
      mid_2[1] = {1'b0,layer_2_2[2247:2240]} - {1'b0, layer_1_2[2247:2240]};
      mid_2[2] = {1'b0,layer_2_2[2255:2248]} - {1'b0, layer_1_2[2255:2248]};
      btm_0[0] = {1'b0,layer_3_0[2239:2232]} - {1'b0, layer_2_0[2239:2232]};
      btm_0[1] = {1'b0,layer_3_0[2247:2240]} - {1'b0, layer_2_0[2247:2240]};
      btm_0[2] = {1'b0,layer_3_0[2255:2248]} - {1'b0, layer_2_0[2255:2248]};
      btm_1[0] = {1'b0,layer_3_1[2239:2232]} - {1'b0, layer_2_1[2239:2232]};
      btm_1[1] = {1'b0,layer_3_1[2247:2240]} - {1'b0, layer_2_1[2247:2240]};
      btm_1[2] = {1'b0,layer_3_1[2255:2248]} - {1'b0, layer_2_1[2255:2248]};
      btm_2[0] = {1'b0,layer_3_2[2239:2232]} - {1'b0, layer_2_2[2239:2232]};
      btm_2[1] = {1'b0,layer_3_2[2247:2240]} - {1'b0, layer_2_2[2247:2240]};
      btm_2[2] = {1'b0,layer_3_2[2255:2248]} - {1'b0, layer_2_2[2255:2248]};
    end
    'd281: begin
      top_0[0] = {1'b0,layer_1_0[2247:2240]} - {1'b0, layer_0_0[2247:2240]};
      top_0[1] = {1'b0,layer_1_0[2255:2248]} - {1'b0, layer_0_0[2255:2248]};
      top_0[2] = {1'b0,layer_1_0[2263:2256]} - {1'b0, layer_0_0[2263:2256]};
      top_1[0] = {1'b0,layer_1_1[2247:2240]} - {1'b0, layer_0_1[2247:2240]};
      top_1[1] = {1'b0,layer_1_1[2255:2248]} - {1'b0, layer_0_1[2255:2248]};
      top_1[2] = {1'b0,layer_1_1[2263:2256]} - {1'b0, layer_0_1[2263:2256]};
      top_2[0] = {1'b0,layer_1_2[2247:2240]} - {1'b0, layer_0_2[2247:2240]};
      top_2[1] = {1'b0,layer_1_2[2255:2248]} - {1'b0, layer_0_2[2255:2248]};
      top_2[2] = {1'b0,layer_1_2[2263:2256]} - {1'b0, layer_0_2[2263:2256]};
      mid_0[0] = {1'b0,layer_2_0[2247:2240]} - {1'b0, layer_1_0[2247:2240]};
      mid_0[1] = {1'b0,layer_2_0[2255:2248]} - {1'b0, layer_1_0[2255:2248]};
      mid_0[2] = {1'b0,layer_2_0[2263:2256]} - {1'b0, layer_1_0[2263:2256]};
      mid_1[0] = {1'b0,layer_2_1[2247:2240]} - {1'b0, layer_1_1[2247:2240]};
      mid_1[1] = {1'b0,layer_2_1[2255:2248]} - {1'b0, layer_1_1[2255:2248]};
      mid_1[2] = {1'b0,layer_2_1[2263:2256]} - {1'b0, layer_1_1[2263:2256]};
      mid_2[0] = {1'b0,layer_2_2[2247:2240]} - {1'b0, layer_1_2[2247:2240]};
      mid_2[1] = {1'b0,layer_2_2[2255:2248]} - {1'b0, layer_1_2[2255:2248]};
      mid_2[2] = {1'b0,layer_2_2[2263:2256]} - {1'b0, layer_1_2[2263:2256]};
      btm_0[0] = {1'b0,layer_3_0[2247:2240]} - {1'b0, layer_2_0[2247:2240]};
      btm_0[1] = {1'b0,layer_3_0[2255:2248]} - {1'b0, layer_2_0[2255:2248]};
      btm_0[2] = {1'b0,layer_3_0[2263:2256]} - {1'b0, layer_2_0[2263:2256]};
      btm_1[0] = {1'b0,layer_3_1[2247:2240]} - {1'b0, layer_2_1[2247:2240]};
      btm_1[1] = {1'b0,layer_3_1[2255:2248]} - {1'b0, layer_2_1[2255:2248]};
      btm_1[2] = {1'b0,layer_3_1[2263:2256]} - {1'b0, layer_2_1[2263:2256]};
      btm_2[0] = {1'b0,layer_3_2[2247:2240]} - {1'b0, layer_2_2[2247:2240]};
      btm_2[1] = {1'b0,layer_3_2[2255:2248]} - {1'b0, layer_2_2[2255:2248]};
      btm_2[2] = {1'b0,layer_3_2[2263:2256]} - {1'b0, layer_2_2[2263:2256]};
    end
    'd282: begin
      top_0[0] = {1'b0,layer_1_0[2255:2248]} - {1'b0, layer_0_0[2255:2248]};
      top_0[1] = {1'b0,layer_1_0[2263:2256]} - {1'b0, layer_0_0[2263:2256]};
      top_0[2] = {1'b0,layer_1_0[2271:2264]} - {1'b0, layer_0_0[2271:2264]};
      top_1[0] = {1'b0,layer_1_1[2255:2248]} - {1'b0, layer_0_1[2255:2248]};
      top_1[1] = {1'b0,layer_1_1[2263:2256]} - {1'b0, layer_0_1[2263:2256]};
      top_1[2] = {1'b0,layer_1_1[2271:2264]} - {1'b0, layer_0_1[2271:2264]};
      top_2[0] = {1'b0,layer_1_2[2255:2248]} - {1'b0, layer_0_2[2255:2248]};
      top_2[1] = {1'b0,layer_1_2[2263:2256]} - {1'b0, layer_0_2[2263:2256]};
      top_2[2] = {1'b0,layer_1_2[2271:2264]} - {1'b0, layer_0_2[2271:2264]};
      mid_0[0] = {1'b0,layer_2_0[2255:2248]} - {1'b0, layer_1_0[2255:2248]};
      mid_0[1] = {1'b0,layer_2_0[2263:2256]} - {1'b0, layer_1_0[2263:2256]};
      mid_0[2] = {1'b0,layer_2_0[2271:2264]} - {1'b0, layer_1_0[2271:2264]};
      mid_1[0] = {1'b0,layer_2_1[2255:2248]} - {1'b0, layer_1_1[2255:2248]};
      mid_1[1] = {1'b0,layer_2_1[2263:2256]} - {1'b0, layer_1_1[2263:2256]};
      mid_1[2] = {1'b0,layer_2_1[2271:2264]} - {1'b0, layer_1_1[2271:2264]};
      mid_2[0] = {1'b0,layer_2_2[2255:2248]} - {1'b0, layer_1_2[2255:2248]};
      mid_2[1] = {1'b0,layer_2_2[2263:2256]} - {1'b0, layer_1_2[2263:2256]};
      mid_2[2] = {1'b0,layer_2_2[2271:2264]} - {1'b0, layer_1_2[2271:2264]};
      btm_0[0] = {1'b0,layer_3_0[2255:2248]} - {1'b0, layer_2_0[2255:2248]};
      btm_0[1] = {1'b0,layer_3_0[2263:2256]} - {1'b0, layer_2_0[2263:2256]};
      btm_0[2] = {1'b0,layer_3_0[2271:2264]} - {1'b0, layer_2_0[2271:2264]};
      btm_1[0] = {1'b0,layer_3_1[2255:2248]} - {1'b0, layer_2_1[2255:2248]};
      btm_1[1] = {1'b0,layer_3_1[2263:2256]} - {1'b0, layer_2_1[2263:2256]};
      btm_1[2] = {1'b0,layer_3_1[2271:2264]} - {1'b0, layer_2_1[2271:2264]};
      btm_2[0] = {1'b0,layer_3_2[2255:2248]} - {1'b0, layer_2_2[2255:2248]};
      btm_2[1] = {1'b0,layer_3_2[2263:2256]} - {1'b0, layer_2_2[2263:2256]};
      btm_2[2] = {1'b0,layer_3_2[2271:2264]} - {1'b0, layer_2_2[2271:2264]};
    end
    'd283: begin
      top_0[0] = {1'b0,layer_1_0[2263:2256]} - {1'b0, layer_0_0[2263:2256]};
      top_0[1] = {1'b0,layer_1_0[2271:2264]} - {1'b0, layer_0_0[2271:2264]};
      top_0[2] = {1'b0,layer_1_0[2279:2272]} - {1'b0, layer_0_0[2279:2272]};
      top_1[0] = {1'b0,layer_1_1[2263:2256]} - {1'b0, layer_0_1[2263:2256]};
      top_1[1] = {1'b0,layer_1_1[2271:2264]} - {1'b0, layer_0_1[2271:2264]};
      top_1[2] = {1'b0,layer_1_1[2279:2272]} - {1'b0, layer_0_1[2279:2272]};
      top_2[0] = {1'b0,layer_1_2[2263:2256]} - {1'b0, layer_0_2[2263:2256]};
      top_2[1] = {1'b0,layer_1_2[2271:2264]} - {1'b0, layer_0_2[2271:2264]};
      top_2[2] = {1'b0,layer_1_2[2279:2272]} - {1'b0, layer_0_2[2279:2272]};
      mid_0[0] = {1'b0,layer_2_0[2263:2256]} - {1'b0, layer_1_0[2263:2256]};
      mid_0[1] = {1'b0,layer_2_0[2271:2264]} - {1'b0, layer_1_0[2271:2264]};
      mid_0[2] = {1'b0,layer_2_0[2279:2272]} - {1'b0, layer_1_0[2279:2272]};
      mid_1[0] = {1'b0,layer_2_1[2263:2256]} - {1'b0, layer_1_1[2263:2256]};
      mid_1[1] = {1'b0,layer_2_1[2271:2264]} - {1'b0, layer_1_1[2271:2264]};
      mid_1[2] = {1'b0,layer_2_1[2279:2272]} - {1'b0, layer_1_1[2279:2272]};
      mid_2[0] = {1'b0,layer_2_2[2263:2256]} - {1'b0, layer_1_2[2263:2256]};
      mid_2[1] = {1'b0,layer_2_2[2271:2264]} - {1'b0, layer_1_2[2271:2264]};
      mid_2[2] = {1'b0,layer_2_2[2279:2272]} - {1'b0, layer_1_2[2279:2272]};
      btm_0[0] = {1'b0,layer_3_0[2263:2256]} - {1'b0, layer_2_0[2263:2256]};
      btm_0[1] = {1'b0,layer_3_0[2271:2264]} - {1'b0, layer_2_0[2271:2264]};
      btm_0[2] = {1'b0,layer_3_0[2279:2272]} - {1'b0, layer_2_0[2279:2272]};
      btm_1[0] = {1'b0,layer_3_1[2263:2256]} - {1'b0, layer_2_1[2263:2256]};
      btm_1[1] = {1'b0,layer_3_1[2271:2264]} - {1'b0, layer_2_1[2271:2264]};
      btm_1[2] = {1'b0,layer_3_1[2279:2272]} - {1'b0, layer_2_1[2279:2272]};
      btm_2[0] = {1'b0,layer_3_2[2263:2256]} - {1'b0, layer_2_2[2263:2256]};
      btm_2[1] = {1'b0,layer_3_2[2271:2264]} - {1'b0, layer_2_2[2271:2264]};
      btm_2[2] = {1'b0,layer_3_2[2279:2272]} - {1'b0, layer_2_2[2279:2272]};
    end
    'd284: begin
      top_0[0] = {1'b0,layer_1_0[2271:2264]} - {1'b0, layer_0_0[2271:2264]};
      top_0[1] = {1'b0,layer_1_0[2279:2272]} - {1'b0, layer_0_0[2279:2272]};
      top_0[2] = {1'b0,layer_1_0[2287:2280]} - {1'b0, layer_0_0[2287:2280]};
      top_1[0] = {1'b0,layer_1_1[2271:2264]} - {1'b0, layer_0_1[2271:2264]};
      top_1[1] = {1'b0,layer_1_1[2279:2272]} - {1'b0, layer_0_1[2279:2272]};
      top_1[2] = {1'b0,layer_1_1[2287:2280]} - {1'b0, layer_0_1[2287:2280]};
      top_2[0] = {1'b0,layer_1_2[2271:2264]} - {1'b0, layer_0_2[2271:2264]};
      top_2[1] = {1'b0,layer_1_2[2279:2272]} - {1'b0, layer_0_2[2279:2272]};
      top_2[2] = {1'b0,layer_1_2[2287:2280]} - {1'b0, layer_0_2[2287:2280]};
      mid_0[0] = {1'b0,layer_2_0[2271:2264]} - {1'b0, layer_1_0[2271:2264]};
      mid_0[1] = {1'b0,layer_2_0[2279:2272]} - {1'b0, layer_1_0[2279:2272]};
      mid_0[2] = {1'b0,layer_2_0[2287:2280]} - {1'b0, layer_1_0[2287:2280]};
      mid_1[0] = {1'b0,layer_2_1[2271:2264]} - {1'b0, layer_1_1[2271:2264]};
      mid_1[1] = {1'b0,layer_2_1[2279:2272]} - {1'b0, layer_1_1[2279:2272]};
      mid_1[2] = {1'b0,layer_2_1[2287:2280]} - {1'b0, layer_1_1[2287:2280]};
      mid_2[0] = {1'b0,layer_2_2[2271:2264]} - {1'b0, layer_1_2[2271:2264]};
      mid_2[1] = {1'b0,layer_2_2[2279:2272]} - {1'b0, layer_1_2[2279:2272]};
      mid_2[2] = {1'b0,layer_2_2[2287:2280]} - {1'b0, layer_1_2[2287:2280]};
      btm_0[0] = {1'b0,layer_3_0[2271:2264]} - {1'b0, layer_2_0[2271:2264]};
      btm_0[1] = {1'b0,layer_3_0[2279:2272]} - {1'b0, layer_2_0[2279:2272]};
      btm_0[2] = {1'b0,layer_3_0[2287:2280]} - {1'b0, layer_2_0[2287:2280]};
      btm_1[0] = {1'b0,layer_3_1[2271:2264]} - {1'b0, layer_2_1[2271:2264]};
      btm_1[1] = {1'b0,layer_3_1[2279:2272]} - {1'b0, layer_2_1[2279:2272]};
      btm_1[2] = {1'b0,layer_3_1[2287:2280]} - {1'b0, layer_2_1[2287:2280]};
      btm_2[0] = {1'b0,layer_3_2[2271:2264]} - {1'b0, layer_2_2[2271:2264]};
      btm_2[1] = {1'b0,layer_3_2[2279:2272]} - {1'b0, layer_2_2[2279:2272]};
      btm_2[2] = {1'b0,layer_3_2[2287:2280]} - {1'b0, layer_2_2[2287:2280]};
    end
    'd285: begin
      top_0[0] = {1'b0,layer_1_0[2279:2272]} - {1'b0, layer_0_0[2279:2272]};
      top_0[1] = {1'b0,layer_1_0[2287:2280]} - {1'b0, layer_0_0[2287:2280]};
      top_0[2] = {1'b0,layer_1_0[2295:2288]} - {1'b0, layer_0_0[2295:2288]};
      top_1[0] = {1'b0,layer_1_1[2279:2272]} - {1'b0, layer_0_1[2279:2272]};
      top_1[1] = {1'b0,layer_1_1[2287:2280]} - {1'b0, layer_0_1[2287:2280]};
      top_1[2] = {1'b0,layer_1_1[2295:2288]} - {1'b0, layer_0_1[2295:2288]};
      top_2[0] = {1'b0,layer_1_2[2279:2272]} - {1'b0, layer_0_2[2279:2272]};
      top_2[1] = {1'b0,layer_1_2[2287:2280]} - {1'b0, layer_0_2[2287:2280]};
      top_2[2] = {1'b0,layer_1_2[2295:2288]} - {1'b0, layer_0_2[2295:2288]};
      mid_0[0] = {1'b0,layer_2_0[2279:2272]} - {1'b0, layer_1_0[2279:2272]};
      mid_0[1] = {1'b0,layer_2_0[2287:2280]} - {1'b0, layer_1_0[2287:2280]};
      mid_0[2] = {1'b0,layer_2_0[2295:2288]} - {1'b0, layer_1_0[2295:2288]};
      mid_1[0] = {1'b0,layer_2_1[2279:2272]} - {1'b0, layer_1_1[2279:2272]};
      mid_1[1] = {1'b0,layer_2_1[2287:2280]} - {1'b0, layer_1_1[2287:2280]};
      mid_1[2] = {1'b0,layer_2_1[2295:2288]} - {1'b0, layer_1_1[2295:2288]};
      mid_2[0] = {1'b0,layer_2_2[2279:2272]} - {1'b0, layer_1_2[2279:2272]};
      mid_2[1] = {1'b0,layer_2_2[2287:2280]} - {1'b0, layer_1_2[2287:2280]};
      mid_2[2] = {1'b0,layer_2_2[2295:2288]} - {1'b0, layer_1_2[2295:2288]};
      btm_0[0] = {1'b0,layer_3_0[2279:2272]} - {1'b0, layer_2_0[2279:2272]};
      btm_0[1] = {1'b0,layer_3_0[2287:2280]} - {1'b0, layer_2_0[2287:2280]};
      btm_0[2] = {1'b0,layer_3_0[2295:2288]} - {1'b0, layer_2_0[2295:2288]};
      btm_1[0] = {1'b0,layer_3_1[2279:2272]} - {1'b0, layer_2_1[2279:2272]};
      btm_1[1] = {1'b0,layer_3_1[2287:2280]} - {1'b0, layer_2_1[2287:2280]};
      btm_1[2] = {1'b0,layer_3_1[2295:2288]} - {1'b0, layer_2_1[2295:2288]};
      btm_2[0] = {1'b0,layer_3_2[2279:2272]} - {1'b0, layer_2_2[2279:2272]};
      btm_2[1] = {1'b0,layer_3_2[2287:2280]} - {1'b0, layer_2_2[2287:2280]};
      btm_2[2] = {1'b0,layer_3_2[2295:2288]} - {1'b0, layer_2_2[2295:2288]};
    end
    'd286: begin
      top_0[0] = {1'b0,layer_1_0[2287:2280]} - {1'b0, layer_0_0[2287:2280]};
      top_0[1] = {1'b0,layer_1_0[2295:2288]} - {1'b0, layer_0_0[2295:2288]};
      top_0[2] = {1'b0,layer_1_0[2303:2296]} - {1'b0, layer_0_0[2303:2296]};
      top_1[0] = {1'b0,layer_1_1[2287:2280]} - {1'b0, layer_0_1[2287:2280]};
      top_1[1] = {1'b0,layer_1_1[2295:2288]} - {1'b0, layer_0_1[2295:2288]};
      top_1[2] = {1'b0,layer_1_1[2303:2296]} - {1'b0, layer_0_1[2303:2296]};
      top_2[0] = {1'b0,layer_1_2[2287:2280]} - {1'b0, layer_0_2[2287:2280]};
      top_2[1] = {1'b0,layer_1_2[2295:2288]} - {1'b0, layer_0_2[2295:2288]};
      top_2[2] = {1'b0,layer_1_2[2303:2296]} - {1'b0, layer_0_2[2303:2296]};
      mid_0[0] = {1'b0,layer_2_0[2287:2280]} - {1'b0, layer_1_0[2287:2280]};
      mid_0[1] = {1'b0,layer_2_0[2295:2288]} - {1'b0, layer_1_0[2295:2288]};
      mid_0[2] = {1'b0,layer_2_0[2303:2296]} - {1'b0, layer_1_0[2303:2296]};
      mid_1[0] = {1'b0,layer_2_1[2287:2280]} - {1'b0, layer_1_1[2287:2280]};
      mid_1[1] = {1'b0,layer_2_1[2295:2288]} - {1'b0, layer_1_1[2295:2288]};
      mid_1[2] = {1'b0,layer_2_1[2303:2296]} - {1'b0, layer_1_1[2303:2296]};
      mid_2[0] = {1'b0,layer_2_2[2287:2280]} - {1'b0, layer_1_2[2287:2280]};
      mid_2[1] = {1'b0,layer_2_2[2295:2288]} - {1'b0, layer_1_2[2295:2288]};
      mid_2[2] = {1'b0,layer_2_2[2303:2296]} - {1'b0, layer_1_2[2303:2296]};
      btm_0[0] = {1'b0,layer_3_0[2287:2280]} - {1'b0, layer_2_0[2287:2280]};
      btm_0[1] = {1'b0,layer_3_0[2295:2288]} - {1'b0, layer_2_0[2295:2288]};
      btm_0[2] = {1'b0,layer_3_0[2303:2296]} - {1'b0, layer_2_0[2303:2296]};
      btm_1[0] = {1'b0,layer_3_1[2287:2280]} - {1'b0, layer_2_1[2287:2280]};
      btm_1[1] = {1'b0,layer_3_1[2295:2288]} - {1'b0, layer_2_1[2295:2288]};
      btm_1[2] = {1'b0,layer_3_1[2303:2296]} - {1'b0, layer_2_1[2303:2296]};
      btm_2[0] = {1'b0,layer_3_2[2287:2280]} - {1'b0, layer_2_2[2287:2280]};
      btm_2[1] = {1'b0,layer_3_2[2295:2288]} - {1'b0, layer_2_2[2295:2288]};
      btm_2[2] = {1'b0,layer_3_2[2303:2296]} - {1'b0, layer_2_2[2303:2296]};
    end
    'd287: begin
      top_0[0] = {1'b0,layer_1_0[2295:2288]} - {1'b0, layer_0_0[2295:2288]};
      top_0[1] = {1'b0,layer_1_0[2303:2296]} - {1'b0, layer_0_0[2303:2296]};
      top_0[2] = {1'b0,layer_1_0[2311:2304]} - {1'b0, layer_0_0[2311:2304]};
      top_1[0] = {1'b0,layer_1_1[2295:2288]} - {1'b0, layer_0_1[2295:2288]};
      top_1[1] = {1'b0,layer_1_1[2303:2296]} - {1'b0, layer_0_1[2303:2296]};
      top_1[2] = {1'b0,layer_1_1[2311:2304]} - {1'b0, layer_0_1[2311:2304]};
      top_2[0] = {1'b0,layer_1_2[2295:2288]} - {1'b0, layer_0_2[2295:2288]};
      top_2[1] = {1'b0,layer_1_2[2303:2296]} - {1'b0, layer_0_2[2303:2296]};
      top_2[2] = {1'b0,layer_1_2[2311:2304]} - {1'b0, layer_0_2[2311:2304]};
      mid_0[0] = {1'b0,layer_2_0[2295:2288]} - {1'b0, layer_1_0[2295:2288]};
      mid_0[1] = {1'b0,layer_2_0[2303:2296]} - {1'b0, layer_1_0[2303:2296]};
      mid_0[2] = {1'b0,layer_2_0[2311:2304]} - {1'b0, layer_1_0[2311:2304]};
      mid_1[0] = {1'b0,layer_2_1[2295:2288]} - {1'b0, layer_1_1[2295:2288]};
      mid_1[1] = {1'b0,layer_2_1[2303:2296]} - {1'b0, layer_1_1[2303:2296]};
      mid_1[2] = {1'b0,layer_2_1[2311:2304]} - {1'b0, layer_1_1[2311:2304]};
      mid_2[0] = {1'b0,layer_2_2[2295:2288]} - {1'b0, layer_1_2[2295:2288]};
      mid_2[1] = {1'b0,layer_2_2[2303:2296]} - {1'b0, layer_1_2[2303:2296]};
      mid_2[2] = {1'b0,layer_2_2[2311:2304]} - {1'b0, layer_1_2[2311:2304]};
      btm_0[0] = {1'b0,layer_3_0[2295:2288]} - {1'b0, layer_2_0[2295:2288]};
      btm_0[1] = {1'b0,layer_3_0[2303:2296]} - {1'b0, layer_2_0[2303:2296]};
      btm_0[2] = {1'b0,layer_3_0[2311:2304]} - {1'b0, layer_2_0[2311:2304]};
      btm_1[0] = {1'b0,layer_3_1[2295:2288]} - {1'b0, layer_2_1[2295:2288]};
      btm_1[1] = {1'b0,layer_3_1[2303:2296]} - {1'b0, layer_2_1[2303:2296]};
      btm_1[2] = {1'b0,layer_3_1[2311:2304]} - {1'b0, layer_2_1[2311:2304]};
      btm_2[0] = {1'b0,layer_3_2[2295:2288]} - {1'b0, layer_2_2[2295:2288]};
      btm_2[1] = {1'b0,layer_3_2[2303:2296]} - {1'b0, layer_2_2[2303:2296]};
      btm_2[2] = {1'b0,layer_3_2[2311:2304]} - {1'b0, layer_2_2[2311:2304]};
    end
    'd288: begin
      top_0[0] = {1'b0,layer_1_0[2303:2296]} - {1'b0, layer_0_0[2303:2296]};
      top_0[1] = {1'b0,layer_1_0[2311:2304]} - {1'b0, layer_0_0[2311:2304]};
      top_0[2] = {1'b0,layer_1_0[2319:2312]} - {1'b0, layer_0_0[2319:2312]};
      top_1[0] = {1'b0,layer_1_1[2303:2296]} - {1'b0, layer_0_1[2303:2296]};
      top_1[1] = {1'b0,layer_1_1[2311:2304]} - {1'b0, layer_0_1[2311:2304]};
      top_1[2] = {1'b0,layer_1_1[2319:2312]} - {1'b0, layer_0_1[2319:2312]};
      top_2[0] = {1'b0,layer_1_2[2303:2296]} - {1'b0, layer_0_2[2303:2296]};
      top_2[1] = {1'b0,layer_1_2[2311:2304]} - {1'b0, layer_0_2[2311:2304]};
      top_2[2] = {1'b0,layer_1_2[2319:2312]} - {1'b0, layer_0_2[2319:2312]};
      mid_0[0] = {1'b0,layer_2_0[2303:2296]} - {1'b0, layer_1_0[2303:2296]};
      mid_0[1] = {1'b0,layer_2_0[2311:2304]} - {1'b0, layer_1_0[2311:2304]};
      mid_0[2] = {1'b0,layer_2_0[2319:2312]} - {1'b0, layer_1_0[2319:2312]};
      mid_1[0] = {1'b0,layer_2_1[2303:2296]} - {1'b0, layer_1_1[2303:2296]};
      mid_1[1] = {1'b0,layer_2_1[2311:2304]} - {1'b0, layer_1_1[2311:2304]};
      mid_1[2] = {1'b0,layer_2_1[2319:2312]} - {1'b0, layer_1_1[2319:2312]};
      mid_2[0] = {1'b0,layer_2_2[2303:2296]} - {1'b0, layer_1_2[2303:2296]};
      mid_2[1] = {1'b0,layer_2_2[2311:2304]} - {1'b0, layer_1_2[2311:2304]};
      mid_2[2] = {1'b0,layer_2_2[2319:2312]} - {1'b0, layer_1_2[2319:2312]};
      btm_0[0] = {1'b0,layer_3_0[2303:2296]} - {1'b0, layer_2_0[2303:2296]};
      btm_0[1] = {1'b0,layer_3_0[2311:2304]} - {1'b0, layer_2_0[2311:2304]};
      btm_0[2] = {1'b0,layer_3_0[2319:2312]} - {1'b0, layer_2_0[2319:2312]};
      btm_1[0] = {1'b0,layer_3_1[2303:2296]} - {1'b0, layer_2_1[2303:2296]};
      btm_1[1] = {1'b0,layer_3_1[2311:2304]} - {1'b0, layer_2_1[2311:2304]};
      btm_1[2] = {1'b0,layer_3_1[2319:2312]} - {1'b0, layer_2_1[2319:2312]};
      btm_2[0] = {1'b0,layer_3_2[2303:2296]} - {1'b0, layer_2_2[2303:2296]};
      btm_2[1] = {1'b0,layer_3_2[2311:2304]} - {1'b0, layer_2_2[2311:2304]};
      btm_2[2] = {1'b0,layer_3_2[2319:2312]} - {1'b0, layer_2_2[2319:2312]};
    end
    'd289: begin
      top_0[0] = {1'b0,layer_1_0[2311:2304]} - {1'b0, layer_0_0[2311:2304]};
      top_0[1] = {1'b0,layer_1_0[2319:2312]} - {1'b0, layer_0_0[2319:2312]};
      top_0[2] = {1'b0,layer_1_0[2327:2320]} - {1'b0, layer_0_0[2327:2320]};
      top_1[0] = {1'b0,layer_1_1[2311:2304]} - {1'b0, layer_0_1[2311:2304]};
      top_1[1] = {1'b0,layer_1_1[2319:2312]} - {1'b0, layer_0_1[2319:2312]};
      top_1[2] = {1'b0,layer_1_1[2327:2320]} - {1'b0, layer_0_1[2327:2320]};
      top_2[0] = {1'b0,layer_1_2[2311:2304]} - {1'b0, layer_0_2[2311:2304]};
      top_2[1] = {1'b0,layer_1_2[2319:2312]} - {1'b0, layer_0_2[2319:2312]};
      top_2[2] = {1'b0,layer_1_2[2327:2320]} - {1'b0, layer_0_2[2327:2320]};
      mid_0[0] = {1'b0,layer_2_0[2311:2304]} - {1'b0, layer_1_0[2311:2304]};
      mid_0[1] = {1'b0,layer_2_0[2319:2312]} - {1'b0, layer_1_0[2319:2312]};
      mid_0[2] = {1'b0,layer_2_0[2327:2320]} - {1'b0, layer_1_0[2327:2320]};
      mid_1[0] = {1'b0,layer_2_1[2311:2304]} - {1'b0, layer_1_1[2311:2304]};
      mid_1[1] = {1'b0,layer_2_1[2319:2312]} - {1'b0, layer_1_1[2319:2312]};
      mid_1[2] = {1'b0,layer_2_1[2327:2320]} - {1'b0, layer_1_1[2327:2320]};
      mid_2[0] = {1'b0,layer_2_2[2311:2304]} - {1'b0, layer_1_2[2311:2304]};
      mid_2[1] = {1'b0,layer_2_2[2319:2312]} - {1'b0, layer_1_2[2319:2312]};
      mid_2[2] = {1'b0,layer_2_2[2327:2320]} - {1'b0, layer_1_2[2327:2320]};
      btm_0[0] = {1'b0,layer_3_0[2311:2304]} - {1'b0, layer_2_0[2311:2304]};
      btm_0[1] = {1'b0,layer_3_0[2319:2312]} - {1'b0, layer_2_0[2319:2312]};
      btm_0[2] = {1'b0,layer_3_0[2327:2320]} - {1'b0, layer_2_0[2327:2320]};
      btm_1[0] = {1'b0,layer_3_1[2311:2304]} - {1'b0, layer_2_1[2311:2304]};
      btm_1[1] = {1'b0,layer_3_1[2319:2312]} - {1'b0, layer_2_1[2319:2312]};
      btm_1[2] = {1'b0,layer_3_1[2327:2320]} - {1'b0, layer_2_1[2327:2320]};
      btm_2[0] = {1'b0,layer_3_2[2311:2304]} - {1'b0, layer_2_2[2311:2304]};
      btm_2[1] = {1'b0,layer_3_2[2319:2312]} - {1'b0, layer_2_2[2319:2312]};
      btm_2[2] = {1'b0,layer_3_2[2327:2320]} - {1'b0, layer_2_2[2327:2320]};
    end
    'd290: begin
      top_0[0] = {1'b0,layer_1_0[2319:2312]} - {1'b0, layer_0_0[2319:2312]};
      top_0[1] = {1'b0,layer_1_0[2327:2320]} - {1'b0, layer_0_0[2327:2320]};
      top_0[2] = {1'b0,layer_1_0[2335:2328]} - {1'b0, layer_0_0[2335:2328]};
      top_1[0] = {1'b0,layer_1_1[2319:2312]} - {1'b0, layer_0_1[2319:2312]};
      top_1[1] = {1'b0,layer_1_1[2327:2320]} - {1'b0, layer_0_1[2327:2320]};
      top_1[2] = {1'b0,layer_1_1[2335:2328]} - {1'b0, layer_0_1[2335:2328]};
      top_2[0] = {1'b0,layer_1_2[2319:2312]} - {1'b0, layer_0_2[2319:2312]};
      top_2[1] = {1'b0,layer_1_2[2327:2320]} - {1'b0, layer_0_2[2327:2320]};
      top_2[2] = {1'b0,layer_1_2[2335:2328]} - {1'b0, layer_0_2[2335:2328]};
      mid_0[0] = {1'b0,layer_2_0[2319:2312]} - {1'b0, layer_1_0[2319:2312]};
      mid_0[1] = {1'b0,layer_2_0[2327:2320]} - {1'b0, layer_1_0[2327:2320]};
      mid_0[2] = {1'b0,layer_2_0[2335:2328]} - {1'b0, layer_1_0[2335:2328]};
      mid_1[0] = {1'b0,layer_2_1[2319:2312]} - {1'b0, layer_1_1[2319:2312]};
      mid_1[1] = {1'b0,layer_2_1[2327:2320]} - {1'b0, layer_1_1[2327:2320]};
      mid_1[2] = {1'b0,layer_2_1[2335:2328]} - {1'b0, layer_1_1[2335:2328]};
      mid_2[0] = {1'b0,layer_2_2[2319:2312]} - {1'b0, layer_1_2[2319:2312]};
      mid_2[1] = {1'b0,layer_2_2[2327:2320]} - {1'b0, layer_1_2[2327:2320]};
      mid_2[2] = {1'b0,layer_2_2[2335:2328]} - {1'b0, layer_1_2[2335:2328]};
      btm_0[0] = {1'b0,layer_3_0[2319:2312]} - {1'b0, layer_2_0[2319:2312]};
      btm_0[1] = {1'b0,layer_3_0[2327:2320]} - {1'b0, layer_2_0[2327:2320]};
      btm_0[2] = {1'b0,layer_3_0[2335:2328]} - {1'b0, layer_2_0[2335:2328]};
      btm_1[0] = {1'b0,layer_3_1[2319:2312]} - {1'b0, layer_2_1[2319:2312]};
      btm_1[1] = {1'b0,layer_3_1[2327:2320]} - {1'b0, layer_2_1[2327:2320]};
      btm_1[2] = {1'b0,layer_3_1[2335:2328]} - {1'b0, layer_2_1[2335:2328]};
      btm_2[0] = {1'b0,layer_3_2[2319:2312]} - {1'b0, layer_2_2[2319:2312]};
      btm_2[1] = {1'b0,layer_3_2[2327:2320]} - {1'b0, layer_2_2[2327:2320]};
      btm_2[2] = {1'b0,layer_3_2[2335:2328]} - {1'b0, layer_2_2[2335:2328]};
    end
    'd291: begin
      top_0[0] = {1'b0,layer_1_0[2327:2320]} - {1'b0, layer_0_0[2327:2320]};
      top_0[1] = {1'b0,layer_1_0[2335:2328]} - {1'b0, layer_0_0[2335:2328]};
      top_0[2] = {1'b0,layer_1_0[2343:2336]} - {1'b0, layer_0_0[2343:2336]};
      top_1[0] = {1'b0,layer_1_1[2327:2320]} - {1'b0, layer_0_1[2327:2320]};
      top_1[1] = {1'b0,layer_1_1[2335:2328]} - {1'b0, layer_0_1[2335:2328]};
      top_1[2] = {1'b0,layer_1_1[2343:2336]} - {1'b0, layer_0_1[2343:2336]};
      top_2[0] = {1'b0,layer_1_2[2327:2320]} - {1'b0, layer_0_2[2327:2320]};
      top_2[1] = {1'b0,layer_1_2[2335:2328]} - {1'b0, layer_0_2[2335:2328]};
      top_2[2] = {1'b0,layer_1_2[2343:2336]} - {1'b0, layer_0_2[2343:2336]};
      mid_0[0] = {1'b0,layer_2_0[2327:2320]} - {1'b0, layer_1_0[2327:2320]};
      mid_0[1] = {1'b0,layer_2_0[2335:2328]} - {1'b0, layer_1_0[2335:2328]};
      mid_0[2] = {1'b0,layer_2_0[2343:2336]} - {1'b0, layer_1_0[2343:2336]};
      mid_1[0] = {1'b0,layer_2_1[2327:2320]} - {1'b0, layer_1_1[2327:2320]};
      mid_1[1] = {1'b0,layer_2_1[2335:2328]} - {1'b0, layer_1_1[2335:2328]};
      mid_1[2] = {1'b0,layer_2_1[2343:2336]} - {1'b0, layer_1_1[2343:2336]};
      mid_2[0] = {1'b0,layer_2_2[2327:2320]} - {1'b0, layer_1_2[2327:2320]};
      mid_2[1] = {1'b0,layer_2_2[2335:2328]} - {1'b0, layer_1_2[2335:2328]};
      mid_2[2] = {1'b0,layer_2_2[2343:2336]} - {1'b0, layer_1_2[2343:2336]};
      btm_0[0] = {1'b0,layer_3_0[2327:2320]} - {1'b0, layer_2_0[2327:2320]};
      btm_0[1] = {1'b0,layer_3_0[2335:2328]} - {1'b0, layer_2_0[2335:2328]};
      btm_0[2] = {1'b0,layer_3_0[2343:2336]} - {1'b0, layer_2_0[2343:2336]};
      btm_1[0] = {1'b0,layer_3_1[2327:2320]} - {1'b0, layer_2_1[2327:2320]};
      btm_1[1] = {1'b0,layer_3_1[2335:2328]} - {1'b0, layer_2_1[2335:2328]};
      btm_1[2] = {1'b0,layer_3_1[2343:2336]} - {1'b0, layer_2_1[2343:2336]};
      btm_2[0] = {1'b0,layer_3_2[2327:2320]} - {1'b0, layer_2_2[2327:2320]};
      btm_2[1] = {1'b0,layer_3_2[2335:2328]} - {1'b0, layer_2_2[2335:2328]};
      btm_2[2] = {1'b0,layer_3_2[2343:2336]} - {1'b0, layer_2_2[2343:2336]};
    end
    'd292: begin
      top_0[0] = {1'b0,layer_1_0[2335:2328]} - {1'b0, layer_0_0[2335:2328]};
      top_0[1] = {1'b0,layer_1_0[2343:2336]} - {1'b0, layer_0_0[2343:2336]};
      top_0[2] = {1'b0,layer_1_0[2351:2344]} - {1'b0, layer_0_0[2351:2344]};
      top_1[0] = {1'b0,layer_1_1[2335:2328]} - {1'b0, layer_0_1[2335:2328]};
      top_1[1] = {1'b0,layer_1_1[2343:2336]} - {1'b0, layer_0_1[2343:2336]};
      top_1[2] = {1'b0,layer_1_1[2351:2344]} - {1'b0, layer_0_1[2351:2344]};
      top_2[0] = {1'b0,layer_1_2[2335:2328]} - {1'b0, layer_0_2[2335:2328]};
      top_2[1] = {1'b0,layer_1_2[2343:2336]} - {1'b0, layer_0_2[2343:2336]};
      top_2[2] = {1'b0,layer_1_2[2351:2344]} - {1'b0, layer_0_2[2351:2344]};
      mid_0[0] = {1'b0,layer_2_0[2335:2328]} - {1'b0, layer_1_0[2335:2328]};
      mid_0[1] = {1'b0,layer_2_0[2343:2336]} - {1'b0, layer_1_0[2343:2336]};
      mid_0[2] = {1'b0,layer_2_0[2351:2344]} - {1'b0, layer_1_0[2351:2344]};
      mid_1[0] = {1'b0,layer_2_1[2335:2328]} - {1'b0, layer_1_1[2335:2328]};
      mid_1[1] = {1'b0,layer_2_1[2343:2336]} - {1'b0, layer_1_1[2343:2336]};
      mid_1[2] = {1'b0,layer_2_1[2351:2344]} - {1'b0, layer_1_1[2351:2344]};
      mid_2[0] = {1'b0,layer_2_2[2335:2328]} - {1'b0, layer_1_2[2335:2328]};
      mid_2[1] = {1'b0,layer_2_2[2343:2336]} - {1'b0, layer_1_2[2343:2336]};
      mid_2[2] = {1'b0,layer_2_2[2351:2344]} - {1'b0, layer_1_2[2351:2344]};
      btm_0[0] = {1'b0,layer_3_0[2335:2328]} - {1'b0, layer_2_0[2335:2328]};
      btm_0[1] = {1'b0,layer_3_0[2343:2336]} - {1'b0, layer_2_0[2343:2336]};
      btm_0[2] = {1'b0,layer_3_0[2351:2344]} - {1'b0, layer_2_0[2351:2344]};
      btm_1[0] = {1'b0,layer_3_1[2335:2328]} - {1'b0, layer_2_1[2335:2328]};
      btm_1[1] = {1'b0,layer_3_1[2343:2336]} - {1'b0, layer_2_1[2343:2336]};
      btm_1[2] = {1'b0,layer_3_1[2351:2344]} - {1'b0, layer_2_1[2351:2344]};
      btm_2[0] = {1'b0,layer_3_2[2335:2328]} - {1'b0, layer_2_2[2335:2328]};
      btm_2[1] = {1'b0,layer_3_2[2343:2336]} - {1'b0, layer_2_2[2343:2336]};
      btm_2[2] = {1'b0,layer_3_2[2351:2344]} - {1'b0, layer_2_2[2351:2344]};
    end
    'd293: begin
      top_0[0] = {1'b0,layer_1_0[2343:2336]} - {1'b0, layer_0_0[2343:2336]};
      top_0[1] = {1'b0,layer_1_0[2351:2344]} - {1'b0, layer_0_0[2351:2344]};
      top_0[2] = {1'b0,layer_1_0[2359:2352]} - {1'b0, layer_0_0[2359:2352]};
      top_1[0] = {1'b0,layer_1_1[2343:2336]} - {1'b0, layer_0_1[2343:2336]};
      top_1[1] = {1'b0,layer_1_1[2351:2344]} - {1'b0, layer_0_1[2351:2344]};
      top_1[2] = {1'b0,layer_1_1[2359:2352]} - {1'b0, layer_0_1[2359:2352]};
      top_2[0] = {1'b0,layer_1_2[2343:2336]} - {1'b0, layer_0_2[2343:2336]};
      top_2[1] = {1'b0,layer_1_2[2351:2344]} - {1'b0, layer_0_2[2351:2344]};
      top_2[2] = {1'b0,layer_1_2[2359:2352]} - {1'b0, layer_0_2[2359:2352]};
      mid_0[0] = {1'b0,layer_2_0[2343:2336]} - {1'b0, layer_1_0[2343:2336]};
      mid_0[1] = {1'b0,layer_2_0[2351:2344]} - {1'b0, layer_1_0[2351:2344]};
      mid_0[2] = {1'b0,layer_2_0[2359:2352]} - {1'b0, layer_1_0[2359:2352]};
      mid_1[0] = {1'b0,layer_2_1[2343:2336]} - {1'b0, layer_1_1[2343:2336]};
      mid_1[1] = {1'b0,layer_2_1[2351:2344]} - {1'b0, layer_1_1[2351:2344]};
      mid_1[2] = {1'b0,layer_2_1[2359:2352]} - {1'b0, layer_1_1[2359:2352]};
      mid_2[0] = {1'b0,layer_2_2[2343:2336]} - {1'b0, layer_1_2[2343:2336]};
      mid_2[1] = {1'b0,layer_2_2[2351:2344]} - {1'b0, layer_1_2[2351:2344]};
      mid_2[2] = {1'b0,layer_2_2[2359:2352]} - {1'b0, layer_1_2[2359:2352]};
      btm_0[0] = {1'b0,layer_3_0[2343:2336]} - {1'b0, layer_2_0[2343:2336]};
      btm_0[1] = {1'b0,layer_3_0[2351:2344]} - {1'b0, layer_2_0[2351:2344]};
      btm_0[2] = {1'b0,layer_3_0[2359:2352]} - {1'b0, layer_2_0[2359:2352]};
      btm_1[0] = {1'b0,layer_3_1[2343:2336]} - {1'b0, layer_2_1[2343:2336]};
      btm_1[1] = {1'b0,layer_3_1[2351:2344]} - {1'b0, layer_2_1[2351:2344]};
      btm_1[2] = {1'b0,layer_3_1[2359:2352]} - {1'b0, layer_2_1[2359:2352]};
      btm_2[0] = {1'b0,layer_3_2[2343:2336]} - {1'b0, layer_2_2[2343:2336]};
      btm_2[1] = {1'b0,layer_3_2[2351:2344]} - {1'b0, layer_2_2[2351:2344]};
      btm_2[2] = {1'b0,layer_3_2[2359:2352]} - {1'b0, layer_2_2[2359:2352]};
    end
    'd294: begin
      top_0[0] = {1'b0,layer_1_0[2351:2344]} - {1'b0, layer_0_0[2351:2344]};
      top_0[1] = {1'b0,layer_1_0[2359:2352]} - {1'b0, layer_0_0[2359:2352]};
      top_0[2] = {1'b0,layer_1_0[2367:2360]} - {1'b0, layer_0_0[2367:2360]};
      top_1[0] = {1'b0,layer_1_1[2351:2344]} - {1'b0, layer_0_1[2351:2344]};
      top_1[1] = {1'b0,layer_1_1[2359:2352]} - {1'b0, layer_0_1[2359:2352]};
      top_1[2] = {1'b0,layer_1_1[2367:2360]} - {1'b0, layer_0_1[2367:2360]};
      top_2[0] = {1'b0,layer_1_2[2351:2344]} - {1'b0, layer_0_2[2351:2344]};
      top_2[1] = {1'b0,layer_1_2[2359:2352]} - {1'b0, layer_0_2[2359:2352]};
      top_2[2] = {1'b0,layer_1_2[2367:2360]} - {1'b0, layer_0_2[2367:2360]};
      mid_0[0] = {1'b0,layer_2_0[2351:2344]} - {1'b0, layer_1_0[2351:2344]};
      mid_0[1] = {1'b0,layer_2_0[2359:2352]} - {1'b0, layer_1_0[2359:2352]};
      mid_0[2] = {1'b0,layer_2_0[2367:2360]} - {1'b0, layer_1_0[2367:2360]};
      mid_1[0] = {1'b0,layer_2_1[2351:2344]} - {1'b0, layer_1_1[2351:2344]};
      mid_1[1] = {1'b0,layer_2_1[2359:2352]} - {1'b0, layer_1_1[2359:2352]};
      mid_1[2] = {1'b0,layer_2_1[2367:2360]} - {1'b0, layer_1_1[2367:2360]};
      mid_2[0] = {1'b0,layer_2_2[2351:2344]} - {1'b0, layer_1_2[2351:2344]};
      mid_2[1] = {1'b0,layer_2_2[2359:2352]} - {1'b0, layer_1_2[2359:2352]};
      mid_2[2] = {1'b0,layer_2_2[2367:2360]} - {1'b0, layer_1_2[2367:2360]};
      btm_0[0] = {1'b0,layer_3_0[2351:2344]} - {1'b0, layer_2_0[2351:2344]};
      btm_0[1] = {1'b0,layer_3_0[2359:2352]} - {1'b0, layer_2_0[2359:2352]};
      btm_0[2] = {1'b0,layer_3_0[2367:2360]} - {1'b0, layer_2_0[2367:2360]};
      btm_1[0] = {1'b0,layer_3_1[2351:2344]} - {1'b0, layer_2_1[2351:2344]};
      btm_1[1] = {1'b0,layer_3_1[2359:2352]} - {1'b0, layer_2_1[2359:2352]};
      btm_1[2] = {1'b0,layer_3_1[2367:2360]} - {1'b0, layer_2_1[2367:2360]};
      btm_2[0] = {1'b0,layer_3_2[2351:2344]} - {1'b0, layer_2_2[2351:2344]};
      btm_2[1] = {1'b0,layer_3_2[2359:2352]} - {1'b0, layer_2_2[2359:2352]};
      btm_2[2] = {1'b0,layer_3_2[2367:2360]} - {1'b0, layer_2_2[2367:2360]};
    end
    'd295: begin
      top_0[0] = {1'b0,layer_1_0[2359:2352]} - {1'b0, layer_0_0[2359:2352]};
      top_0[1] = {1'b0,layer_1_0[2367:2360]} - {1'b0, layer_0_0[2367:2360]};
      top_0[2] = {1'b0,layer_1_0[2375:2368]} - {1'b0, layer_0_0[2375:2368]};
      top_1[0] = {1'b0,layer_1_1[2359:2352]} - {1'b0, layer_0_1[2359:2352]};
      top_1[1] = {1'b0,layer_1_1[2367:2360]} - {1'b0, layer_0_1[2367:2360]};
      top_1[2] = {1'b0,layer_1_1[2375:2368]} - {1'b0, layer_0_1[2375:2368]};
      top_2[0] = {1'b0,layer_1_2[2359:2352]} - {1'b0, layer_0_2[2359:2352]};
      top_2[1] = {1'b0,layer_1_2[2367:2360]} - {1'b0, layer_0_2[2367:2360]};
      top_2[2] = {1'b0,layer_1_2[2375:2368]} - {1'b0, layer_0_2[2375:2368]};
      mid_0[0] = {1'b0,layer_2_0[2359:2352]} - {1'b0, layer_1_0[2359:2352]};
      mid_0[1] = {1'b0,layer_2_0[2367:2360]} - {1'b0, layer_1_0[2367:2360]};
      mid_0[2] = {1'b0,layer_2_0[2375:2368]} - {1'b0, layer_1_0[2375:2368]};
      mid_1[0] = {1'b0,layer_2_1[2359:2352]} - {1'b0, layer_1_1[2359:2352]};
      mid_1[1] = {1'b0,layer_2_1[2367:2360]} - {1'b0, layer_1_1[2367:2360]};
      mid_1[2] = {1'b0,layer_2_1[2375:2368]} - {1'b0, layer_1_1[2375:2368]};
      mid_2[0] = {1'b0,layer_2_2[2359:2352]} - {1'b0, layer_1_2[2359:2352]};
      mid_2[1] = {1'b0,layer_2_2[2367:2360]} - {1'b0, layer_1_2[2367:2360]};
      mid_2[2] = {1'b0,layer_2_2[2375:2368]} - {1'b0, layer_1_2[2375:2368]};
      btm_0[0] = {1'b0,layer_3_0[2359:2352]} - {1'b0, layer_2_0[2359:2352]};
      btm_0[1] = {1'b0,layer_3_0[2367:2360]} - {1'b0, layer_2_0[2367:2360]};
      btm_0[2] = {1'b0,layer_3_0[2375:2368]} - {1'b0, layer_2_0[2375:2368]};
      btm_1[0] = {1'b0,layer_3_1[2359:2352]} - {1'b0, layer_2_1[2359:2352]};
      btm_1[1] = {1'b0,layer_3_1[2367:2360]} - {1'b0, layer_2_1[2367:2360]};
      btm_1[2] = {1'b0,layer_3_1[2375:2368]} - {1'b0, layer_2_1[2375:2368]};
      btm_2[0] = {1'b0,layer_3_2[2359:2352]} - {1'b0, layer_2_2[2359:2352]};
      btm_2[1] = {1'b0,layer_3_2[2367:2360]} - {1'b0, layer_2_2[2367:2360]};
      btm_2[2] = {1'b0,layer_3_2[2375:2368]} - {1'b0, layer_2_2[2375:2368]};
    end
    'd296: begin
      top_0[0] = {1'b0,layer_1_0[2367:2360]} - {1'b0, layer_0_0[2367:2360]};
      top_0[1] = {1'b0,layer_1_0[2375:2368]} - {1'b0, layer_0_0[2375:2368]};
      top_0[2] = {1'b0,layer_1_0[2383:2376]} - {1'b0, layer_0_0[2383:2376]};
      top_1[0] = {1'b0,layer_1_1[2367:2360]} - {1'b0, layer_0_1[2367:2360]};
      top_1[1] = {1'b0,layer_1_1[2375:2368]} - {1'b0, layer_0_1[2375:2368]};
      top_1[2] = {1'b0,layer_1_1[2383:2376]} - {1'b0, layer_0_1[2383:2376]};
      top_2[0] = {1'b0,layer_1_2[2367:2360]} - {1'b0, layer_0_2[2367:2360]};
      top_2[1] = {1'b0,layer_1_2[2375:2368]} - {1'b0, layer_0_2[2375:2368]};
      top_2[2] = {1'b0,layer_1_2[2383:2376]} - {1'b0, layer_0_2[2383:2376]};
      mid_0[0] = {1'b0,layer_2_0[2367:2360]} - {1'b0, layer_1_0[2367:2360]};
      mid_0[1] = {1'b0,layer_2_0[2375:2368]} - {1'b0, layer_1_0[2375:2368]};
      mid_0[2] = {1'b0,layer_2_0[2383:2376]} - {1'b0, layer_1_0[2383:2376]};
      mid_1[0] = {1'b0,layer_2_1[2367:2360]} - {1'b0, layer_1_1[2367:2360]};
      mid_1[1] = {1'b0,layer_2_1[2375:2368]} - {1'b0, layer_1_1[2375:2368]};
      mid_1[2] = {1'b0,layer_2_1[2383:2376]} - {1'b0, layer_1_1[2383:2376]};
      mid_2[0] = {1'b0,layer_2_2[2367:2360]} - {1'b0, layer_1_2[2367:2360]};
      mid_2[1] = {1'b0,layer_2_2[2375:2368]} - {1'b0, layer_1_2[2375:2368]};
      mid_2[2] = {1'b0,layer_2_2[2383:2376]} - {1'b0, layer_1_2[2383:2376]};
      btm_0[0] = {1'b0,layer_3_0[2367:2360]} - {1'b0, layer_2_0[2367:2360]};
      btm_0[1] = {1'b0,layer_3_0[2375:2368]} - {1'b0, layer_2_0[2375:2368]};
      btm_0[2] = {1'b0,layer_3_0[2383:2376]} - {1'b0, layer_2_0[2383:2376]};
      btm_1[0] = {1'b0,layer_3_1[2367:2360]} - {1'b0, layer_2_1[2367:2360]};
      btm_1[1] = {1'b0,layer_3_1[2375:2368]} - {1'b0, layer_2_1[2375:2368]};
      btm_1[2] = {1'b0,layer_3_1[2383:2376]} - {1'b0, layer_2_1[2383:2376]};
      btm_2[0] = {1'b0,layer_3_2[2367:2360]} - {1'b0, layer_2_2[2367:2360]};
      btm_2[1] = {1'b0,layer_3_2[2375:2368]} - {1'b0, layer_2_2[2375:2368]};
      btm_2[2] = {1'b0,layer_3_2[2383:2376]} - {1'b0, layer_2_2[2383:2376]};
    end
    'd297: begin
      top_0[0] = {1'b0,layer_1_0[2375:2368]} - {1'b0, layer_0_0[2375:2368]};
      top_0[1] = {1'b0,layer_1_0[2383:2376]} - {1'b0, layer_0_0[2383:2376]};
      top_0[2] = {1'b0,layer_1_0[2391:2384]} - {1'b0, layer_0_0[2391:2384]};
      top_1[0] = {1'b0,layer_1_1[2375:2368]} - {1'b0, layer_0_1[2375:2368]};
      top_1[1] = {1'b0,layer_1_1[2383:2376]} - {1'b0, layer_0_1[2383:2376]};
      top_1[2] = {1'b0,layer_1_1[2391:2384]} - {1'b0, layer_0_1[2391:2384]};
      top_2[0] = {1'b0,layer_1_2[2375:2368]} - {1'b0, layer_0_2[2375:2368]};
      top_2[1] = {1'b0,layer_1_2[2383:2376]} - {1'b0, layer_0_2[2383:2376]};
      top_2[2] = {1'b0,layer_1_2[2391:2384]} - {1'b0, layer_0_2[2391:2384]};
      mid_0[0] = {1'b0,layer_2_0[2375:2368]} - {1'b0, layer_1_0[2375:2368]};
      mid_0[1] = {1'b0,layer_2_0[2383:2376]} - {1'b0, layer_1_0[2383:2376]};
      mid_0[2] = {1'b0,layer_2_0[2391:2384]} - {1'b0, layer_1_0[2391:2384]};
      mid_1[0] = {1'b0,layer_2_1[2375:2368]} - {1'b0, layer_1_1[2375:2368]};
      mid_1[1] = {1'b0,layer_2_1[2383:2376]} - {1'b0, layer_1_1[2383:2376]};
      mid_1[2] = {1'b0,layer_2_1[2391:2384]} - {1'b0, layer_1_1[2391:2384]};
      mid_2[0] = {1'b0,layer_2_2[2375:2368]} - {1'b0, layer_1_2[2375:2368]};
      mid_2[1] = {1'b0,layer_2_2[2383:2376]} - {1'b0, layer_1_2[2383:2376]};
      mid_2[2] = {1'b0,layer_2_2[2391:2384]} - {1'b0, layer_1_2[2391:2384]};
      btm_0[0] = {1'b0,layer_3_0[2375:2368]} - {1'b0, layer_2_0[2375:2368]};
      btm_0[1] = {1'b0,layer_3_0[2383:2376]} - {1'b0, layer_2_0[2383:2376]};
      btm_0[2] = {1'b0,layer_3_0[2391:2384]} - {1'b0, layer_2_0[2391:2384]};
      btm_1[0] = {1'b0,layer_3_1[2375:2368]} - {1'b0, layer_2_1[2375:2368]};
      btm_1[1] = {1'b0,layer_3_1[2383:2376]} - {1'b0, layer_2_1[2383:2376]};
      btm_1[2] = {1'b0,layer_3_1[2391:2384]} - {1'b0, layer_2_1[2391:2384]};
      btm_2[0] = {1'b0,layer_3_2[2375:2368]} - {1'b0, layer_2_2[2375:2368]};
      btm_2[1] = {1'b0,layer_3_2[2383:2376]} - {1'b0, layer_2_2[2383:2376]};
      btm_2[2] = {1'b0,layer_3_2[2391:2384]} - {1'b0, layer_2_2[2391:2384]};
    end
    'd298: begin
      top_0[0] = {1'b0,layer_1_0[2383:2376]} - {1'b0, layer_0_0[2383:2376]};
      top_0[1] = {1'b0,layer_1_0[2391:2384]} - {1'b0, layer_0_0[2391:2384]};
      top_0[2] = {1'b0,layer_1_0[2399:2392]} - {1'b0, layer_0_0[2399:2392]};
      top_1[0] = {1'b0,layer_1_1[2383:2376]} - {1'b0, layer_0_1[2383:2376]};
      top_1[1] = {1'b0,layer_1_1[2391:2384]} - {1'b0, layer_0_1[2391:2384]};
      top_1[2] = {1'b0,layer_1_1[2399:2392]} - {1'b0, layer_0_1[2399:2392]};
      top_2[0] = {1'b0,layer_1_2[2383:2376]} - {1'b0, layer_0_2[2383:2376]};
      top_2[1] = {1'b0,layer_1_2[2391:2384]} - {1'b0, layer_0_2[2391:2384]};
      top_2[2] = {1'b0,layer_1_2[2399:2392]} - {1'b0, layer_0_2[2399:2392]};
      mid_0[0] = {1'b0,layer_2_0[2383:2376]} - {1'b0, layer_1_0[2383:2376]};
      mid_0[1] = {1'b0,layer_2_0[2391:2384]} - {1'b0, layer_1_0[2391:2384]};
      mid_0[2] = {1'b0,layer_2_0[2399:2392]} - {1'b0, layer_1_0[2399:2392]};
      mid_1[0] = {1'b0,layer_2_1[2383:2376]} - {1'b0, layer_1_1[2383:2376]};
      mid_1[1] = {1'b0,layer_2_1[2391:2384]} - {1'b0, layer_1_1[2391:2384]};
      mid_1[2] = {1'b0,layer_2_1[2399:2392]} - {1'b0, layer_1_1[2399:2392]};
      mid_2[0] = {1'b0,layer_2_2[2383:2376]} - {1'b0, layer_1_2[2383:2376]};
      mid_2[1] = {1'b0,layer_2_2[2391:2384]} - {1'b0, layer_1_2[2391:2384]};
      mid_2[2] = {1'b0,layer_2_2[2399:2392]} - {1'b0, layer_1_2[2399:2392]};
      btm_0[0] = {1'b0,layer_3_0[2383:2376]} - {1'b0, layer_2_0[2383:2376]};
      btm_0[1] = {1'b0,layer_3_0[2391:2384]} - {1'b0, layer_2_0[2391:2384]};
      btm_0[2] = {1'b0,layer_3_0[2399:2392]} - {1'b0, layer_2_0[2399:2392]};
      btm_1[0] = {1'b0,layer_3_1[2383:2376]} - {1'b0, layer_2_1[2383:2376]};
      btm_1[1] = {1'b0,layer_3_1[2391:2384]} - {1'b0, layer_2_1[2391:2384]};
      btm_1[2] = {1'b0,layer_3_1[2399:2392]} - {1'b0, layer_2_1[2399:2392]};
      btm_2[0] = {1'b0,layer_3_2[2383:2376]} - {1'b0, layer_2_2[2383:2376]};
      btm_2[1] = {1'b0,layer_3_2[2391:2384]} - {1'b0, layer_2_2[2391:2384]};
      btm_2[2] = {1'b0,layer_3_2[2399:2392]} - {1'b0, layer_2_2[2399:2392]};
    end
    'd299: begin
      top_0[0] = {1'b0,layer_1_0[2391:2384]} - {1'b0, layer_0_0[2391:2384]};
      top_0[1] = {1'b0,layer_1_0[2399:2392]} - {1'b0, layer_0_0[2399:2392]};
      top_0[2] = {1'b0,layer_1_0[2407:2400]} - {1'b0, layer_0_0[2407:2400]};
      top_1[0] = {1'b0,layer_1_1[2391:2384]} - {1'b0, layer_0_1[2391:2384]};
      top_1[1] = {1'b0,layer_1_1[2399:2392]} - {1'b0, layer_0_1[2399:2392]};
      top_1[2] = {1'b0,layer_1_1[2407:2400]} - {1'b0, layer_0_1[2407:2400]};
      top_2[0] = {1'b0,layer_1_2[2391:2384]} - {1'b0, layer_0_2[2391:2384]};
      top_2[1] = {1'b0,layer_1_2[2399:2392]} - {1'b0, layer_0_2[2399:2392]};
      top_2[2] = {1'b0,layer_1_2[2407:2400]} - {1'b0, layer_0_2[2407:2400]};
      mid_0[0] = {1'b0,layer_2_0[2391:2384]} - {1'b0, layer_1_0[2391:2384]};
      mid_0[1] = {1'b0,layer_2_0[2399:2392]} - {1'b0, layer_1_0[2399:2392]};
      mid_0[2] = {1'b0,layer_2_0[2407:2400]} - {1'b0, layer_1_0[2407:2400]};
      mid_1[0] = {1'b0,layer_2_1[2391:2384]} - {1'b0, layer_1_1[2391:2384]};
      mid_1[1] = {1'b0,layer_2_1[2399:2392]} - {1'b0, layer_1_1[2399:2392]};
      mid_1[2] = {1'b0,layer_2_1[2407:2400]} - {1'b0, layer_1_1[2407:2400]};
      mid_2[0] = {1'b0,layer_2_2[2391:2384]} - {1'b0, layer_1_2[2391:2384]};
      mid_2[1] = {1'b0,layer_2_2[2399:2392]} - {1'b0, layer_1_2[2399:2392]};
      mid_2[2] = {1'b0,layer_2_2[2407:2400]} - {1'b0, layer_1_2[2407:2400]};
      btm_0[0] = {1'b0,layer_3_0[2391:2384]} - {1'b0, layer_2_0[2391:2384]};
      btm_0[1] = {1'b0,layer_3_0[2399:2392]} - {1'b0, layer_2_0[2399:2392]};
      btm_0[2] = {1'b0,layer_3_0[2407:2400]} - {1'b0, layer_2_0[2407:2400]};
      btm_1[0] = {1'b0,layer_3_1[2391:2384]} - {1'b0, layer_2_1[2391:2384]};
      btm_1[1] = {1'b0,layer_3_1[2399:2392]} - {1'b0, layer_2_1[2399:2392]};
      btm_1[2] = {1'b0,layer_3_1[2407:2400]} - {1'b0, layer_2_1[2407:2400]};
      btm_2[0] = {1'b0,layer_3_2[2391:2384]} - {1'b0, layer_2_2[2391:2384]};
      btm_2[1] = {1'b0,layer_3_2[2399:2392]} - {1'b0, layer_2_2[2399:2392]};
      btm_2[2] = {1'b0,layer_3_2[2407:2400]} - {1'b0, layer_2_2[2407:2400]};
    end
    'd300: begin
      top_0[0] = {1'b0,layer_1_0[2399:2392]} - {1'b0, layer_0_0[2399:2392]};
      top_0[1] = {1'b0,layer_1_0[2407:2400]} - {1'b0, layer_0_0[2407:2400]};
      top_0[2] = {1'b0,layer_1_0[2415:2408]} - {1'b0, layer_0_0[2415:2408]};
      top_1[0] = {1'b0,layer_1_1[2399:2392]} - {1'b0, layer_0_1[2399:2392]};
      top_1[1] = {1'b0,layer_1_1[2407:2400]} - {1'b0, layer_0_1[2407:2400]};
      top_1[2] = {1'b0,layer_1_1[2415:2408]} - {1'b0, layer_0_1[2415:2408]};
      top_2[0] = {1'b0,layer_1_2[2399:2392]} - {1'b0, layer_0_2[2399:2392]};
      top_2[1] = {1'b0,layer_1_2[2407:2400]} - {1'b0, layer_0_2[2407:2400]};
      top_2[2] = {1'b0,layer_1_2[2415:2408]} - {1'b0, layer_0_2[2415:2408]};
      mid_0[0] = {1'b0,layer_2_0[2399:2392]} - {1'b0, layer_1_0[2399:2392]};
      mid_0[1] = {1'b0,layer_2_0[2407:2400]} - {1'b0, layer_1_0[2407:2400]};
      mid_0[2] = {1'b0,layer_2_0[2415:2408]} - {1'b0, layer_1_0[2415:2408]};
      mid_1[0] = {1'b0,layer_2_1[2399:2392]} - {1'b0, layer_1_1[2399:2392]};
      mid_1[1] = {1'b0,layer_2_1[2407:2400]} - {1'b0, layer_1_1[2407:2400]};
      mid_1[2] = {1'b0,layer_2_1[2415:2408]} - {1'b0, layer_1_1[2415:2408]};
      mid_2[0] = {1'b0,layer_2_2[2399:2392]} - {1'b0, layer_1_2[2399:2392]};
      mid_2[1] = {1'b0,layer_2_2[2407:2400]} - {1'b0, layer_1_2[2407:2400]};
      mid_2[2] = {1'b0,layer_2_2[2415:2408]} - {1'b0, layer_1_2[2415:2408]};
      btm_0[0] = {1'b0,layer_3_0[2399:2392]} - {1'b0, layer_2_0[2399:2392]};
      btm_0[1] = {1'b0,layer_3_0[2407:2400]} - {1'b0, layer_2_0[2407:2400]};
      btm_0[2] = {1'b0,layer_3_0[2415:2408]} - {1'b0, layer_2_0[2415:2408]};
      btm_1[0] = {1'b0,layer_3_1[2399:2392]} - {1'b0, layer_2_1[2399:2392]};
      btm_1[1] = {1'b0,layer_3_1[2407:2400]} - {1'b0, layer_2_1[2407:2400]};
      btm_1[2] = {1'b0,layer_3_1[2415:2408]} - {1'b0, layer_2_1[2415:2408]};
      btm_2[0] = {1'b0,layer_3_2[2399:2392]} - {1'b0, layer_2_2[2399:2392]};
      btm_2[1] = {1'b0,layer_3_2[2407:2400]} - {1'b0, layer_2_2[2407:2400]};
      btm_2[2] = {1'b0,layer_3_2[2415:2408]} - {1'b0, layer_2_2[2415:2408]};
    end
    'd301: begin
      top_0[0] = {1'b0,layer_1_0[2407:2400]} - {1'b0, layer_0_0[2407:2400]};
      top_0[1] = {1'b0,layer_1_0[2415:2408]} - {1'b0, layer_0_0[2415:2408]};
      top_0[2] = {1'b0,layer_1_0[2423:2416]} - {1'b0, layer_0_0[2423:2416]};
      top_1[0] = {1'b0,layer_1_1[2407:2400]} - {1'b0, layer_0_1[2407:2400]};
      top_1[1] = {1'b0,layer_1_1[2415:2408]} - {1'b0, layer_0_1[2415:2408]};
      top_1[2] = {1'b0,layer_1_1[2423:2416]} - {1'b0, layer_0_1[2423:2416]};
      top_2[0] = {1'b0,layer_1_2[2407:2400]} - {1'b0, layer_0_2[2407:2400]};
      top_2[1] = {1'b0,layer_1_2[2415:2408]} - {1'b0, layer_0_2[2415:2408]};
      top_2[2] = {1'b0,layer_1_2[2423:2416]} - {1'b0, layer_0_2[2423:2416]};
      mid_0[0] = {1'b0,layer_2_0[2407:2400]} - {1'b0, layer_1_0[2407:2400]};
      mid_0[1] = {1'b0,layer_2_0[2415:2408]} - {1'b0, layer_1_0[2415:2408]};
      mid_0[2] = {1'b0,layer_2_0[2423:2416]} - {1'b0, layer_1_0[2423:2416]};
      mid_1[0] = {1'b0,layer_2_1[2407:2400]} - {1'b0, layer_1_1[2407:2400]};
      mid_1[1] = {1'b0,layer_2_1[2415:2408]} - {1'b0, layer_1_1[2415:2408]};
      mid_1[2] = {1'b0,layer_2_1[2423:2416]} - {1'b0, layer_1_1[2423:2416]};
      mid_2[0] = {1'b0,layer_2_2[2407:2400]} - {1'b0, layer_1_2[2407:2400]};
      mid_2[1] = {1'b0,layer_2_2[2415:2408]} - {1'b0, layer_1_2[2415:2408]};
      mid_2[2] = {1'b0,layer_2_2[2423:2416]} - {1'b0, layer_1_2[2423:2416]};
      btm_0[0] = {1'b0,layer_3_0[2407:2400]} - {1'b0, layer_2_0[2407:2400]};
      btm_0[1] = {1'b0,layer_3_0[2415:2408]} - {1'b0, layer_2_0[2415:2408]};
      btm_0[2] = {1'b0,layer_3_0[2423:2416]} - {1'b0, layer_2_0[2423:2416]};
      btm_1[0] = {1'b0,layer_3_1[2407:2400]} - {1'b0, layer_2_1[2407:2400]};
      btm_1[1] = {1'b0,layer_3_1[2415:2408]} - {1'b0, layer_2_1[2415:2408]};
      btm_1[2] = {1'b0,layer_3_1[2423:2416]} - {1'b0, layer_2_1[2423:2416]};
      btm_2[0] = {1'b0,layer_3_2[2407:2400]} - {1'b0, layer_2_2[2407:2400]};
      btm_2[1] = {1'b0,layer_3_2[2415:2408]} - {1'b0, layer_2_2[2415:2408]};
      btm_2[2] = {1'b0,layer_3_2[2423:2416]} - {1'b0, layer_2_2[2423:2416]};
    end
    'd302: begin
      top_0[0] = {1'b0,layer_1_0[2415:2408]} - {1'b0, layer_0_0[2415:2408]};
      top_0[1] = {1'b0,layer_1_0[2423:2416]} - {1'b0, layer_0_0[2423:2416]};
      top_0[2] = {1'b0,layer_1_0[2431:2424]} - {1'b0, layer_0_0[2431:2424]};
      top_1[0] = {1'b0,layer_1_1[2415:2408]} - {1'b0, layer_0_1[2415:2408]};
      top_1[1] = {1'b0,layer_1_1[2423:2416]} - {1'b0, layer_0_1[2423:2416]};
      top_1[2] = {1'b0,layer_1_1[2431:2424]} - {1'b0, layer_0_1[2431:2424]};
      top_2[0] = {1'b0,layer_1_2[2415:2408]} - {1'b0, layer_0_2[2415:2408]};
      top_2[1] = {1'b0,layer_1_2[2423:2416]} - {1'b0, layer_0_2[2423:2416]};
      top_2[2] = {1'b0,layer_1_2[2431:2424]} - {1'b0, layer_0_2[2431:2424]};
      mid_0[0] = {1'b0,layer_2_0[2415:2408]} - {1'b0, layer_1_0[2415:2408]};
      mid_0[1] = {1'b0,layer_2_0[2423:2416]} - {1'b0, layer_1_0[2423:2416]};
      mid_0[2] = {1'b0,layer_2_0[2431:2424]} - {1'b0, layer_1_0[2431:2424]};
      mid_1[0] = {1'b0,layer_2_1[2415:2408]} - {1'b0, layer_1_1[2415:2408]};
      mid_1[1] = {1'b0,layer_2_1[2423:2416]} - {1'b0, layer_1_1[2423:2416]};
      mid_1[2] = {1'b0,layer_2_1[2431:2424]} - {1'b0, layer_1_1[2431:2424]};
      mid_2[0] = {1'b0,layer_2_2[2415:2408]} - {1'b0, layer_1_2[2415:2408]};
      mid_2[1] = {1'b0,layer_2_2[2423:2416]} - {1'b0, layer_1_2[2423:2416]};
      mid_2[2] = {1'b0,layer_2_2[2431:2424]} - {1'b0, layer_1_2[2431:2424]};
      btm_0[0] = {1'b0,layer_3_0[2415:2408]} - {1'b0, layer_2_0[2415:2408]};
      btm_0[1] = {1'b0,layer_3_0[2423:2416]} - {1'b0, layer_2_0[2423:2416]};
      btm_0[2] = {1'b0,layer_3_0[2431:2424]} - {1'b0, layer_2_0[2431:2424]};
      btm_1[0] = {1'b0,layer_3_1[2415:2408]} - {1'b0, layer_2_1[2415:2408]};
      btm_1[1] = {1'b0,layer_3_1[2423:2416]} - {1'b0, layer_2_1[2423:2416]};
      btm_1[2] = {1'b0,layer_3_1[2431:2424]} - {1'b0, layer_2_1[2431:2424]};
      btm_2[0] = {1'b0,layer_3_2[2415:2408]} - {1'b0, layer_2_2[2415:2408]};
      btm_2[1] = {1'b0,layer_3_2[2423:2416]} - {1'b0, layer_2_2[2423:2416]};
      btm_2[2] = {1'b0,layer_3_2[2431:2424]} - {1'b0, layer_2_2[2431:2424]};
    end
    'd303: begin
      top_0[0] = {1'b0,layer_1_0[2423:2416]} - {1'b0, layer_0_0[2423:2416]};
      top_0[1] = {1'b0,layer_1_0[2431:2424]} - {1'b0, layer_0_0[2431:2424]};
      top_0[2] = {1'b0,layer_1_0[2439:2432]} - {1'b0, layer_0_0[2439:2432]};
      top_1[0] = {1'b0,layer_1_1[2423:2416]} - {1'b0, layer_0_1[2423:2416]};
      top_1[1] = {1'b0,layer_1_1[2431:2424]} - {1'b0, layer_0_1[2431:2424]};
      top_1[2] = {1'b0,layer_1_1[2439:2432]} - {1'b0, layer_0_1[2439:2432]};
      top_2[0] = {1'b0,layer_1_2[2423:2416]} - {1'b0, layer_0_2[2423:2416]};
      top_2[1] = {1'b0,layer_1_2[2431:2424]} - {1'b0, layer_0_2[2431:2424]};
      top_2[2] = {1'b0,layer_1_2[2439:2432]} - {1'b0, layer_0_2[2439:2432]};
      mid_0[0] = {1'b0,layer_2_0[2423:2416]} - {1'b0, layer_1_0[2423:2416]};
      mid_0[1] = {1'b0,layer_2_0[2431:2424]} - {1'b0, layer_1_0[2431:2424]};
      mid_0[2] = {1'b0,layer_2_0[2439:2432]} - {1'b0, layer_1_0[2439:2432]};
      mid_1[0] = {1'b0,layer_2_1[2423:2416]} - {1'b0, layer_1_1[2423:2416]};
      mid_1[1] = {1'b0,layer_2_1[2431:2424]} - {1'b0, layer_1_1[2431:2424]};
      mid_1[2] = {1'b0,layer_2_1[2439:2432]} - {1'b0, layer_1_1[2439:2432]};
      mid_2[0] = {1'b0,layer_2_2[2423:2416]} - {1'b0, layer_1_2[2423:2416]};
      mid_2[1] = {1'b0,layer_2_2[2431:2424]} - {1'b0, layer_1_2[2431:2424]};
      mid_2[2] = {1'b0,layer_2_2[2439:2432]} - {1'b0, layer_1_2[2439:2432]};
      btm_0[0] = {1'b0,layer_3_0[2423:2416]} - {1'b0, layer_2_0[2423:2416]};
      btm_0[1] = {1'b0,layer_3_0[2431:2424]} - {1'b0, layer_2_0[2431:2424]};
      btm_0[2] = {1'b0,layer_3_0[2439:2432]} - {1'b0, layer_2_0[2439:2432]};
      btm_1[0] = {1'b0,layer_3_1[2423:2416]} - {1'b0, layer_2_1[2423:2416]};
      btm_1[1] = {1'b0,layer_3_1[2431:2424]} - {1'b0, layer_2_1[2431:2424]};
      btm_1[2] = {1'b0,layer_3_1[2439:2432]} - {1'b0, layer_2_1[2439:2432]};
      btm_2[0] = {1'b0,layer_3_2[2423:2416]} - {1'b0, layer_2_2[2423:2416]};
      btm_2[1] = {1'b0,layer_3_2[2431:2424]} - {1'b0, layer_2_2[2431:2424]};
      btm_2[2] = {1'b0,layer_3_2[2439:2432]} - {1'b0, layer_2_2[2439:2432]};
    end
    'd304: begin
      top_0[0] = {1'b0,layer_1_0[2431:2424]} - {1'b0, layer_0_0[2431:2424]};
      top_0[1] = {1'b0,layer_1_0[2439:2432]} - {1'b0, layer_0_0[2439:2432]};
      top_0[2] = {1'b0,layer_1_0[2447:2440]} - {1'b0, layer_0_0[2447:2440]};
      top_1[0] = {1'b0,layer_1_1[2431:2424]} - {1'b0, layer_0_1[2431:2424]};
      top_1[1] = {1'b0,layer_1_1[2439:2432]} - {1'b0, layer_0_1[2439:2432]};
      top_1[2] = {1'b0,layer_1_1[2447:2440]} - {1'b0, layer_0_1[2447:2440]};
      top_2[0] = {1'b0,layer_1_2[2431:2424]} - {1'b0, layer_0_2[2431:2424]};
      top_2[1] = {1'b0,layer_1_2[2439:2432]} - {1'b0, layer_0_2[2439:2432]};
      top_2[2] = {1'b0,layer_1_2[2447:2440]} - {1'b0, layer_0_2[2447:2440]};
      mid_0[0] = {1'b0,layer_2_0[2431:2424]} - {1'b0, layer_1_0[2431:2424]};
      mid_0[1] = {1'b0,layer_2_0[2439:2432]} - {1'b0, layer_1_0[2439:2432]};
      mid_0[2] = {1'b0,layer_2_0[2447:2440]} - {1'b0, layer_1_0[2447:2440]};
      mid_1[0] = {1'b0,layer_2_1[2431:2424]} - {1'b0, layer_1_1[2431:2424]};
      mid_1[1] = {1'b0,layer_2_1[2439:2432]} - {1'b0, layer_1_1[2439:2432]};
      mid_1[2] = {1'b0,layer_2_1[2447:2440]} - {1'b0, layer_1_1[2447:2440]};
      mid_2[0] = {1'b0,layer_2_2[2431:2424]} - {1'b0, layer_1_2[2431:2424]};
      mid_2[1] = {1'b0,layer_2_2[2439:2432]} - {1'b0, layer_1_2[2439:2432]};
      mid_2[2] = {1'b0,layer_2_2[2447:2440]} - {1'b0, layer_1_2[2447:2440]};
      btm_0[0] = {1'b0,layer_3_0[2431:2424]} - {1'b0, layer_2_0[2431:2424]};
      btm_0[1] = {1'b0,layer_3_0[2439:2432]} - {1'b0, layer_2_0[2439:2432]};
      btm_0[2] = {1'b0,layer_3_0[2447:2440]} - {1'b0, layer_2_0[2447:2440]};
      btm_1[0] = {1'b0,layer_3_1[2431:2424]} - {1'b0, layer_2_1[2431:2424]};
      btm_1[1] = {1'b0,layer_3_1[2439:2432]} - {1'b0, layer_2_1[2439:2432]};
      btm_1[2] = {1'b0,layer_3_1[2447:2440]} - {1'b0, layer_2_1[2447:2440]};
      btm_2[0] = {1'b0,layer_3_2[2431:2424]} - {1'b0, layer_2_2[2431:2424]};
      btm_2[1] = {1'b0,layer_3_2[2439:2432]} - {1'b0, layer_2_2[2439:2432]};
      btm_2[2] = {1'b0,layer_3_2[2447:2440]} - {1'b0, layer_2_2[2447:2440]};
    end
    'd305: begin
      top_0[0] = {1'b0,layer_1_0[2439:2432]} - {1'b0, layer_0_0[2439:2432]};
      top_0[1] = {1'b0,layer_1_0[2447:2440]} - {1'b0, layer_0_0[2447:2440]};
      top_0[2] = {1'b0,layer_1_0[2455:2448]} - {1'b0, layer_0_0[2455:2448]};
      top_1[0] = {1'b0,layer_1_1[2439:2432]} - {1'b0, layer_0_1[2439:2432]};
      top_1[1] = {1'b0,layer_1_1[2447:2440]} - {1'b0, layer_0_1[2447:2440]};
      top_1[2] = {1'b0,layer_1_1[2455:2448]} - {1'b0, layer_0_1[2455:2448]};
      top_2[0] = {1'b0,layer_1_2[2439:2432]} - {1'b0, layer_0_2[2439:2432]};
      top_2[1] = {1'b0,layer_1_2[2447:2440]} - {1'b0, layer_0_2[2447:2440]};
      top_2[2] = {1'b0,layer_1_2[2455:2448]} - {1'b0, layer_0_2[2455:2448]};
      mid_0[0] = {1'b0,layer_2_0[2439:2432]} - {1'b0, layer_1_0[2439:2432]};
      mid_0[1] = {1'b0,layer_2_0[2447:2440]} - {1'b0, layer_1_0[2447:2440]};
      mid_0[2] = {1'b0,layer_2_0[2455:2448]} - {1'b0, layer_1_0[2455:2448]};
      mid_1[0] = {1'b0,layer_2_1[2439:2432]} - {1'b0, layer_1_1[2439:2432]};
      mid_1[1] = {1'b0,layer_2_1[2447:2440]} - {1'b0, layer_1_1[2447:2440]};
      mid_1[2] = {1'b0,layer_2_1[2455:2448]} - {1'b0, layer_1_1[2455:2448]};
      mid_2[0] = {1'b0,layer_2_2[2439:2432]} - {1'b0, layer_1_2[2439:2432]};
      mid_2[1] = {1'b0,layer_2_2[2447:2440]} - {1'b0, layer_1_2[2447:2440]};
      mid_2[2] = {1'b0,layer_2_2[2455:2448]} - {1'b0, layer_1_2[2455:2448]};
      btm_0[0] = {1'b0,layer_3_0[2439:2432]} - {1'b0, layer_2_0[2439:2432]};
      btm_0[1] = {1'b0,layer_3_0[2447:2440]} - {1'b0, layer_2_0[2447:2440]};
      btm_0[2] = {1'b0,layer_3_0[2455:2448]} - {1'b0, layer_2_0[2455:2448]};
      btm_1[0] = {1'b0,layer_3_1[2439:2432]} - {1'b0, layer_2_1[2439:2432]};
      btm_1[1] = {1'b0,layer_3_1[2447:2440]} - {1'b0, layer_2_1[2447:2440]};
      btm_1[2] = {1'b0,layer_3_1[2455:2448]} - {1'b0, layer_2_1[2455:2448]};
      btm_2[0] = {1'b0,layer_3_2[2439:2432]} - {1'b0, layer_2_2[2439:2432]};
      btm_2[1] = {1'b0,layer_3_2[2447:2440]} - {1'b0, layer_2_2[2447:2440]};
      btm_2[2] = {1'b0,layer_3_2[2455:2448]} - {1'b0, layer_2_2[2455:2448]};
    end
    'd306: begin
      top_0[0] = {1'b0,layer_1_0[2447:2440]} - {1'b0, layer_0_0[2447:2440]};
      top_0[1] = {1'b0,layer_1_0[2455:2448]} - {1'b0, layer_0_0[2455:2448]};
      top_0[2] = {1'b0,layer_1_0[2463:2456]} - {1'b0, layer_0_0[2463:2456]};
      top_1[0] = {1'b0,layer_1_1[2447:2440]} - {1'b0, layer_0_1[2447:2440]};
      top_1[1] = {1'b0,layer_1_1[2455:2448]} - {1'b0, layer_0_1[2455:2448]};
      top_1[2] = {1'b0,layer_1_1[2463:2456]} - {1'b0, layer_0_1[2463:2456]};
      top_2[0] = {1'b0,layer_1_2[2447:2440]} - {1'b0, layer_0_2[2447:2440]};
      top_2[1] = {1'b0,layer_1_2[2455:2448]} - {1'b0, layer_0_2[2455:2448]};
      top_2[2] = {1'b0,layer_1_2[2463:2456]} - {1'b0, layer_0_2[2463:2456]};
      mid_0[0] = {1'b0,layer_2_0[2447:2440]} - {1'b0, layer_1_0[2447:2440]};
      mid_0[1] = {1'b0,layer_2_0[2455:2448]} - {1'b0, layer_1_0[2455:2448]};
      mid_0[2] = {1'b0,layer_2_0[2463:2456]} - {1'b0, layer_1_0[2463:2456]};
      mid_1[0] = {1'b0,layer_2_1[2447:2440]} - {1'b0, layer_1_1[2447:2440]};
      mid_1[1] = {1'b0,layer_2_1[2455:2448]} - {1'b0, layer_1_1[2455:2448]};
      mid_1[2] = {1'b0,layer_2_1[2463:2456]} - {1'b0, layer_1_1[2463:2456]};
      mid_2[0] = {1'b0,layer_2_2[2447:2440]} - {1'b0, layer_1_2[2447:2440]};
      mid_2[1] = {1'b0,layer_2_2[2455:2448]} - {1'b0, layer_1_2[2455:2448]};
      mid_2[2] = {1'b0,layer_2_2[2463:2456]} - {1'b0, layer_1_2[2463:2456]};
      btm_0[0] = {1'b0,layer_3_0[2447:2440]} - {1'b0, layer_2_0[2447:2440]};
      btm_0[1] = {1'b0,layer_3_0[2455:2448]} - {1'b0, layer_2_0[2455:2448]};
      btm_0[2] = {1'b0,layer_3_0[2463:2456]} - {1'b0, layer_2_0[2463:2456]};
      btm_1[0] = {1'b0,layer_3_1[2447:2440]} - {1'b0, layer_2_1[2447:2440]};
      btm_1[1] = {1'b0,layer_3_1[2455:2448]} - {1'b0, layer_2_1[2455:2448]};
      btm_1[2] = {1'b0,layer_3_1[2463:2456]} - {1'b0, layer_2_1[2463:2456]};
      btm_2[0] = {1'b0,layer_3_2[2447:2440]} - {1'b0, layer_2_2[2447:2440]};
      btm_2[1] = {1'b0,layer_3_2[2455:2448]} - {1'b0, layer_2_2[2455:2448]};
      btm_2[2] = {1'b0,layer_3_2[2463:2456]} - {1'b0, layer_2_2[2463:2456]};
    end
    'd307: begin
      top_0[0] = {1'b0,layer_1_0[2455:2448]} - {1'b0, layer_0_0[2455:2448]};
      top_0[1] = {1'b0,layer_1_0[2463:2456]} - {1'b0, layer_0_0[2463:2456]};
      top_0[2] = {1'b0,layer_1_0[2471:2464]} - {1'b0, layer_0_0[2471:2464]};
      top_1[0] = {1'b0,layer_1_1[2455:2448]} - {1'b0, layer_0_1[2455:2448]};
      top_1[1] = {1'b0,layer_1_1[2463:2456]} - {1'b0, layer_0_1[2463:2456]};
      top_1[2] = {1'b0,layer_1_1[2471:2464]} - {1'b0, layer_0_1[2471:2464]};
      top_2[0] = {1'b0,layer_1_2[2455:2448]} - {1'b0, layer_0_2[2455:2448]};
      top_2[1] = {1'b0,layer_1_2[2463:2456]} - {1'b0, layer_0_2[2463:2456]};
      top_2[2] = {1'b0,layer_1_2[2471:2464]} - {1'b0, layer_0_2[2471:2464]};
      mid_0[0] = {1'b0,layer_2_0[2455:2448]} - {1'b0, layer_1_0[2455:2448]};
      mid_0[1] = {1'b0,layer_2_0[2463:2456]} - {1'b0, layer_1_0[2463:2456]};
      mid_0[2] = {1'b0,layer_2_0[2471:2464]} - {1'b0, layer_1_0[2471:2464]};
      mid_1[0] = {1'b0,layer_2_1[2455:2448]} - {1'b0, layer_1_1[2455:2448]};
      mid_1[1] = {1'b0,layer_2_1[2463:2456]} - {1'b0, layer_1_1[2463:2456]};
      mid_1[2] = {1'b0,layer_2_1[2471:2464]} - {1'b0, layer_1_1[2471:2464]};
      mid_2[0] = {1'b0,layer_2_2[2455:2448]} - {1'b0, layer_1_2[2455:2448]};
      mid_2[1] = {1'b0,layer_2_2[2463:2456]} - {1'b0, layer_1_2[2463:2456]};
      mid_2[2] = {1'b0,layer_2_2[2471:2464]} - {1'b0, layer_1_2[2471:2464]};
      btm_0[0] = {1'b0,layer_3_0[2455:2448]} - {1'b0, layer_2_0[2455:2448]};
      btm_0[1] = {1'b0,layer_3_0[2463:2456]} - {1'b0, layer_2_0[2463:2456]};
      btm_0[2] = {1'b0,layer_3_0[2471:2464]} - {1'b0, layer_2_0[2471:2464]};
      btm_1[0] = {1'b0,layer_3_1[2455:2448]} - {1'b0, layer_2_1[2455:2448]};
      btm_1[1] = {1'b0,layer_3_1[2463:2456]} - {1'b0, layer_2_1[2463:2456]};
      btm_1[2] = {1'b0,layer_3_1[2471:2464]} - {1'b0, layer_2_1[2471:2464]};
      btm_2[0] = {1'b0,layer_3_2[2455:2448]} - {1'b0, layer_2_2[2455:2448]};
      btm_2[1] = {1'b0,layer_3_2[2463:2456]} - {1'b0, layer_2_2[2463:2456]};
      btm_2[2] = {1'b0,layer_3_2[2471:2464]} - {1'b0, layer_2_2[2471:2464]};
    end
    'd308: begin
      top_0[0] = {1'b0,layer_1_0[2463:2456]} - {1'b0, layer_0_0[2463:2456]};
      top_0[1] = {1'b0,layer_1_0[2471:2464]} - {1'b0, layer_0_0[2471:2464]};
      top_0[2] = {1'b0,layer_1_0[2479:2472]} - {1'b0, layer_0_0[2479:2472]};
      top_1[0] = {1'b0,layer_1_1[2463:2456]} - {1'b0, layer_0_1[2463:2456]};
      top_1[1] = {1'b0,layer_1_1[2471:2464]} - {1'b0, layer_0_1[2471:2464]};
      top_1[2] = {1'b0,layer_1_1[2479:2472]} - {1'b0, layer_0_1[2479:2472]};
      top_2[0] = {1'b0,layer_1_2[2463:2456]} - {1'b0, layer_0_2[2463:2456]};
      top_2[1] = {1'b0,layer_1_2[2471:2464]} - {1'b0, layer_0_2[2471:2464]};
      top_2[2] = {1'b0,layer_1_2[2479:2472]} - {1'b0, layer_0_2[2479:2472]};
      mid_0[0] = {1'b0,layer_2_0[2463:2456]} - {1'b0, layer_1_0[2463:2456]};
      mid_0[1] = {1'b0,layer_2_0[2471:2464]} - {1'b0, layer_1_0[2471:2464]};
      mid_0[2] = {1'b0,layer_2_0[2479:2472]} - {1'b0, layer_1_0[2479:2472]};
      mid_1[0] = {1'b0,layer_2_1[2463:2456]} - {1'b0, layer_1_1[2463:2456]};
      mid_1[1] = {1'b0,layer_2_1[2471:2464]} - {1'b0, layer_1_1[2471:2464]};
      mid_1[2] = {1'b0,layer_2_1[2479:2472]} - {1'b0, layer_1_1[2479:2472]};
      mid_2[0] = {1'b0,layer_2_2[2463:2456]} - {1'b0, layer_1_2[2463:2456]};
      mid_2[1] = {1'b0,layer_2_2[2471:2464]} - {1'b0, layer_1_2[2471:2464]};
      mid_2[2] = {1'b0,layer_2_2[2479:2472]} - {1'b0, layer_1_2[2479:2472]};
      btm_0[0] = {1'b0,layer_3_0[2463:2456]} - {1'b0, layer_2_0[2463:2456]};
      btm_0[1] = {1'b0,layer_3_0[2471:2464]} - {1'b0, layer_2_0[2471:2464]};
      btm_0[2] = {1'b0,layer_3_0[2479:2472]} - {1'b0, layer_2_0[2479:2472]};
      btm_1[0] = {1'b0,layer_3_1[2463:2456]} - {1'b0, layer_2_1[2463:2456]};
      btm_1[1] = {1'b0,layer_3_1[2471:2464]} - {1'b0, layer_2_1[2471:2464]};
      btm_1[2] = {1'b0,layer_3_1[2479:2472]} - {1'b0, layer_2_1[2479:2472]};
      btm_2[0] = {1'b0,layer_3_2[2463:2456]} - {1'b0, layer_2_2[2463:2456]};
      btm_2[1] = {1'b0,layer_3_2[2471:2464]} - {1'b0, layer_2_2[2471:2464]};
      btm_2[2] = {1'b0,layer_3_2[2479:2472]} - {1'b0, layer_2_2[2479:2472]};
    end
    'd309: begin
      top_0[0] = {1'b0,layer_1_0[2471:2464]} - {1'b0, layer_0_0[2471:2464]};
      top_0[1] = {1'b0,layer_1_0[2479:2472]} - {1'b0, layer_0_0[2479:2472]};
      top_0[2] = {1'b0,layer_1_0[2487:2480]} - {1'b0, layer_0_0[2487:2480]};
      top_1[0] = {1'b0,layer_1_1[2471:2464]} - {1'b0, layer_0_1[2471:2464]};
      top_1[1] = {1'b0,layer_1_1[2479:2472]} - {1'b0, layer_0_1[2479:2472]};
      top_1[2] = {1'b0,layer_1_1[2487:2480]} - {1'b0, layer_0_1[2487:2480]};
      top_2[0] = {1'b0,layer_1_2[2471:2464]} - {1'b0, layer_0_2[2471:2464]};
      top_2[1] = {1'b0,layer_1_2[2479:2472]} - {1'b0, layer_0_2[2479:2472]};
      top_2[2] = {1'b0,layer_1_2[2487:2480]} - {1'b0, layer_0_2[2487:2480]};
      mid_0[0] = {1'b0,layer_2_0[2471:2464]} - {1'b0, layer_1_0[2471:2464]};
      mid_0[1] = {1'b0,layer_2_0[2479:2472]} - {1'b0, layer_1_0[2479:2472]};
      mid_0[2] = {1'b0,layer_2_0[2487:2480]} - {1'b0, layer_1_0[2487:2480]};
      mid_1[0] = {1'b0,layer_2_1[2471:2464]} - {1'b0, layer_1_1[2471:2464]};
      mid_1[1] = {1'b0,layer_2_1[2479:2472]} - {1'b0, layer_1_1[2479:2472]};
      mid_1[2] = {1'b0,layer_2_1[2487:2480]} - {1'b0, layer_1_1[2487:2480]};
      mid_2[0] = {1'b0,layer_2_2[2471:2464]} - {1'b0, layer_1_2[2471:2464]};
      mid_2[1] = {1'b0,layer_2_2[2479:2472]} - {1'b0, layer_1_2[2479:2472]};
      mid_2[2] = {1'b0,layer_2_2[2487:2480]} - {1'b0, layer_1_2[2487:2480]};
      btm_0[0] = {1'b0,layer_3_0[2471:2464]} - {1'b0, layer_2_0[2471:2464]};
      btm_0[1] = {1'b0,layer_3_0[2479:2472]} - {1'b0, layer_2_0[2479:2472]};
      btm_0[2] = {1'b0,layer_3_0[2487:2480]} - {1'b0, layer_2_0[2487:2480]};
      btm_1[0] = {1'b0,layer_3_1[2471:2464]} - {1'b0, layer_2_1[2471:2464]};
      btm_1[1] = {1'b0,layer_3_1[2479:2472]} - {1'b0, layer_2_1[2479:2472]};
      btm_1[2] = {1'b0,layer_3_1[2487:2480]} - {1'b0, layer_2_1[2487:2480]};
      btm_2[0] = {1'b0,layer_3_2[2471:2464]} - {1'b0, layer_2_2[2471:2464]};
      btm_2[1] = {1'b0,layer_3_2[2479:2472]} - {1'b0, layer_2_2[2479:2472]};
      btm_2[2] = {1'b0,layer_3_2[2487:2480]} - {1'b0, layer_2_2[2487:2480]};
    end
    'd310: begin
      top_0[0] = {1'b0,layer_1_0[2479:2472]} - {1'b0, layer_0_0[2479:2472]};
      top_0[1] = {1'b0,layer_1_0[2487:2480]} - {1'b0, layer_0_0[2487:2480]};
      top_0[2] = {1'b0,layer_1_0[2495:2488]} - {1'b0, layer_0_0[2495:2488]};
      top_1[0] = {1'b0,layer_1_1[2479:2472]} - {1'b0, layer_0_1[2479:2472]};
      top_1[1] = {1'b0,layer_1_1[2487:2480]} - {1'b0, layer_0_1[2487:2480]};
      top_1[2] = {1'b0,layer_1_1[2495:2488]} - {1'b0, layer_0_1[2495:2488]};
      top_2[0] = {1'b0,layer_1_2[2479:2472]} - {1'b0, layer_0_2[2479:2472]};
      top_2[1] = {1'b0,layer_1_2[2487:2480]} - {1'b0, layer_0_2[2487:2480]};
      top_2[2] = {1'b0,layer_1_2[2495:2488]} - {1'b0, layer_0_2[2495:2488]};
      mid_0[0] = {1'b0,layer_2_0[2479:2472]} - {1'b0, layer_1_0[2479:2472]};
      mid_0[1] = {1'b0,layer_2_0[2487:2480]} - {1'b0, layer_1_0[2487:2480]};
      mid_0[2] = {1'b0,layer_2_0[2495:2488]} - {1'b0, layer_1_0[2495:2488]};
      mid_1[0] = {1'b0,layer_2_1[2479:2472]} - {1'b0, layer_1_1[2479:2472]};
      mid_1[1] = {1'b0,layer_2_1[2487:2480]} - {1'b0, layer_1_1[2487:2480]};
      mid_1[2] = {1'b0,layer_2_1[2495:2488]} - {1'b0, layer_1_1[2495:2488]};
      mid_2[0] = {1'b0,layer_2_2[2479:2472]} - {1'b0, layer_1_2[2479:2472]};
      mid_2[1] = {1'b0,layer_2_2[2487:2480]} - {1'b0, layer_1_2[2487:2480]};
      mid_2[2] = {1'b0,layer_2_2[2495:2488]} - {1'b0, layer_1_2[2495:2488]};
      btm_0[0] = {1'b0,layer_3_0[2479:2472]} - {1'b0, layer_2_0[2479:2472]};
      btm_0[1] = {1'b0,layer_3_0[2487:2480]} - {1'b0, layer_2_0[2487:2480]};
      btm_0[2] = {1'b0,layer_3_0[2495:2488]} - {1'b0, layer_2_0[2495:2488]};
      btm_1[0] = {1'b0,layer_3_1[2479:2472]} - {1'b0, layer_2_1[2479:2472]};
      btm_1[1] = {1'b0,layer_3_1[2487:2480]} - {1'b0, layer_2_1[2487:2480]};
      btm_1[2] = {1'b0,layer_3_1[2495:2488]} - {1'b0, layer_2_1[2495:2488]};
      btm_2[0] = {1'b0,layer_3_2[2479:2472]} - {1'b0, layer_2_2[2479:2472]};
      btm_2[1] = {1'b0,layer_3_2[2487:2480]} - {1'b0, layer_2_2[2487:2480]};
      btm_2[2] = {1'b0,layer_3_2[2495:2488]} - {1'b0, layer_2_2[2495:2488]};
    end
    'd311: begin
      top_0[0] = {1'b0,layer_1_0[2487:2480]} - {1'b0, layer_0_0[2487:2480]};
      top_0[1] = {1'b0,layer_1_0[2495:2488]} - {1'b0, layer_0_0[2495:2488]};
      top_0[2] = {1'b0,layer_1_0[2503:2496]} - {1'b0, layer_0_0[2503:2496]};
      top_1[0] = {1'b0,layer_1_1[2487:2480]} - {1'b0, layer_0_1[2487:2480]};
      top_1[1] = {1'b0,layer_1_1[2495:2488]} - {1'b0, layer_0_1[2495:2488]};
      top_1[2] = {1'b0,layer_1_1[2503:2496]} - {1'b0, layer_0_1[2503:2496]};
      top_2[0] = {1'b0,layer_1_2[2487:2480]} - {1'b0, layer_0_2[2487:2480]};
      top_2[1] = {1'b0,layer_1_2[2495:2488]} - {1'b0, layer_0_2[2495:2488]};
      top_2[2] = {1'b0,layer_1_2[2503:2496]} - {1'b0, layer_0_2[2503:2496]};
      mid_0[0] = {1'b0,layer_2_0[2487:2480]} - {1'b0, layer_1_0[2487:2480]};
      mid_0[1] = {1'b0,layer_2_0[2495:2488]} - {1'b0, layer_1_0[2495:2488]};
      mid_0[2] = {1'b0,layer_2_0[2503:2496]} - {1'b0, layer_1_0[2503:2496]};
      mid_1[0] = {1'b0,layer_2_1[2487:2480]} - {1'b0, layer_1_1[2487:2480]};
      mid_1[1] = {1'b0,layer_2_1[2495:2488]} - {1'b0, layer_1_1[2495:2488]};
      mid_1[2] = {1'b0,layer_2_1[2503:2496]} - {1'b0, layer_1_1[2503:2496]};
      mid_2[0] = {1'b0,layer_2_2[2487:2480]} - {1'b0, layer_1_2[2487:2480]};
      mid_2[1] = {1'b0,layer_2_2[2495:2488]} - {1'b0, layer_1_2[2495:2488]};
      mid_2[2] = {1'b0,layer_2_2[2503:2496]} - {1'b0, layer_1_2[2503:2496]};
      btm_0[0] = {1'b0,layer_3_0[2487:2480]} - {1'b0, layer_2_0[2487:2480]};
      btm_0[1] = {1'b0,layer_3_0[2495:2488]} - {1'b0, layer_2_0[2495:2488]};
      btm_0[2] = {1'b0,layer_3_0[2503:2496]} - {1'b0, layer_2_0[2503:2496]};
      btm_1[0] = {1'b0,layer_3_1[2487:2480]} - {1'b0, layer_2_1[2487:2480]};
      btm_1[1] = {1'b0,layer_3_1[2495:2488]} - {1'b0, layer_2_1[2495:2488]};
      btm_1[2] = {1'b0,layer_3_1[2503:2496]} - {1'b0, layer_2_1[2503:2496]};
      btm_2[0] = {1'b0,layer_3_2[2487:2480]} - {1'b0, layer_2_2[2487:2480]};
      btm_2[1] = {1'b0,layer_3_2[2495:2488]} - {1'b0, layer_2_2[2495:2488]};
      btm_2[2] = {1'b0,layer_3_2[2503:2496]} - {1'b0, layer_2_2[2503:2496]};
    end
    'd312: begin
      top_0[0] = {1'b0,layer_1_0[2495:2488]} - {1'b0, layer_0_0[2495:2488]};
      top_0[1] = {1'b0,layer_1_0[2503:2496]} - {1'b0, layer_0_0[2503:2496]};
      top_0[2] = {1'b0,layer_1_0[2511:2504]} - {1'b0, layer_0_0[2511:2504]};
      top_1[0] = {1'b0,layer_1_1[2495:2488]} - {1'b0, layer_0_1[2495:2488]};
      top_1[1] = {1'b0,layer_1_1[2503:2496]} - {1'b0, layer_0_1[2503:2496]};
      top_1[2] = {1'b0,layer_1_1[2511:2504]} - {1'b0, layer_0_1[2511:2504]};
      top_2[0] = {1'b0,layer_1_2[2495:2488]} - {1'b0, layer_0_2[2495:2488]};
      top_2[1] = {1'b0,layer_1_2[2503:2496]} - {1'b0, layer_0_2[2503:2496]};
      top_2[2] = {1'b0,layer_1_2[2511:2504]} - {1'b0, layer_0_2[2511:2504]};
      mid_0[0] = {1'b0,layer_2_0[2495:2488]} - {1'b0, layer_1_0[2495:2488]};
      mid_0[1] = {1'b0,layer_2_0[2503:2496]} - {1'b0, layer_1_0[2503:2496]};
      mid_0[2] = {1'b0,layer_2_0[2511:2504]} - {1'b0, layer_1_0[2511:2504]};
      mid_1[0] = {1'b0,layer_2_1[2495:2488]} - {1'b0, layer_1_1[2495:2488]};
      mid_1[1] = {1'b0,layer_2_1[2503:2496]} - {1'b0, layer_1_1[2503:2496]};
      mid_1[2] = {1'b0,layer_2_1[2511:2504]} - {1'b0, layer_1_1[2511:2504]};
      mid_2[0] = {1'b0,layer_2_2[2495:2488]} - {1'b0, layer_1_2[2495:2488]};
      mid_2[1] = {1'b0,layer_2_2[2503:2496]} - {1'b0, layer_1_2[2503:2496]};
      mid_2[2] = {1'b0,layer_2_2[2511:2504]} - {1'b0, layer_1_2[2511:2504]};
      btm_0[0] = {1'b0,layer_3_0[2495:2488]} - {1'b0, layer_2_0[2495:2488]};
      btm_0[1] = {1'b0,layer_3_0[2503:2496]} - {1'b0, layer_2_0[2503:2496]};
      btm_0[2] = {1'b0,layer_3_0[2511:2504]} - {1'b0, layer_2_0[2511:2504]};
      btm_1[0] = {1'b0,layer_3_1[2495:2488]} - {1'b0, layer_2_1[2495:2488]};
      btm_1[1] = {1'b0,layer_3_1[2503:2496]} - {1'b0, layer_2_1[2503:2496]};
      btm_1[2] = {1'b0,layer_3_1[2511:2504]} - {1'b0, layer_2_1[2511:2504]};
      btm_2[0] = {1'b0,layer_3_2[2495:2488]} - {1'b0, layer_2_2[2495:2488]};
      btm_2[1] = {1'b0,layer_3_2[2503:2496]} - {1'b0, layer_2_2[2503:2496]};
      btm_2[2] = {1'b0,layer_3_2[2511:2504]} - {1'b0, layer_2_2[2511:2504]};
    end
    'd313: begin
      top_0[0] = {1'b0,layer_1_0[2503:2496]} - {1'b0, layer_0_0[2503:2496]};
      top_0[1] = {1'b0,layer_1_0[2511:2504]} - {1'b0, layer_0_0[2511:2504]};
      top_0[2] = {1'b0,layer_1_0[2519:2512]} - {1'b0, layer_0_0[2519:2512]};
      top_1[0] = {1'b0,layer_1_1[2503:2496]} - {1'b0, layer_0_1[2503:2496]};
      top_1[1] = {1'b0,layer_1_1[2511:2504]} - {1'b0, layer_0_1[2511:2504]};
      top_1[2] = {1'b0,layer_1_1[2519:2512]} - {1'b0, layer_0_1[2519:2512]};
      top_2[0] = {1'b0,layer_1_2[2503:2496]} - {1'b0, layer_0_2[2503:2496]};
      top_2[1] = {1'b0,layer_1_2[2511:2504]} - {1'b0, layer_0_2[2511:2504]};
      top_2[2] = {1'b0,layer_1_2[2519:2512]} - {1'b0, layer_0_2[2519:2512]};
      mid_0[0] = {1'b0,layer_2_0[2503:2496]} - {1'b0, layer_1_0[2503:2496]};
      mid_0[1] = {1'b0,layer_2_0[2511:2504]} - {1'b0, layer_1_0[2511:2504]};
      mid_0[2] = {1'b0,layer_2_0[2519:2512]} - {1'b0, layer_1_0[2519:2512]};
      mid_1[0] = {1'b0,layer_2_1[2503:2496]} - {1'b0, layer_1_1[2503:2496]};
      mid_1[1] = {1'b0,layer_2_1[2511:2504]} - {1'b0, layer_1_1[2511:2504]};
      mid_1[2] = {1'b0,layer_2_1[2519:2512]} - {1'b0, layer_1_1[2519:2512]};
      mid_2[0] = {1'b0,layer_2_2[2503:2496]} - {1'b0, layer_1_2[2503:2496]};
      mid_2[1] = {1'b0,layer_2_2[2511:2504]} - {1'b0, layer_1_2[2511:2504]};
      mid_2[2] = {1'b0,layer_2_2[2519:2512]} - {1'b0, layer_1_2[2519:2512]};
      btm_0[0] = {1'b0,layer_3_0[2503:2496]} - {1'b0, layer_2_0[2503:2496]};
      btm_0[1] = {1'b0,layer_3_0[2511:2504]} - {1'b0, layer_2_0[2511:2504]};
      btm_0[2] = {1'b0,layer_3_0[2519:2512]} - {1'b0, layer_2_0[2519:2512]};
      btm_1[0] = {1'b0,layer_3_1[2503:2496]} - {1'b0, layer_2_1[2503:2496]};
      btm_1[1] = {1'b0,layer_3_1[2511:2504]} - {1'b0, layer_2_1[2511:2504]};
      btm_1[2] = {1'b0,layer_3_1[2519:2512]} - {1'b0, layer_2_1[2519:2512]};
      btm_2[0] = {1'b0,layer_3_2[2503:2496]} - {1'b0, layer_2_2[2503:2496]};
      btm_2[1] = {1'b0,layer_3_2[2511:2504]} - {1'b0, layer_2_2[2511:2504]};
      btm_2[2] = {1'b0,layer_3_2[2519:2512]} - {1'b0, layer_2_2[2519:2512]};
    end
    'd314: begin
      top_0[0] = {1'b0,layer_1_0[2511:2504]} - {1'b0, layer_0_0[2511:2504]};
      top_0[1] = {1'b0,layer_1_0[2519:2512]} - {1'b0, layer_0_0[2519:2512]};
      top_0[2] = {1'b0,layer_1_0[2527:2520]} - {1'b0, layer_0_0[2527:2520]};
      top_1[0] = {1'b0,layer_1_1[2511:2504]} - {1'b0, layer_0_1[2511:2504]};
      top_1[1] = {1'b0,layer_1_1[2519:2512]} - {1'b0, layer_0_1[2519:2512]};
      top_1[2] = {1'b0,layer_1_1[2527:2520]} - {1'b0, layer_0_1[2527:2520]};
      top_2[0] = {1'b0,layer_1_2[2511:2504]} - {1'b0, layer_0_2[2511:2504]};
      top_2[1] = {1'b0,layer_1_2[2519:2512]} - {1'b0, layer_0_2[2519:2512]};
      top_2[2] = {1'b0,layer_1_2[2527:2520]} - {1'b0, layer_0_2[2527:2520]};
      mid_0[0] = {1'b0,layer_2_0[2511:2504]} - {1'b0, layer_1_0[2511:2504]};
      mid_0[1] = {1'b0,layer_2_0[2519:2512]} - {1'b0, layer_1_0[2519:2512]};
      mid_0[2] = {1'b0,layer_2_0[2527:2520]} - {1'b0, layer_1_0[2527:2520]};
      mid_1[0] = {1'b0,layer_2_1[2511:2504]} - {1'b0, layer_1_1[2511:2504]};
      mid_1[1] = {1'b0,layer_2_1[2519:2512]} - {1'b0, layer_1_1[2519:2512]};
      mid_1[2] = {1'b0,layer_2_1[2527:2520]} - {1'b0, layer_1_1[2527:2520]};
      mid_2[0] = {1'b0,layer_2_2[2511:2504]} - {1'b0, layer_1_2[2511:2504]};
      mid_2[1] = {1'b0,layer_2_2[2519:2512]} - {1'b0, layer_1_2[2519:2512]};
      mid_2[2] = {1'b0,layer_2_2[2527:2520]} - {1'b0, layer_1_2[2527:2520]};
      btm_0[0] = {1'b0,layer_3_0[2511:2504]} - {1'b0, layer_2_0[2511:2504]};
      btm_0[1] = {1'b0,layer_3_0[2519:2512]} - {1'b0, layer_2_0[2519:2512]};
      btm_0[2] = {1'b0,layer_3_0[2527:2520]} - {1'b0, layer_2_0[2527:2520]};
      btm_1[0] = {1'b0,layer_3_1[2511:2504]} - {1'b0, layer_2_1[2511:2504]};
      btm_1[1] = {1'b0,layer_3_1[2519:2512]} - {1'b0, layer_2_1[2519:2512]};
      btm_1[2] = {1'b0,layer_3_1[2527:2520]} - {1'b0, layer_2_1[2527:2520]};
      btm_2[0] = {1'b0,layer_3_2[2511:2504]} - {1'b0, layer_2_2[2511:2504]};
      btm_2[1] = {1'b0,layer_3_2[2519:2512]} - {1'b0, layer_2_2[2519:2512]};
      btm_2[2] = {1'b0,layer_3_2[2527:2520]} - {1'b0, layer_2_2[2527:2520]};
    end
    'd315: begin
      top_0[0] = {1'b0,layer_1_0[2519:2512]} - {1'b0, layer_0_0[2519:2512]};
      top_0[1] = {1'b0,layer_1_0[2527:2520]} - {1'b0, layer_0_0[2527:2520]};
      top_0[2] = {1'b0,layer_1_0[2535:2528]} - {1'b0, layer_0_0[2535:2528]};
      top_1[0] = {1'b0,layer_1_1[2519:2512]} - {1'b0, layer_0_1[2519:2512]};
      top_1[1] = {1'b0,layer_1_1[2527:2520]} - {1'b0, layer_0_1[2527:2520]};
      top_1[2] = {1'b0,layer_1_1[2535:2528]} - {1'b0, layer_0_1[2535:2528]};
      top_2[0] = {1'b0,layer_1_2[2519:2512]} - {1'b0, layer_0_2[2519:2512]};
      top_2[1] = {1'b0,layer_1_2[2527:2520]} - {1'b0, layer_0_2[2527:2520]};
      top_2[2] = {1'b0,layer_1_2[2535:2528]} - {1'b0, layer_0_2[2535:2528]};
      mid_0[0] = {1'b0,layer_2_0[2519:2512]} - {1'b0, layer_1_0[2519:2512]};
      mid_0[1] = {1'b0,layer_2_0[2527:2520]} - {1'b0, layer_1_0[2527:2520]};
      mid_0[2] = {1'b0,layer_2_0[2535:2528]} - {1'b0, layer_1_0[2535:2528]};
      mid_1[0] = {1'b0,layer_2_1[2519:2512]} - {1'b0, layer_1_1[2519:2512]};
      mid_1[1] = {1'b0,layer_2_1[2527:2520]} - {1'b0, layer_1_1[2527:2520]};
      mid_1[2] = {1'b0,layer_2_1[2535:2528]} - {1'b0, layer_1_1[2535:2528]};
      mid_2[0] = {1'b0,layer_2_2[2519:2512]} - {1'b0, layer_1_2[2519:2512]};
      mid_2[1] = {1'b0,layer_2_2[2527:2520]} - {1'b0, layer_1_2[2527:2520]};
      mid_2[2] = {1'b0,layer_2_2[2535:2528]} - {1'b0, layer_1_2[2535:2528]};
      btm_0[0] = {1'b0,layer_3_0[2519:2512]} - {1'b0, layer_2_0[2519:2512]};
      btm_0[1] = {1'b0,layer_3_0[2527:2520]} - {1'b0, layer_2_0[2527:2520]};
      btm_0[2] = {1'b0,layer_3_0[2535:2528]} - {1'b0, layer_2_0[2535:2528]};
      btm_1[0] = {1'b0,layer_3_1[2519:2512]} - {1'b0, layer_2_1[2519:2512]};
      btm_1[1] = {1'b0,layer_3_1[2527:2520]} - {1'b0, layer_2_1[2527:2520]};
      btm_1[2] = {1'b0,layer_3_1[2535:2528]} - {1'b0, layer_2_1[2535:2528]};
      btm_2[0] = {1'b0,layer_3_2[2519:2512]} - {1'b0, layer_2_2[2519:2512]};
      btm_2[1] = {1'b0,layer_3_2[2527:2520]} - {1'b0, layer_2_2[2527:2520]};
      btm_2[2] = {1'b0,layer_3_2[2535:2528]} - {1'b0, layer_2_2[2535:2528]};
    end
    'd316: begin
      top_0[0] = {1'b0,layer_1_0[2527:2520]} - {1'b0, layer_0_0[2527:2520]};
      top_0[1] = {1'b0,layer_1_0[2535:2528]} - {1'b0, layer_0_0[2535:2528]};
      top_0[2] = {1'b0,layer_1_0[2543:2536]} - {1'b0, layer_0_0[2543:2536]};
      top_1[0] = {1'b0,layer_1_1[2527:2520]} - {1'b0, layer_0_1[2527:2520]};
      top_1[1] = {1'b0,layer_1_1[2535:2528]} - {1'b0, layer_0_1[2535:2528]};
      top_1[2] = {1'b0,layer_1_1[2543:2536]} - {1'b0, layer_0_1[2543:2536]};
      top_2[0] = {1'b0,layer_1_2[2527:2520]} - {1'b0, layer_0_2[2527:2520]};
      top_2[1] = {1'b0,layer_1_2[2535:2528]} - {1'b0, layer_0_2[2535:2528]};
      top_2[2] = {1'b0,layer_1_2[2543:2536]} - {1'b0, layer_0_2[2543:2536]};
      mid_0[0] = {1'b0,layer_2_0[2527:2520]} - {1'b0, layer_1_0[2527:2520]};
      mid_0[1] = {1'b0,layer_2_0[2535:2528]} - {1'b0, layer_1_0[2535:2528]};
      mid_0[2] = {1'b0,layer_2_0[2543:2536]} - {1'b0, layer_1_0[2543:2536]};
      mid_1[0] = {1'b0,layer_2_1[2527:2520]} - {1'b0, layer_1_1[2527:2520]};
      mid_1[1] = {1'b0,layer_2_1[2535:2528]} - {1'b0, layer_1_1[2535:2528]};
      mid_1[2] = {1'b0,layer_2_1[2543:2536]} - {1'b0, layer_1_1[2543:2536]};
      mid_2[0] = {1'b0,layer_2_2[2527:2520]} - {1'b0, layer_1_2[2527:2520]};
      mid_2[1] = {1'b0,layer_2_2[2535:2528]} - {1'b0, layer_1_2[2535:2528]};
      mid_2[2] = {1'b0,layer_2_2[2543:2536]} - {1'b0, layer_1_2[2543:2536]};
      btm_0[0] = {1'b0,layer_3_0[2527:2520]} - {1'b0, layer_2_0[2527:2520]};
      btm_0[1] = {1'b0,layer_3_0[2535:2528]} - {1'b0, layer_2_0[2535:2528]};
      btm_0[2] = {1'b0,layer_3_0[2543:2536]} - {1'b0, layer_2_0[2543:2536]};
      btm_1[0] = {1'b0,layer_3_1[2527:2520]} - {1'b0, layer_2_1[2527:2520]};
      btm_1[1] = {1'b0,layer_3_1[2535:2528]} - {1'b0, layer_2_1[2535:2528]};
      btm_1[2] = {1'b0,layer_3_1[2543:2536]} - {1'b0, layer_2_1[2543:2536]};
      btm_2[0] = {1'b0,layer_3_2[2527:2520]} - {1'b0, layer_2_2[2527:2520]};
      btm_2[1] = {1'b0,layer_3_2[2535:2528]} - {1'b0, layer_2_2[2535:2528]};
      btm_2[2] = {1'b0,layer_3_2[2543:2536]} - {1'b0, layer_2_2[2543:2536]};
    end
    'd317: begin
      top_0[0] = {1'b0,layer_1_0[2535:2528]} - {1'b0, layer_0_0[2535:2528]};
      top_0[1] = {1'b0,layer_1_0[2543:2536]} - {1'b0, layer_0_0[2543:2536]};
      top_0[2] = {1'b0,layer_1_0[2551:2544]} - {1'b0, layer_0_0[2551:2544]};
      top_1[0] = {1'b0,layer_1_1[2535:2528]} - {1'b0, layer_0_1[2535:2528]};
      top_1[1] = {1'b0,layer_1_1[2543:2536]} - {1'b0, layer_0_1[2543:2536]};
      top_1[2] = {1'b0,layer_1_1[2551:2544]} - {1'b0, layer_0_1[2551:2544]};
      top_2[0] = {1'b0,layer_1_2[2535:2528]} - {1'b0, layer_0_2[2535:2528]};
      top_2[1] = {1'b0,layer_1_2[2543:2536]} - {1'b0, layer_0_2[2543:2536]};
      top_2[2] = {1'b0,layer_1_2[2551:2544]} - {1'b0, layer_0_2[2551:2544]};
      mid_0[0] = {1'b0,layer_2_0[2535:2528]} - {1'b0, layer_1_0[2535:2528]};
      mid_0[1] = {1'b0,layer_2_0[2543:2536]} - {1'b0, layer_1_0[2543:2536]};
      mid_0[2] = {1'b0,layer_2_0[2551:2544]} - {1'b0, layer_1_0[2551:2544]};
      mid_1[0] = {1'b0,layer_2_1[2535:2528]} - {1'b0, layer_1_1[2535:2528]};
      mid_1[1] = {1'b0,layer_2_1[2543:2536]} - {1'b0, layer_1_1[2543:2536]};
      mid_1[2] = {1'b0,layer_2_1[2551:2544]} - {1'b0, layer_1_1[2551:2544]};
      mid_2[0] = {1'b0,layer_2_2[2535:2528]} - {1'b0, layer_1_2[2535:2528]};
      mid_2[1] = {1'b0,layer_2_2[2543:2536]} - {1'b0, layer_1_2[2543:2536]};
      mid_2[2] = {1'b0,layer_2_2[2551:2544]} - {1'b0, layer_1_2[2551:2544]};
      btm_0[0] = {1'b0,layer_3_0[2535:2528]} - {1'b0, layer_2_0[2535:2528]};
      btm_0[1] = {1'b0,layer_3_0[2543:2536]} - {1'b0, layer_2_0[2543:2536]};
      btm_0[2] = {1'b0,layer_3_0[2551:2544]} - {1'b0, layer_2_0[2551:2544]};
      btm_1[0] = {1'b0,layer_3_1[2535:2528]} - {1'b0, layer_2_1[2535:2528]};
      btm_1[1] = {1'b0,layer_3_1[2543:2536]} - {1'b0, layer_2_1[2543:2536]};
      btm_1[2] = {1'b0,layer_3_1[2551:2544]} - {1'b0, layer_2_1[2551:2544]};
      btm_2[0] = {1'b0,layer_3_2[2535:2528]} - {1'b0, layer_2_2[2535:2528]};
      btm_2[1] = {1'b0,layer_3_2[2543:2536]} - {1'b0, layer_2_2[2543:2536]};
      btm_2[2] = {1'b0,layer_3_2[2551:2544]} - {1'b0, layer_2_2[2551:2544]};
    end
    'd318: begin
      top_0[0] = {1'b0,layer_1_0[2543:2536]} - {1'b0, layer_0_0[2543:2536]};
      top_0[1] = {1'b0,layer_1_0[2551:2544]} - {1'b0, layer_0_0[2551:2544]};
      top_0[2] = {1'b0,layer_1_0[2559:2552]} - {1'b0, layer_0_0[2559:2552]};
      top_1[0] = {1'b0,layer_1_1[2543:2536]} - {1'b0, layer_0_1[2543:2536]};
      top_1[1] = {1'b0,layer_1_1[2551:2544]} - {1'b0, layer_0_1[2551:2544]};
      top_1[2] = {1'b0,layer_1_1[2559:2552]} - {1'b0, layer_0_1[2559:2552]};
      top_2[0] = {1'b0,layer_1_2[2543:2536]} - {1'b0, layer_0_2[2543:2536]};
      top_2[1] = {1'b0,layer_1_2[2551:2544]} - {1'b0, layer_0_2[2551:2544]};
      top_2[2] = {1'b0,layer_1_2[2559:2552]} - {1'b0, layer_0_2[2559:2552]};
      mid_0[0] = {1'b0,layer_2_0[2543:2536]} - {1'b0, layer_1_0[2543:2536]};
      mid_0[1] = {1'b0,layer_2_0[2551:2544]} - {1'b0, layer_1_0[2551:2544]};
      mid_0[2] = {1'b0,layer_2_0[2559:2552]} - {1'b0, layer_1_0[2559:2552]};
      mid_1[0] = {1'b0,layer_2_1[2543:2536]} - {1'b0, layer_1_1[2543:2536]};
      mid_1[1] = {1'b0,layer_2_1[2551:2544]} - {1'b0, layer_1_1[2551:2544]};
      mid_1[2] = {1'b0,layer_2_1[2559:2552]} - {1'b0, layer_1_1[2559:2552]};
      mid_2[0] = {1'b0,layer_2_2[2543:2536]} - {1'b0, layer_1_2[2543:2536]};
      mid_2[1] = {1'b0,layer_2_2[2551:2544]} - {1'b0, layer_1_2[2551:2544]};
      mid_2[2] = {1'b0,layer_2_2[2559:2552]} - {1'b0, layer_1_2[2559:2552]};
      btm_0[0] = {1'b0,layer_3_0[2543:2536]} - {1'b0, layer_2_0[2543:2536]};
      btm_0[1] = {1'b0,layer_3_0[2551:2544]} - {1'b0, layer_2_0[2551:2544]};
      btm_0[2] = {1'b0,layer_3_0[2559:2552]} - {1'b0, layer_2_0[2559:2552]};
      btm_1[0] = {1'b0,layer_3_1[2543:2536]} - {1'b0, layer_2_1[2543:2536]};
      btm_1[1] = {1'b0,layer_3_1[2551:2544]} - {1'b0, layer_2_1[2551:2544]};
      btm_1[2] = {1'b0,layer_3_1[2559:2552]} - {1'b0, layer_2_1[2559:2552]};
      btm_2[0] = {1'b0,layer_3_2[2543:2536]} - {1'b0, layer_2_2[2543:2536]};
      btm_2[1] = {1'b0,layer_3_2[2551:2544]} - {1'b0, layer_2_2[2551:2544]};
      btm_2[2] = {1'b0,layer_3_2[2559:2552]} - {1'b0, layer_2_2[2559:2552]};
    end
    'd319: begin
      top_0[0] = {1'b0,layer_1_0[2551:2544]} - {1'b0, layer_0_0[2551:2544]};
      top_0[1] = {1'b0,layer_1_0[2559:2552]} - {1'b0, layer_0_0[2559:2552]};
      top_0[2] = {1'b0,layer_1_0[2567:2560]} - {1'b0, layer_0_0[2567:2560]};
      top_1[0] = {1'b0,layer_1_1[2551:2544]} - {1'b0, layer_0_1[2551:2544]};
      top_1[1] = {1'b0,layer_1_1[2559:2552]} - {1'b0, layer_0_1[2559:2552]};
      top_1[2] = {1'b0,layer_1_1[2567:2560]} - {1'b0, layer_0_1[2567:2560]};
      top_2[0] = {1'b0,layer_1_2[2551:2544]} - {1'b0, layer_0_2[2551:2544]};
      top_2[1] = {1'b0,layer_1_2[2559:2552]} - {1'b0, layer_0_2[2559:2552]};
      top_2[2] = {1'b0,layer_1_2[2567:2560]} - {1'b0, layer_0_2[2567:2560]};
      mid_0[0] = {1'b0,layer_2_0[2551:2544]} - {1'b0, layer_1_0[2551:2544]};
      mid_0[1] = {1'b0,layer_2_0[2559:2552]} - {1'b0, layer_1_0[2559:2552]};
      mid_0[2] = {1'b0,layer_2_0[2567:2560]} - {1'b0, layer_1_0[2567:2560]};
      mid_1[0] = {1'b0,layer_2_1[2551:2544]} - {1'b0, layer_1_1[2551:2544]};
      mid_1[1] = {1'b0,layer_2_1[2559:2552]} - {1'b0, layer_1_1[2559:2552]};
      mid_1[2] = {1'b0,layer_2_1[2567:2560]} - {1'b0, layer_1_1[2567:2560]};
      mid_2[0] = {1'b0,layer_2_2[2551:2544]} - {1'b0, layer_1_2[2551:2544]};
      mid_2[1] = {1'b0,layer_2_2[2559:2552]} - {1'b0, layer_1_2[2559:2552]};
      mid_2[2] = {1'b0,layer_2_2[2567:2560]} - {1'b0, layer_1_2[2567:2560]};
      btm_0[0] = {1'b0,layer_3_0[2551:2544]} - {1'b0, layer_2_0[2551:2544]};
      btm_0[1] = {1'b0,layer_3_0[2559:2552]} - {1'b0, layer_2_0[2559:2552]};
      btm_0[2] = {1'b0,layer_3_0[2567:2560]} - {1'b0, layer_2_0[2567:2560]};
      btm_1[0] = {1'b0,layer_3_1[2551:2544]} - {1'b0, layer_2_1[2551:2544]};
      btm_1[1] = {1'b0,layer_3_1[2559:2552]} - {1'b0, layer_2_1[2559:2552]};
      btm_1[2] = {1'b0,layer_3_1[2567:2560]} - {1'b0, layer_2_1[2567:2560]};
      btm_2[0] = {1'b0,layer_3_2[2551:2544]} - {1'b0, layer_2_2[2551:2544]};
      btm_2[1] = {1'b0,layer_3_2[2559:2552]} - {1'b0, layer_2_2[2559:2552]};
      btm_2[2] = {1'b0,layer_3_2[2567:2560]} - {1'b0, layer_2_2[2567:2560]};
    end
    'd320: begin
      top_0[0] = {1'b0,layer_1_0[2559:2552]} - {1'b0, layer_0_0[2559:2552]};
      top_0[1] = {1'b0,layer_1_0[2567:2560]} - {1'b0, layer_0_0[2567:2560]};
      top_0[2] = {1'b0,layer_1_0[2575:2568]} - {1'b0, layer_0_0[2575:2568]};
      top_1[0] = {1'b0,layer_1_1[2559:2552]} - {1'b0, layer_0_1[2559:2552]};
      top_1[1] = {1'b0,layer_1_1[2567:2560]} - {1'b0, layer_0_1[2567:2560]};
      top_1[2] = {1'b0,layer_1_1[2575:2568]} - {1'b0, layer_0_1[2575:2568]};
      top_2[0] = {1'b0,layer_1_2[2559:2552]} - {1'b0, layer_0_2[2559:2552]};
      top_2[1] = {1'b0,layer_1_2[2567:2560]} - {1'b0, layer_0_2[2567:2560]};
      top_2[2] = {1'b0,layer_1_2[2575:2568]} - {1'b0, layer_0_2[2575:2568]};
      mid_0[0] = {1'b0,layer_2_0[2559:2552]} - {1'b0, layer_1_0[2559:2552]};
      mid_0[1] = {1'b0,layer_2_0[2567:2560]} - {1'b0, layer_1_0[2567:2560]};
      mid_0[2] = {1'b0,layer_2_0[2575:2568]} - {1'b0, layer_1_0[2575:2568]};
      mid_1[0] = {1'b0,layer_2_1[2559:2552]} - {1'b0, layer_1_1[2559:2552]};
      mid_1[1] = {1'b0,layer_2_1[2567:2560]} - {1'b0, layer_1_1[2567:2560]};
      mid_1[2] = {1'b0,layer_2_1[2575:2568]} - {1'b0, layer_1_1[2575:2568]};
      mid_2[0] = {1'b0,layer_2_2[2559:2552]} - {1'b0, layer_1_2[2559:2552]};
      mid_2[1] = {1'b0,layer_2_2[2567:2560]} - {1'b0, layer_1_2[2567:2560]};
      mid_2[2] = {1'b0,layer_2_2[2575:2568]} - {1'b0, layer_1_2[2575:2568]};
      btm_0[0] = {1'b0,layer_3_0[2559:2552]} - {1'b0, layer_2_0[2559:2552]};
      btm_0[1] = {1'b0,layer_3_0[2567:2560]} - {1'b0, layer_2_0[2567:2560]};
      btm_0[2] = {1'b0,layer_3_0[2575:2568]} - {1'b0, layer_2_0[2575:2568]};
      btm_1[0] = {1'b0,layer_3_1[2559:2552]} - {1'b0, layer_2_1[2559:2552]};
      btm_1[1] = {1'b0,layer_3_1[2567:2560]} - {1'b0, layer_2_1[2567:2560]};
      btm_1[2] = {1'b0,layer_3_1[2575:2568]} - {1'b0, layer_2_1[2575:2568]};
      btm_2[0] = {1'b0,layer_3_2[2559:2552]} - {1'b0, layer_2_2[2559:2552]};
      btm_2[1] = {1'b0,layer_3_2[2567:2560]} - {1'b0, layer_2_2[2567:2560]};
      btm_2[2] = {1'b0,layer_3_2[2575:2568]} - {1'b0, layer_2_2[2575:2568]};
    end
    'd321: begin
      top_0[0] = {1'b0,layer_1_0[2567:2560]} - {1'b0, layer_0_0[2567:2560]};
      top_0[1] = {1'b0,layer_1_0[2575:2568]} - {1'b0, layer_0_0[2575:2568]};
      top_0[2] = {1'b0,layer_1_0[2583:2576]} - {1'b0, layer_0_0[2583:2576]};
      top_1[0] = {1'b0,layer_1_1[2567:2560]} - {1'b0, layer_0_1[2567:2560]};
      top_1[1] = {1'b0,layer_1_1[2575:2568]} - {1'b0, layer_0_1[2575:2568]};
      top_1[2] = {1'b0,layer_1_1[2583:2576]} - {1'b0, layer_0_1[2583:2576]};
      top_2[0] = {1'b0,layer_1_2[2567:2560]} - {1'b0, layer_0_2[2567:2560]};
      top_2[1] = {1'b0,layer_1_2[2575:2568]} - {1'b0, layer_0_2[2575:2568]};
      top_2[2] = {1'b0,layer_1_2[2583:2576]} - {1'b0, layer_0_2[2583:2576]};
      mid_0[0] = {1'b0,layer_2_0[2567:2560]} - {1'b0, layer_1_0[2567:2560]};
      mid_0[1] = {1'b0,layer_2_0[2575:2568]} - {1'b0, layer_1_0[2575:2568]};
      mid_0[2] = {1'b0,layer_2_0[2583:2576]} - {1'b0, layer_1_0[2583:2576]};
      mid_1[0] = {1'b0,layer_2_1[2567:2560]} - {1'b0, layer_1_1[2567:2560]};
      mid_1[1] = {1'b0,layer_2_1[2575:2568]} - {1'b0, layer_1_1[2575:2568]};
      mid_1[2] = {1'b0,layer_2_1[2583:2576]} - {1'b0, layer_1_1[2583:2576]};
      mid_2[0] = {1'b0,layer_2_2[2567:2560]} - {1'b0, layer_1_2[2567:2560]};
      mid_2[1] = {1'b0,layer_2_2[2575:2568]} - {1'b0, layer_1_2[2575:2568]};
      mid_2[2] = {1'b0,layer_2_2[2583:2576]} - {1'b0, layer_1_2[2583:2576]};
      btm_0[0] = {1'b0,layer_3_0[2567:2560]} - {1'b0, layer_2_0[2567:2560]};
      btm_0[1] = {1'b0,layer_3_0[2575:2568]} - {1'b0, layer_2_0[2575:2568]};
      btm_0[2] = {1'b0,layer_3_0[2583:2576]} - {1'b0, layer_2_0[2583:2576]};
      btm_1[0] = {1'b0,layer_3_1[2567:2560]} - {1'b0, layer_2_1[2567:2560]};
      btm_1[1] = {1'b0,layer_3_1[2575:2568]} - {1'b0, layer_2_1[2575:2568]};
      btm_1[2] = {1'b0,layer_3_1[2583:2576]} - {1'b0, layer_2_1[2583:2576]};
      btm_2[0] = {1'b0,layer_3_2[2567:2560]} - {1'b0, layer_2_2[2567:2560]};
      btm_2[1] = {1'b0,layer_3_2[2575:2568]} - {1'b0, layer_2_2[2575:2568]};
      btm_2[2] = {1'b0,layer_3_2[2583:2576]} - {1'b0, layer_2_2[2583:2576]};
    end
    'd322: begin
      top_0[0] = {1'b0,layer_1_0[2575:2568]} - {1'b0, layer_0_0[2575:2568]};
      top_0[1] = {1'b0,layer_1_0[2583:2576]} - {1'b0, layer_0_0[2583:2576]};
      top_0[2] = {1'b0,layer_1_0[2591:2584]} - {1'b0, layer_0_0[2591:2584]};
      top_1[0] = {1'b0,layer_1_1[2575:2568]} - {1'b0, layer_0_1[2575:2568]};
      top_1[1] = {1'b0,layer_1_1[2583:2576]} - {1'b0, layer_0_1[2583:2576]};
      top_1[2] = {1'b0,layer_1_1[2591:2584]} - {1'b0, layer_0_1[2591:2584]};
      top_2[0] = {1'b0,layer_1_2[2575:2568]} - {1'b0, layer_0_2[2575:2568]};
      top_2[1] = {1'b0,layer_1_2[2583:2576]} - {1'b0, layer_0_2[2583:2576]};
      top_2[2] = {1'b0,layer_1_2[2591:2584]} - {1'b0, layer_0_2[2591:2584]};
      mid_0[0] = {1'b0,layer_2_0[2575:2568]} - {1'b0, layer_1_0[2575:2568]};
      mid_0[1] = {1'b0,layer_2_0[2583:2576]} - {1'b0, layer_1_0[2583:2576]};
      mid_0[2] = {1'b0,layer_2_0[2591:2584]} - {1'b0, layer_1_0[2591:2584]};
      mid_1[0] = {1'b0,layer_2_1[2575:2568]} - {1'b0, layer_1_1[2575:2568]};
      mid_1[1] = {1'b0,layer_2_1[2583:2576]} - {1'b0, layer_1_1[2583:2576]};
      mid_1[2] = {1'b0,layer_2_1[2591:2584]} - {1'b0, layer_1_1[2591:2584]};
      mid_2[0] = {1'b0,layer_2_2[2575:2568]} - {1'b0, layer_1_2[2575:2568]};
      mid_2[1] = {1'b0,layer_2_2[2583:2576]} - {1'b0, layer_1_2[2583:2576]};
      mid_2[2] = {1'b0,layer_2_2[2591:2584]} - {1'b0, layer_1_2[2591:2584]};
      btm_0[0] = {1'b0,layer_3_0[2575:2568]} - {1'b0, layer_2_0[2575:2568]};
      btm_0[1] = {1'b0,layer_3_0[2583:2576]} - {1'b0, layer_2_0[2583:2576]};
      btm_0[2] = {1'b0,layer_3_0[2591:2584]} - {1'b0, layer_2_0[2591:2584]};
      btm_1[0] = {1'b0,layer_3_1[2575:2568]} - {1'b0, layer_2_1[2575:2568]};
      btm_1[1] = {1'b0,layer_3_1[2583:2576]} - {1'b0, layer_2_1[2583:2576]};
      btm_1[2] = {1'b0,layer_3_1[2591:2584]} - {1'b0, layer_2_1[2591:2584]};
      btm_2[0] = {1'b0,layer_3_2[2575:2568]} - {1'b0, layer_2_2[2575:2568]};
      btm_2[1] = {1'b0,layer_3_2[2583:2576]} - {1'b0, layer_2_2[2583:2576]};
      btm_2[2] = {1'b0,layer_3_2[2591:2584]} - {1'b0, layer_2_2[2591:2584]};
    end
    'd323: begin
      top_0[0] = {1'b0,layer_1_0[2583:2576]} - {1'b0, layer_0_0[2583:2576]};
      top_0[1] = {1'b0,layer_1_0[2591:2584]} - {1'b0, layer_0_0[2591:2584]};
      top_0[2] = {1'b0,layer_1_0[2599:2592]} - {1'b0, layer_0_0[2599:2592]};
      top_1[0] = {1'b0,layer_1_1[2583:2576]} - {1'b0, layer_0_1[2583:2576]};
      top_1[1] = {1'b0,layer_1_1[2591:2584]} - {1'b0, layer_0_1[2591:2584]};
      top_1[2] = {1'b0,layer_1_1[2599:2592]} - {1'b0, layer_0_1[2599:2592]};
      top_2[0] = {1'b0,layer_1_2[2583:2576]} - {1'b0, layer_0_2[2583:2576]};
      top_2[1] = {1'b0,layer_1_2[2591:2584]} - {1'b0, layer_0_2[2591:2584]};
      top_2[2] = {1'b0,layer_1_2[2599:2592]} - {1'b0, layer_0_2[2599:2592]};
      mid_0[0] = {1'b0,layer_2_0[2583:2576]} - {1'b0, layer_1_0[2583:2576]};
      mid_0[1] = {1'b0,layer_2_0[2591:2584]} - {1'b0, layer_1_0[2591:2584]};
      mid_0[2] = {1'b0,layer_2_0[2599:2592]} - {1'b0, layer_1_0[2599:2592]};
      mid_1[0] = {1'b0,layer_2_1[2583:2576]} - {1'b0, layer_1_1[2583:2576]};
      mid_1[1] = {1'b0,layer_2_1[2591:2584]} - {1'b0, layer_1_1[2591:2584]};
      mid_1[2] = {1'b0,layer_2_1[2599:2592]} - {1'b0, layer_1_1[2599:2592]};
      mid_2[0] = {1'b0,layer_2_2[2583:2576]} - {1'b0, layer_1_2[2583:2576]};
      mid_2[1] = {1'b0,layer_2_2[2591:2584]} - {1'b0, layer_1_2[2591:2584]};
      mid_2[2] = {1'b0,layer_2_2[2599:2592]} - {1'b0, layer_1_2[2599:2592]};
      btm_0[0] = {1'b0,layer_3_0[2583:2576]} - {1'b0, layer_2_0[2583:2576]};
      btm_0[1] = {1'b0,layer_3_0[2591:2584]} - {1'b0, layer_2_0[2591:2584]};
      btm_0[2] = {1'b0,layer_3_0[2599:2592]} - {1'b0, layer_2_0[2599:2592]};
      btm_1[0] = {1'b0,layer_3_1[2583:2576]} - {1'b0, layer_2_1[2583:2576]};
      btm_1[1] = {1'b0,layer_3_1[2591:2584]} - {1'b0, layer_2_1[2591:2584]};
      btm_1[2] = {1'b0,layer_3_1[2599:2592]} - {1'b0, layer_2_1[2599:2592]};
      btm_2[0] = {1'b0,layer_3_2[2583:2576]} - {1'b0, layer_2_2[2583:2576]};
      btm_2[1] = {1'b0,layer_3_2[2591:2584]} - {1'b0, layer_2_2[2591:2584]};
      btm_2[2] = {1'b0,layer_3_2[2599:2592]} - {1'b0, layer_2_2[2599:2592]};
    end
    'd324: begin
      top_0[0] = {1'b0,layer_1_0[2591:2584]} - {1'b0, layer_0_0[2591:2584]};
      top_0[1] = {1'b0,layer_1_0[2599:2592]} - {1'b0, layer_0_0[2599:2592]};
      top_0[2] = {1'b0,layer_1_0[2607:2600]} - {1'b0, layer_0_0[2607:2600]};
      top_1[0] = {1'b0,layer_1_1[2591:2584]} - {1'b0, layer_0_1[2591:2584]};
      top_1[1] = {1'b0,layer_1_1[2599:2592]} - {1'b0, layer_0_1[2599:2592]};
      top_1[2] = {1'b0,layer_1_1[2607:2600]} - {1'b0, layer_0_1[2607:2600]};
      top_2[0] = {1'b0,layer_1_2[2591:2584]} - {1'b0, layer_0_2[2591:2584]};
      top_2[1] = {1'b0,layer_1_2[2599:2592]} - {1'b0, layer_0_2[2599:2592]};
      top_2[2] = {1'b0,layer_1_2[2607:2600]} - {1'b0, layer_0_2[2607:2600]};
      mid_0[0] = {1'b0,layer_2_0[2591:2584]} - {1'b0, layer_1_0[2591:2584]};
      mid_0[1] = {1'b0,layer_2_0[2599:2592]} - {1'b0, layer_1_0[2599:2592]};
      mid_0[2] = {1'b0,layer_2_0[2607:2600]} - {1'b0, layer_1_0[2607:2600]};
      mid_1[0] = {1'b0,layer_2_1[2591:2584]} - {1'b0, layer_1_1[2591:2584]};
      mid_1[1] = {1'b0,layer_2_1[2599:2592]} - {1'b0, layer_1_1[2599:2592]};
      mid_1[2] = {1'b0,layer_2_1[2607:2600]} - {1'b0, layer_1_1[2607:2600]};
      mid_2[0] = {1'b0,layer_2_2[2591:2584]} - {1'b0, layer_1_2[2591:2584]};
      mid_2[1] = {1'b0,layer_2_2[2599:2592]} - {1'b0, layer_1_2[2599:2592]};
      mid_2[2] = {1'b0,layer_2_2[2607:2600]} - {1'b0, layer_1_2[2607:2600]};
      btm_0[0] = {1'b0,layer_3_0[2591:2584]} - {1'b0, layer_2_0[2591:2584]};
      btm_0[1] = {1'b0,layer_3_0[2599:2592]} - {1'b0, layer_2_0[2599:2592]};
      btm_0[2] = {1'b0,layer_3_0[2607:2600]} - {1'b0, layer_2_0[2607:2600]};
      btm_1[0] = {1'b0,layer_3_1[2591:2584]} - {1'b0, layer_2_1[2591:2584]};
      btm_1[1] = {1'b0,layer_3_1[2599:2592]} - {1'b0, layer_2_1[2599:2592]};
      btm_1[2] = {1'b0,layer_3_1[2607:2600]} - {1'b0, layer_2_1[2607:2600]};
      btm_2[0] = {1'b0,layer_3_2[2591:2584]} - {1'b0, layer_2_2[2591:2584]};
      btm_2[1] = {1'b0,layer_3_2[2599:2592]} - {1'b0, layer_2_2[2599:2592]};
      btm_2[2] = {1'b0,layer_3_2[2607:2600]} - {1'b0, layer_2_2[2607:2600]};
    end
    'd325: begin
      top_0[0] = {1'b0,layer_1_0[2599:2592]} - {1'b0, layer_0_0[2599:2592]};
      top_0[1] = {1'b0,layer_1_0[2607:2600]} - {1'b0, layer_0_0[2607:2600]};
      top_0[2] = {1'b0,layer_1_0[2615:2608]} - {1'b0, layer_0_0[2615:2608]};
      top_1[0] = {1'b0,layer_1_1[2599:2592]} - {1'b0, layer_0_1[2599:2592]};
      top_1[1] = {1'b0,layer_1_1[2607:2600]} - {1'b0, layer_0_1[2607:2600]};
      top_1[2] = {1'b0,layer_1_1[2615:2608]} - {1'b0, layer_0_1[2615:2608]};
      top_2[0] = {1'b0,layer_1_2[2599:2592]} - {1'b0, layer_0_2[2599:2592]};
      top_2[1] = {1'b0,layer_1_2[2607:2600]} - {1'b0, layer_0_2[2607:2600]};
      top_2[2] = {1'b0,layer_1_2[2615:2608]} - {1'b0, layer_0_2[2615:2608]};
      mid_0[0] = {1'b0,layer_2_0[2599:2592]} - {1'b0, layer_1_0[2599:2592]};
      mid_0[1] = {1'b0,layer_2_0[2607:2600]} - {1'b0, layer_1_0[2607:2600]};
      mid_0[2] = {1'b0,layer_2_0[2615:2608]} - {1'b0, layer_1_0[2615:2608]};
      mid_1[0] = {1'b0,layer_2_1[2599:2592]} - {1'b0, layer_1_1[2599:2592]};
      mid_1[1] = {1'b0,layer_2_1[2607:2600]} - {1'b0, layer_1_1[2607:2600]};
      mid_1[2] = {1'b0,layer_2_1[2615:2608]} - {1'b0, layer_1_1[2615:2608]};
      mid_2[0] = {1'b0,layer_2_2[2599:2592]} - {1'b0, layer_1_2[2599:2592]};
      mid_2[1] = {1'b0,layer_2_2[2607:2600]} - {1'b0, layer_1_2[2607:2600]};
      mid_2[2] = {1'b0,layer_2_2[2615:2608]} - {1'b0, layer_1_2[2615:2608]};
      btm_0[0] = {1'b0,layer_3_0[2599:2592]} - {1'b0, layer_2_0[2599:2592]};
      btm_0[1] = {1'b0,layer_3_0[2607:2600]} - {1'b0, layer_2_0[2607:2600]};
      btm_0[2] = {1'b0,layer_3_0[2615:2608]} - {1'b0, layer_2_0[2615:2608]};
      btm_1[0] = {1'b0,layer_3_1[2599:2592]} - {1'b0, layer_2_1[2599:2592]};
      btm_1[1] = {1'b0,layer_3_1[2607:2600]} - {1'b0, layer_2_1[2607:2600]};
      btm_1[2] = {1'b0,layer_3_1[2615:2608]} - {1'b0, layer_2_1[2615:2608]};
      btm_2[0] = {1'b0,layer_3_2[2599:2592]} - {1'b0, layer_2_2[2599:2592]};
      btm_2[1] = {1'b0,layer_3_2[2607:2600]} - {1'b0, layer_2_2[2607:2600]};
      btm_2[2] = {1'b0,layer_3_2[2615:2608]} - {1'b0, layer_2_2[2615:2608]};
    end
    'd326: begin
      top_0[0] = {1'b0,layer_1_0[2607:2600]} - {1'b0, layer_0_0[2607:2600]};
      top_0[1] = {1'b0,layer_1_0[2615:2608]} - {1'b0, layer_0_0[2615:2608]};
      top_0[2] = {1'b0,layer_1_0[2623:2616]} - {1'b0, layer_0_0[2623:2616]};
      top_1[0] = {1'b0,layer_1_1[2607:2600]} - {1'b0, layer_0_1[2607:2600]};
      top_1[1] = {1'b0,layer_1_1[2615:2608]} - {1'b0, layer_0_1[2615:2608]};
      top_1[2] = {1'b0,layer_1_1[2623:2616]} - {1'b0, layer_0_1[2623:2616]};
      top_2[0] = {1'b0,layer_1_2[2607:2600]} - {1'b0, layer_0_2[2607:2600]};
      top_2[1] = {1'b0,layer_1_2[2615:2608]} - {1'b0, layer_0_2[2615:2608]};
      top_2[2] = {1'b0,layer_1_2[2623:2616]} - {1'b0, layer_0_2[2623:2616]};
      mid_0[0] = {1'b0,layer_2_0[2607:2600]} - {1'b0, layer_1_0[2607:2600]};
      mid_0[1] = {1'b0,layer_2_0[2615:2608]} - {1'b0, layer_1_0[2615:2608]};
      mid_0[2] = {1'b0,layer_2_0[2623:2616]} - {1'b0, layer_1_0[2623:2616]};
      mid_1[0] = {1'b0,layer_2_1[2607:2600]} - {1'b0, layer_1_1[2607:2600]};
      mid_1[1] = {1'b0,layer_2_1[2615:2608]} - {1'b0, layer_1_1[2615:2608]};
      mid_1[2] = {1'b0,layer_2_1[2623:2616]} - {1'b0, layer_1_1[2623:2616]};
      mid_2[0] = {1'b0,layer_2_2[2607:2600]} - {1'b0, layer_1_2[2607:2600]};
      mid_2[1] = {1'b0,layer_2_2[2615:2608]} - {1'b0, layer_1_2[2615:2608]};
      mid_2[2] = {1'b0,layer_2_2[2623:2616]} - {1'b0, layer_1_2[2623:2616]};
      btm_0[0] = {1'b0,layer_3_0[2607:2600]} - {1'b0, layer_2_0[2607:2600]};
      btm_0[1] = {1'b0,layer_3_0[2615:2608]} - {1'b0, layer_2_0[2615:2608]};
      btm_0[2] = {1'b0,layer_3_0[2623:2616]} - {1'b0, layer_2_0[2623:2616]};
      btm_1[0] = {1'b0,layer_3_1[2607:2600]} - {1'b0, layer_2_1[2607:2600]};
      btm_1[1] = {1'b0,layer_3_1[2615:2608]} - {1'b0, layer_2_1[2615:2608]};
      btm_1[2] = {1'b0,layer_3_1[2623:2616]} - {1'b0, layer_2_1[2623:2616]};
      btm_2[0] = {1'b0,layer_3_2[2607:2600]} - {1'b0, layer_2_2[2607:2600]};
      btm_2[1] = {1'b0,layer_3_2[2615:2608]} - {1'b0, layer_2_2[2615:2608]};
      btm_2[2] = {1'b0,layer_3_2[2623:2616]} - {1'b0, layer_2_2[2623:2616]};
    end
    'd327: begin
      top_0[0] = {1'b0,layer_1_0[2615:2608]} - {1'b0, layer_0_0[2615:2608]};
      top_0[1] = {1'b0,layer_1_0[2623:2616]} - {1'b0, layer_0_0[2623:2616]};
      top_0[2] = {1'b0,layer_1_0[2631:2624]} - {1'b0, layer_0_0[2631:2624]};
      top_1[0] = {1'b0,layer_1_1[2615:2608]} - {1'b0, layer_0_1[2615:2608]};
      top_1[1] = {1'b0,layer_1_1[2623:2616]} - {1'b0, layer_0_1[2623:2616]};
      top_1[2] = {1'b0,layer_1_1[2631:2624]} - {1'b0, layer_0_1[2631:2624]};
      top_2[0] = {1'b0,layer_1_2[2615:2608]} - {1'b0, layer_0_2[2615:2608]};
      top_2[1] = {1'b0,layer_1_2[2623:2616]} - {1'b0, layer_0_2[2623:2616]};
      top_2[2] = {1'b0,layer_1_2[2631:2624]} - {1'b0, layer_0_2[2631:2624]};
      mid_0[0] = {1'b0,layer_2_0[2615:2608]} - {1'b0, layer_1_0[2615:2608]};
      mid_0[1] = {1'b0,layer_2_0[2623:2616]} - {1'b0, layer_1_0[2623:2616]};
      mid_0[2] = {1'b0,layer_2_0[2631:2624]} - {1'b0, layer_1_0[2631:2624]};
      mid_1[0] = {1'b0,layer_2_1[2615:2608]} - {1'b0, layer_1_1[2615:2608]};
      mid_1[1] = {1'b0,layer_2_1[2623:2616]} - {1'b0, layer_1_1[2623:2616]};
      mid_1[2] = {1'b0,layer_2_1[2631:2624]} - {1'b0, layer_1_1[2631:2624]};
      mid_2[0] = {1'b0,layer_2_2[2615:2608]} - {1'b0, layer_1_2[2615:2608]};
      mid_2[1] = {1'b0,layer_2_2[2623:2616]} - {1'b0, layer_1_2[2623:2616]};
      mid_2[2] = {1'b0,layer_2_2[2631:2624]} - {1'b0, layer_1_2[2631:2624]};
      btm_0[0] = {1'b0,layer_3_0[2615:2608]} - {1'b0, layer_2_0[2615:2608]};
      btm_0[1] = {1'b0,layer_3_0[2623:2616]} - {1'b0, layer_2_0[2623:2616]};
      btm_0[2] = {1'b0,layer_3_0[2631:2624]} - {1'b0, layer_2_0[2631:2624]};
      btm_1[0] = {1'b0,layer_3_1[2615:2608]} - {1'b0, layer_2_1[2615:2608]};
      btm_1[1] = {1'b0,layer_3_1[2623:2616]} - {1'b0, layer_2_1[2623:2616]};
      btm_1[2] = {1'b0,layer_3_1[2631:2624]} - {1'b0, layer_2_1[2631:2624]};
      btm_2[0] = {1'b0,layer_3_2[2615:2608]} - {1'b0, layer_2_2[2615:2608]};
      btm_2[1] = {1'b0,layer_3_2[2623:2616]} - {1'b0, layer_2_2[2623:2616]};
      btm_2[2] = {1'b0,layer_3_2[2631:2624]} - {1'b0, layer_2_2[2631:2624]};
    end
    'd328: begin
      top_0[0] = {1'b0,layer_1_0[2623:2616]} - {1'b0, layer_0_0[2623:2616]};
      top_0[1] = {1'b0,layer_1_0[2631:2624]} - {1'b0, layer_0_0[2631:2624]};
      top_0[2] = {1'b0,layer_1_0[2639:2632]} - {1'b0, layer_0_0[2639:2632]};
      top_1[0] = {1'b0,layer_1_1[2623:2616]} - {1'b0, layer_0_1[2623:2616]};
      top_1[1] = {1'b0,layer_1_1[2631:2624]} - {1'b0, layer_0_1[2631:2624]};
      top_1[2] = {1'b0,layer_1_1[2639:2632]} - {1'b0, layer_0_1[2639:2632]};
      top_2[0] = {1'b0,layer_1_2[2623:2616]} - {1'b0, layer_0_2[2623:2616]};
      top_2[1] = {1'b0,layer_1_2[2631:2624]} - {1'b0, layer_0_2[2631:2624]};
      top_2[2] = {1'b0,layer_1_2[2639:2632]} - {1'b0, layer_0_2[2639:2632]};
      mid_0[0] = {1'b0,layer_2_0[2623:2616]} - {1'b0, layer_1_0[2623:2616]};
      mid_0[1] = {1'b0,layer_2_0[2631:2624]} - {1'b0, layer_1_0[2631:2624]};
      mid_0[2] = {1'b0,layer_2_0[2639:2632]} - {1'b0, layer_1_0[2639:2632]};
      mid_1[0] = {1'b0,layer_2_1[2623:2616]} - {1'b0, layer_1_1[2623:2616]};
      mid_1[1] = {1'b0,layer_2_1[2631:2624]} - {1'b0, layer_1_1[2631:2624]};
      mid_1[2] = {1'b0,layer_2_1[2639:2632]} - {1'b0, layer_1_1[2639:2632]};
      mid_2[0] = {1'b0,layer_2_2[2623:2616]} - {1'b0, layer_1_2[2623:2616]};
      mid_2[1] = {1'b0,layer_2_2[2631:2624]} - {1'b0, layer_1_2[2631:2624]};
      mid_2[2] = {1'b0,layer_2_2[2639:2632]} - {1'b0, layer_1_2[2639:2632]};
      btm_0[0] = {1'b0,layer_3_0[2623:2616]} - {1'b0, layer_2_0[2623:2616]};
      btm_0[1] = {1'b0,layer_3_0[2631:2624]} - {1'b0, layer_2_0[2631:2624]};
      btm_0[2] = {1'b0,layer_3_0[2639:2632]} - {1'b0, layer_2_0[2639:2632]};
      btm_1[0] = {1'b0,layer_3_1[2623:2616]} - {1'b0, layer_2_1[2623:2616]};
      btm_1[1] = {1'b0,layer_3_1[2631:2624]} - {1'b0, layer_2_1[2631:2624]};
      btm_1[2] = {1'b0,layer_3_1[2639:2632]} - {1'b0, layer_2_1[2639:2632]};
      btm_2[0] = {1'b0,layer_3_2[2623:2616]} - {1'b0, layer_2_2[2623:2616]};
      btm_2[1] = {1'b0,layer_3_2[2631:2624]} - {1'b0, layer_2_2[2631:2624]};
      btm_2[2] = {1'b0,layer_3_2[2639:2632]} - {1'b0, layer_2_2[2639:2632]};
    end
    'd329: begin
      top_0[0] = {1'b0,layer_1_0[2631:2624]} - {1'b0, layer_0_0[2631:2624]};
      top_0[1] = {1'b0,layer_1_0[2639:2632]} - {1'b0, layer_0_0[2639:2632]};
      top_0[2] = {1'b0,layer_1_0[2647:2640]} - {1'b0, layer_0_0[2647:2640]};
      top_1[0] = {1'b0,layer_1_1[2631:2624]} - {1'b0, layer_0_1[2631:2624]};
      top_1[1] = {1'b0,layer_1_1[2639:2632]} - {1'b0, layer_0_1[2639:2632]};
      top_1[2] = {1'b0,layer_1_1[2647:2640]} - {1'b0, layer_0_1[2647:2640]};
      top_2[0] = {1'b0,layer_1_2[2631:2624]} - {1'b0, layer_0_2[2631:2624]};
      top_2[1] = {1'b0,layer_1_2[2639:2632]} - {1'b0, layer_0_2[2639:2632]};
      top_2[2] = {1'b0,layer_1_2[2647:2640]} - {1'b0, layer_0_2[2647:2640]};
      mid_0[0] = {1'b0,layer_2_0[2631:2624]} - {1'b0, layer_1_0[2631:2624]};
      mid_0[1] = {1'b0,layer_2_0[2639:2632]} - {1'b0, layer_1_0[2639:2632]};
      mid_0[2] = {1'b0,layer_2_0[2647:2640]} - {1'b0, layer_1_0[2647:2640]};
      mid_1[0] = {1'b0,layer_2_1[2631:2624]} - {1'b0, layer_1_1[2631:2624]};
      mid_1[1] = {1'b0,layer_2_1[2639:2632]} - {1'b0, layer_1_1[2639:2632]};
      mid_1[2] = {1'b0,layer_2_1[2647:2640]} - {1'b0, layer_1_1[2647:2640]};
      mid_2[0] = {1'b0,layer_2_2[2631:2624]} - {1'b0, layer_1_2[2631:2624]};
      mid_2[1] = {1'b0,layer_2_2[2639:2632]} - {1'b0, layer_1_2[2639:2632]};
      mid_2[2] = {1'b0,layer_2_2[2647:2640]} - {1'b0, layer_1_2[2647:2640]};
      btm_0[0] = {1'b0,layer_3_0[2631:2624]} - {1'b0, layer_2_0[2631:2624]};
      btm_0[1] = {1'b0,layer_3_0[2639:2632]} - {1'b0, layer_2_0[2639:2632]};
      btm_0[2] = {1'b0,layer_3_0[2647:2640]} - {1'b0, layer_2_0[2647:2640]};
      btm_1[0] = {1'b0,layer_3_1[2631:2624]} - {1'b0, layer_2_1[2631:2624]};
      btm_1[1] = {1'b0,layer_3_1[2639:2632]} - {1'b0, layer_2_1[2639:2632]};
      btm_1[2] = {1'b0,layer_3_1[2647:2640]} - {1'b0, layer_2_1[2647:2640]};
      btm_2[0] = {1'b0,layer_3_2[2631:2624]} - {1'b0, layer_2_2[2631:2624]};
      btm_2[1] = {1'b0,layer_3_2[2639:2632]} - {1'b0, layer_2_2[2639:2632]};
      btm_2[2] = {1'b0,layer_3_2[2647:2640]} - {1'b0, layer_2_2[2647:2640]};
    end
    'd330: begin
      top_0[0] = {1'b0,layer_1_0[2639:2632]} - {1'b0, layer_0_0[2639:2632]};
      top_0[1] = {1'b0,layer_1_0[2647:2640]} - {1'b0, layer_0_0[2647:2640]};
      top_0[2] = {1'b0,layer_1_0[2655:2648]} - {1'b0, layer_0_0[2655:2648]};
      top_1[0] = {1'b0,layer_1_1[2639:2632]} - {1'b0, layer_0_1[2639:2632]};
      top_1[1] = {1'b0,layer_1_1[2647:2640]} - {1'b0, layer_0_1[2647:2640]};
      top_1[2] = {1'b0,layer_1_1[2655:2648]} - {1'b0, layer_0_1[2655:2648]};
      top_2[0] = {1'b0,layer_1_2[2639:2632]} - {1'b0, layer_0_2[2639:2632]};
      top_2[1] = {1'b0,layer_1_2[2647:2640]} - {1'b0, layer_0_2[2647:2640]};
      top_2[2] = {1'b0,layer_1_2[2655:2648]} - {1'b0, layer_0_2[2655:2648]};
      mid_0[0] = {1'b0,layer_2_0[2639:2632]} - {1'b0, layer_1_0[2639:2632]};
      mid_0[1] = {1'b0,layer_2_0[2647:2640]} - {1'b0, layer_1_0[2647:2640]};
      mid_0[2] = {1'b0,layer_2_0[2655:2648]} - {1'b0, layer_1_0[2655:2648]};
      mid_1[0] = {1'b0,layer_2_1[2639:2632]} - {1'b0, layer_1_1[2639:2632]};
      mid_1[1] = {1'b0,layer_2_1[2647:2640]} - {1'b0, layer_1_1[2647:2640]};
      mid_1[2] = {1'b0,layer_2_1[2655:2648]} - {1'b0, layer_1_1[2655:2648]};
      mid_2[0] = {1'b0,layer_2_2[2639:2632]} - {1'b0, layer_1_2[2639:2632]};
      mid_2[1] = {1'b0,layer_2_2[2647:2640]} - {1'b0, layer_1_2[2647:2640]};
      mid_2[2] = {1'b0,layer_2_2[2655:2648]} - {1'b0, layer_1_2[2655:2648]};
      btm_0[0] = {1'b0,layer_3_0[2639:2632]} - {1'b0, layer_2_0[2639:2632]};
      btm_0[1] = {1'b0,layer_3_0[2647:2640]} - {1'b0, layer_2_0[2647:2640]};
      btm_0[2] = {1'b0,layer_3_0[2655:2648]} - {1'b0, layer_2_0[2655:2648]};
      btm_1[0] = {1'b0,layer_3_1[2639:2632]} - {1'b0, layer_2_1[2639:2632]};
      btm_1[1] = {1'b0,layer_3_1[2647:2640]} - {1'b0, layer_2_1[2647:2640]};
      btm_1[2] = {1'b0,layer_3_1[2655:2648]} - {1'b0, layer_2_1[2655:2648]};
      btm_2[0] = {1'b0,layer_3_2[2639:2632]} - {1'b0, layer_2_2[2639:2632]};
      btm_2[1] = {1'b0,layer_3_2[2647:2640]} - {1'b0, layer_2_2[2647:2640]};
      btm_2[2] = {1'b0,layer_3_2[2655:2648]} - {1'b0, layer_2_2[2655:2648]};
    end
    'd331: begin
      top_0[0] = {1'b0,layer_1_0[2647:2640]} - {1'b0, layer_0_0[2647:2640]};
      top_0[1] = {1'b0,layer_1_0[2655:2648]} - {1'b0, layer_0_0[2655:2648]};
      top_0[2] = {1'b0,layer_1_0[2663:2656]} - {1'b0, layer_0_0[2663:2656]};
      top_1[0] = {1'b0,layer_1_1[2647:2640]} - {1'b0, layer_0_1[2647:2640]};
      top_1[1] = {1'b0,layer_1_1[2655:2648]} - {1'b0, layer_0_1[2655:2648]};
      top_1[2] = {1'b0,layer_1_1[2663:2656]} - {1'b0, layer_0_1[2663:2656]};
      top_2[0] = {1'b0,layer_1_2[2647:2640]} - {1'b0, layer_0_2[2647:2640]};
      top_2[1] = {1'b0,layer_1_2[2655:2648]} - {1'b0, layer_0_2[2655:2648]};
      top_2[2] = {1'b0,layer_1_2[2663:2656]} - {1'b0, layer_0_2[2663:2656]};
      mid_0[0] = {1'b0,layer_2_0[2647:2640]} - {1'b0, layer_1_0[2647:2640]};
      mid_0[1] = {1'b0,layer_2_0[2655:2648]} - {1'b0, layer_1_0[2655:2648]};
      mid_0[2] = {1'b0,layer_2_0[2663:2656]} - {1'b0, layer_1_0[2663:2656]};
      mid_1[0] = {1'b0,layer_2_1[2647:2640]} - {1'b0, layer_1_1[2647:2640]};
      mid_1[1] = {1'b0,layer_2_1[2655:2648]} - {1'b0, layer_1_1[2655:2648]};
      mid_1[2] = {1'b0,layer_2_1[2663:2656]} - {1'b0, layer_1_1[2663:2656]};
      mid_2[0] = {1'b0,layer_2_2[2647:2640]} - {1'b0, layer_1_2[2647:2640]};
      mid_2[1] = {1'b0,layer_2_2[2655:2648]} - {1'b0, layer_1_2[2655:2648]};
      mid_2[2] = {1'b0,layer_2_2[2663:2656]} - {1'b0, layer_1_2[2663:2656]};
      btm_0[0] = {1'b0,layer_3_0[2647:2640]} - {1'b0, layer_2_0[2647:2640]};
      btm_0[1] = {1'b0,layer_3_0[2655:2648]} - {1'b0, layer_2_0[2655:2648]};
      btm_0[2] = {1'b0,layer_3_0[2663:2656]} - {1'b0, layer_2_0[2663:2656]};
      btm_1[0] = {1'b0,layer_3_1[2647:2640]} - {1'b0, layer_2_1[2647:2640]};
      btm_1[1] = {1'b0,layer_3_1[2655:2648]} - {1'b0, layer_2_1[2655:2648]};
      btm_1[2] = {1'b0,layer_3_1[2663:2656]} - {1'b0, layer_2_1[2663:2656]};
      btm_2[0] = {1'b0,layer_3_2[2647:2640]} - {1'b0, layer_2_2[2647:2640]};
      btm_2[1] = {1'b0,layer_3_2[2655:2648]} - {1'b0, layer_2_2[2655:2648]};
      btm_2[2] = {1'b0,layer_3_2[2663:2656]} - {1'b0, layer_2_2[2663:2656]};
    end
    'd332: begin
      top_0[0] = {1'b0,layer_1_0[2655:2648]} - {1'b0, layer_0_0[2655:2648]};
      top_0[1] = {1'b0,layer_1_0[2663:2656]} - {1'b0, layer_0_0[2663:2656]};
      top_0[2] = {1'b0,layer_1_0[2671:2664]} - {1'b0, layer_0_0[2671:2664]};
      top_1[0] = {1'b0,layer_1_1[2655:2648]} - {1'b0, layer_0_1[2655:2648]};
      top_1[1] = {1'b0,layer_1_1[2663:2656]} - {1'b0, layer_0_1[2663:2656]};
      top_1[2] = {1'b0,layer_1_1[2671:2664]} - {1'b0, layer_0_1[2671:2664]};
      top_2[0] = {1'b0,layer_1_2[2655:2648]} - {1'b0, layer_0_2[2655:2648]};
      top_2[1] = {1'b0,layer_1_2[2663:2656]} - {1'b0, layer_0_2[2663:2656]};
      top_2[2] = {1'b0,layer_1_2[2671:2664]} - {1'b0, layer_0_2[2671:2664]};
      mid_0[0] = {1'b0,layer_2_0[2655:2648]} - {1'b0, layer_1_0[2655:2648]};
      mid_0[1] = {1'b0,layer_2_0[2663:2656]} - {1'b0, layer_1_0[2663:2656]};
      mid_0[2] = {1'b0,layer_2_0[2671:2664]} - {1'b0, layer_1_0[2671:2664]};
      mid_1[0] = {1'b0,layer_2_1[2655:2648]} - {1'b0, layer_1_1[2655:2648]};
      mid_1[1] = {1'b0,layer_2_1[2663:2656]} - {1'b0, layer_1_1[2663:2656]};
      mid_1[2] = {1'b0,layer_2_1[2671:2664]} - {1'b0, layer_1_1[2671:2664]};
      mid_2[0] = {1'b0,layer_2_2[2655:2648]} - {1'b0, layer_1_2[2655:2648]};
      mid_2[1] = {1'b0,layer_2_2[2663:2656]} - {1'b0, layer_1_2[2663:2656]};
      mid_2[2] = {1'b0,layer_2_2[2671:2664]} - {1'b0, layer_1_2[2671:2664]};
      btm_0[0] = {1'b0,layer_3_0[2655:2648]} - {1'b0, layer_2_0[2655:2648]};
      btm_0[1] = {1'b0,layer_3_0[2663:2656]} - {1'b0, layer_2_0[2663:2656]};
      btm_0[2] = {1'b0,layer_3_0[2671:2664]} - {1'b0, layer_2_0[2671:2664]};
      btm_1[0] = {1'b0,layer_3_1[2655:2648]} - {1'b0, layer_2_1[2655:2648]};
      btm_1[1] = {1'b0,layer_3_1[2663:2656]} - {1'b0, layer_2_1[2663:2656]};
      btm_1[2] = {1'b0,layer_3_1[2671:2664]} - {1'b0, layer_2_1[2671:2664]};
      btm_2[0] = {1'b0,layer_3_2[2655:2648]} - {1'b0, layer_2_2[2655:2648]};
      btm_2[1] = {1'b0,layer_3_2[2663:2656]} - {1'b0, layer_2_2[2663:2656]};
      btm_2[2] = {1'b0,layer_3_2[2671:2664]} - {1'b0, layer_2_2[2671:2664]};
    end
    'd333: begin
      top_0[0] = {1'b0,layer_1_0[2663:2656]} - {1'b0, layer_0_0[2663:2656]};
      top_0[1] = {1'b0,layer_1_0[2671:2664]} - {1'b0, layer_0_0[2671:2664]};
      top_0[2] = {1'b0,layer_1_0[2679:2672]} - {1'b0, layer_0_0[2679:2672]};
      top_1[0] = {1'b0,layer_1_1[2663:2656]} - {1'b0, layer_0_1[2663:2656]};
      top_1[1] = {1'b0,layer_1_1[2671:2664]} - {1'b0, layer_0_1[2671:2664]};
      top_1[2] = {1'b0,layer_1_1[2679:2672]} - {1'b0, layer_0_1[2679:2672]};
      top_2[0] = {1'b0,layer_1_2[2663:2656]} - {1'b0, layer_0_2[2663:2656]};
      top_2[1] = {1'b0,layer_1_2[2671:2664]} - {1'b0, layer_0_2[2671:2664]};
      top_2[2] = {1'b0,layer_1_2[2679:2672]} - {1'b0, layer_0_2[2679:2672]};
      mid_0[0] = {1'b0,layer_2_0[2663:2656]} - {1'b0, layer_1_0[2663:2656]};
      mid_0[1] = {1'b0,layer_2_0[2671:2664]} - {1'b0, layer_1_0[2671:2664]};
      mid_0[2] = {1'b0,layer_2_0[2679:2672]} - {1'b0, layer_1_0[2679:2672]};
      mid_1[0] = {1'b0,layer_2_1[2663:2656]} - {1'b0, layer_1_1[2663:2656]};
      mid_1[1] = {1'b0,layer_2_1[2671:2664]} - {1'b0, layer_1_1[2671:2664]};
      mid_1[2] = {1'b0,layer_2_1[2679:2672]} - {1'b0, layer_1_1[2679:2672]};
      mid_2[0] = {1'b0,layer_2_2[2663:2656]} - {1'b0, layer_1_2[2663:2656]};
      mid_2[1] = {1'b0,layer_2_2[2671:2664]} - {1'b0, layer_1_2[2671:2664]};
      mid_2[2] = {1'b0,layer_2_2[2679:2672]} - {1'b0, layer_1_2[2679:2672]};
      btm_0[0] = {1'b0,layer_3_0[2663:2656]} - {1'b0, layer_2_0[2663:2656]};
      btm_0[1] = {1'b0,layer_3_0[2671:2664]} - {1'b0, layer_2_0[2671:2664]};
      btm_0[2] = {1'b0,layer_3_0[2679:2672]} - {1'b0, layer_2_0[2679:2672]};
      btm_1[0] = {1'b0,layer_3_1[2663:2656]} - {1'b0, layer_2_1[2663:2656]};
      btm_1[1] = {1'b0,layer_3_1[2671:2664]} - {1'b0, layer_2_1[2671:2664]};
      btm_1[2] = {1'b0,layer_3_1[2679:2672]} - {1'b0, layer_2_1[2679:2672]};
      btm_2[0] = {1'b0,layer_3_2[2663:2656]} - {1'b0, layer_2_2[2663:2656]};
      btm_2[1] = {1'b0,layer_3_2[2671:2664]} - {1'b0, layer_2_2[2671:2664]};
      btm_2[2] = {1'b0,layer_3_2[2679:2672]} - {1'b0, layer_2_2[2679:2672]};
    end
    'd334: begin
      top_0[0] = {1'b0,layer_1_0[2671:2664]} - {1'b0, layer_0_0[2671:2664]};
      top_0[1] = {1'b0,layer_1_0[2679:2672]} - {1'b0, layer_0_0[2679:2672]};
      top_0[2] = {1'b0,layer_1_0[2687:2680]} - {1'b0, layer_0_0[2687:2680]};
      top_1[0] = {1'b0,layer_1_1[2671:2664]} - {1'b0, layer_0_1[2671:2664]};
      top_1[1] = {1'b0,layer_1_1[2679:2672]} - {1'b0, layer_0_1[2679:2672]};
      top_1[2] = {1'b0,layer_1_1[2687:2680]} - {1'b0, layer_0_1[2687:2680]};
      top_2[0] = {1'b0,layer_1_2[2671:2664]} - {1'b0, layer_0_2[2671:2664]};
      top_2[1] = {1'b0,layer_1_2[2679:2672]} - {1'b0, layer_0_2[2679:2672]};
      top_2[2] = {1'b0,layer_1_2[2687:2680]} - {1'b0, layer_0_2[2687:2680]};
      mid_0[0] = {1'b0,layer_2_0[2671:2664]} - {1'b0, layer_1_0[2671:2664]};
      mid_0[1] = {1'b0,layer_2_0[2679:2672]} - {1'b0, layer_1_0[2679:2672]};
      mid_0[2] = {1'b0,layer_2_0[2687:2680]} - {1'b0, layer_1_0[2687:2680]};
      mid_1[0] = {1'b0,layer_2_1[2671:2664]} - {1'b0, layer_1_1[2671:2664]};
      mid_1[1] = {1'b0,layer_2_1[2679:2672]} - {1'b0, layer_1_1[2679:2672]};
      mid_1[2] = {1'b0,layer_2_1[2687:2680]} - {1'b0, layer_1_1[2687:2680]};
      mid_2[0] = {1'b0,layer_2_2[2671:2664]} - {1'b0, layer_1_2[2671:2664]};
      mid_2[1] = {1'b0,layer_2_2[2679:2672]} - {1'b0, layer_1_2[2679:2672]};
      mid_2[2] = {1'b0,layer_2_2[2687:2680]} - {1'b0, layer_1_2[2687:2680]};
      btm_0[0] = {1'b0,layer_3_0[2671:2664]} - {1'b0, layer_2_0[2671:2664]};
      btm_0[1] = {1'b0,layer_3_0[2679:2672]} - {1'b0, layer_2_0[2679:2672]};
      btm_0[2] = {1'b0,layer_3_0[2687:2680]} - {1'b0, layer_2_0[2687:2680]};
      btm_1[0] = {1'b0,layer_3_1[2671:2664]} - {1'b0, layer_2_1[2671:2664]};
      btm_1[1] = {1'b0,layer_3_1[2679:2672]} - {1'b0, layer_2_1[2679:2672]};
      btm_1[2] = {1'b0,layer_3_1[2687:2680]} - {1'b0, layer_2_1[2687:2680]};
      btm_2[0] = {1'b0,layer_3_2[2671:2664]} - {1'b0, layer_2_2[2671:2664]};
      btm_2[1] = {1'b0,layer_3_2[2679:2672]} - {1'b0, layer_2_2[2679:2672]};
      btm_2[2] = {1'b0,layer_3_2[2687:2680]} - {1'b0, layer_2_2[2687:2680]};
    end
    'd335: begin
      top_0[0] = {1'b0,layer_1_0[2679:2672]} - {1'b0, layer_0_0[2679:2672]};
      top_0[1] = {1'b0,layer_1_0[2687:2680]} - {1'b0, layer_0_0[2687:2680]};
      top_0[2] = {1'b0,layer_1_0[2695:2688]} - {1'b0, layer_0_0[2695:2688]};
      top_1[0] = {1'b0,layer_1_1[2679:2672]} - {1'b0, layer_0_1[2679:2672]};
      top_1[1] = {1'b0,layer_1_1[2687:2680]} - {1'b0, layer_0_1[2687:2680]};
      top_1[2] = {1'b0,layer_1_1[2695:2688]} - {1'b0, layer_0_1[2695:2688]};
      top_2[0] = {1'b0,layer_1_2[2679:2672]} - {1'b0, layer_0_2[2679:2672]};
      top_2[1] = {1'b0,layer_1_2[2687:2680]} - {1'b0, layer_0_2[2687:2680]};
      top_2[2] = {1'b0,layer_1_2[2695:2688]} - {1'b0, layer_0_2[2695:2688]};
      mid_0[0] = {1'b0,layer_2_0[2679:2672]} - {1'b0, layer_1_0[2679:2672]};
      mid_0[1] = {1'b0,layer_2_0[2687:2680]} - {1'b0, layer_1_0[2687:2680]};
      mid_0[2] = {1'b0,layer_2_0[2695:2688]} - {1'b0, layer_1_0[2695:2688]};
      mid_1[0] = {1'b0,layer_2_1[2679:2672]} - {1'b0, layer_1_1[2679:2672]};
      mid_1[1] = {1'b0,layer_2_1[2687:2680]} - {1'b0, layer_1_1[2687:2680]};
      mid_1[2] = {1'b0,layer_2_1[2695:2688]} - {1'b0, layer_1_1[2695:2688]};
      mid_2[0] = {1'b0,layer_2_2[2679:2672]} - {1'b0, layer_1_2[2679:2672]};
      mid_2[1] = {1'b0,layer_2_2[2687:2680]} - {1'b0, layer_1_2[2687:2680]};
      mid_2[2] = {1'b0,layer_2_2[2695:2688]} - {1'b0, layer_1_2[2695:2688]};
      btm_0[0] = {1'b0,layer_3_0[2679:2672]} - {1'b0, layer_2_0[2679:2672]};
      btm_0[1] = {1'b0,layer_3_0[2687:2680]} - {1'b0, layer_2_0[2687:2680]};
      btm_0[2] = {1'b0,layer_3_0[2695:2688]} - {1'b0, layer_2_0[2695:2688]};
      btm_1[0] = {1'b0,layer_3_1[2679:2672]} - {1'b0, layer_2_1[2679:2672]};
      btm_1[1] = {1'b0,layer_3_1[2687:2680]} - {1'b0, layer_2_1[2687:2680]};
      btm_1[2] = {1'b0,layer_3_1[2695:2688]} - {1'b0, layer_2_1[2695:2688]};
      btm_2[0] = {1'b0,layer_3_2[2679:2672]} - {1'b0, layer_2_2[2679:2672]};
      btm_2[1] = {1'b0,layer_3_2[2687:2680]} - {1'b0, layer_2_2[2687:2680]};
      btm_2[2] = {1'b0,layer_3_2[2695:2688]} - {1'b0, layer_2_2[2695:2688]};
    end
    'd336: begin
      top_0[0] = {1'b0,layer_1_0[2687:2680]} - {1'b0, layer_0_0[2687:2680]};
      top_0[1] = {1'b0,layer_1_0[2695:2688]} - {1'b0, layer_0_0[2695:2688]};
      top_0[2] = {1'b0,layer_1_0[2703:2696]} - {1'b0, layer_0_0[2703:2696]};
      top_1[0] = {1'b0,layer_1_1[2687:2680]} - {1'b0, layer_0_1[2687:2680]};
      top_1[1] = {1'b0,layer_1_1[2695:2688]} - {1'b0, layer_0_1[2695:2688]};
      top_1[2] = {1'b0,layer_1_1[2703:2696]} - {1'b0, layer_0_1[2703:2696]};
      top_2[0] = {1'b0,layer_1_2[2687:2680]} - {1'b0, layer_0_2[2687:2680]};
      top_2[1] = {1'b0,layer_1_2[2695:2688]} - {1'b0, layer_0_2[2695:2688]};
      top_2[2] = {1'b0,layer_1_2[2703:2696]} - {1'b0, layer_0_2[2703:2696]};
      mid_0[0] = {1'b0,layer_2_0[2687:2680]} - {1'b0, layer_1_0[2687:2680]};
      mid_0[1] = {1'b0,layer_2_0[2695:2688]} - {1'b0, layer_1_0[2695:2688]};
      mid_0[2] = {1'b0,layer_2_0[2703:2696]} - {1'b0, layer_1_0[2703:2696]};
      mid_1[0] = {1'b0,layer_2_1[2687:2680]} - {1'b0, layer_1_1[2687:2680]};
      mid_1[1] = {1'b0,layer_2_1[2695:2688]} - {1'b0, layer_1_1[2695:2688]};
      mid_1[2] = {1'b0,layer_2_1[2703:2696]} - {1'b0, layer_1_1[2703:2696]};
      mid_2[0] = {1'b0,layer_2_2[2687:2680]} - {1'b0, layer_1_2[2687:2680]};
      mid_2[1] = {1'b0,layer_2_2[2695:2688]} - {1'b0, layer_1_2[2695:2688]};
      mid_2[2] = {1'b0,layer_2_2[2703:2696]} - {1'b0, layer_1_2[2703:2696]};
      btm_0[0] = {1'b0,layer_3_0[2687:2680]} - {1'b0, layer_2_0[2687:2680]};
      btm_0[1] = {1'b0,layer_3_0[2695:2688]} - {1'b0, layer_2_0[2695:2688]};
      btm_0[2] = {1'b0,layer_3_0[2703:2696]} - {1'b0, layer_2_0[2703:2696]};
      btm_1[0] = {1'b0,layer_3_1[2687:2680]} - {1'b0, layer_2_1[2687:2680]};
      btm_1[1] = {1'b0,layer_3_1[2695:2688]} - {1'b0, layer_2_1[2695:2688]};
      btm_1[2] = {1'b0,layer_3_1[2703:2696]} - {1'b0, layer_2_1[2703:2696]};
      btm_2[0] = {1'b0,layer_3_2[2687:2680]} - {1'b0, layer_2_2[2687:2680]};
      btm_2[1] = {1'b0,layer_3_2[2695:2688]} - {1'b0, layer_2_2[2695:2688]};
      btm_2[2] = {1'b0,layer_3_2[2703:2696]} - {1'b0, layer_2_2[2703:2696]};
    end
    'd337: begin
      top_0[0] = {1'b0,layer_1_0[2695:2688]} - {1'b0, layer_0_0[2695:2688]};
      top_0[1] = {1'b0,layer_1_0[2703:2696]} - {1'b0, layer_0_0[2703:2696]};
      top_0[2] = {1'b0,layer_1_0[2711:2704]} - {1'b0, layer_0_0[2711:2704]};
      top_1[0] = {1'b0,layer_1_1[2695:2688]} - {1'b0, layer_0_1[2695:2688]};
      top_1[1] = {1'b0,layer_1_1[2703:2696]} - {1'b0, layer_0_1[2703:2696]};
      top_1[2] = {1'b0,layer_1_1[2711:2704]} - {1'b0, layer_0_1[2711:2704]};
      top_2[0] = {1'b0,layer_1_2[2695:2688]} - {1'b0, layer_0_2[2695:2688]};
      top_2[1] = {1'b0,layer_1_2[2703:2696]} - {1'b0, layer_0_2[2703:2696]};
      top_2[2] = {1'b0,layer_1_2[2711:2704]} - {1'b0, layer_0_2[2711:2704]};
      mid_0[0] = {1'b0,layer_2_0[2695:2688]} - {1'b0, layer_1_0[2695:2688]};
      mid_0[1] = {1'b0,layer_2_0[2703:2696]} - {1'b0, layer_1_0[2703:2696]};
      mid_0[2] = {1'b0,layer_2_0[2711:2704]} - {1'b0, layer_1_0[2711:2704]};
      mid_1[0] = {1'b0,layer_2_1[2695:2688]} - {1'b0, layer_1_1[2695:2688]};
      mid_1[1] = {1'b0,layer_2_1[2703:2696]} - {1'b0, layer_1_1[2703:2696]};
      mid_1[2] = {1'b0,layer_2_1[2711:2704]} - {1'b0, layer_1_1[2711:2704]};
      mid_2[0] = {1'b0,layer_2_2[2695:2688]} - {1'b0, layer_1_2[2695:2688]};
      mid_2[1] = {1'b0,layer_2_2[2703:2696]} - {1'b0, layer_1_2[2703:2696]};
      mid_2[2] = {1'b0,layer_2_2[2711:2704]} - {1'b0, layer_1_2[2711:2704]};
      btm_0[0] = {1'b0,layer_3_0[2695:2688]} - {1'b0, layer_2_0[2695:2688]};
      btm_0[1] = {1'b0,layer_3_0[2703:2696]} - {1'b0, layer_2_0[2703:2696]};
      btm_0[2] = {1'b0,layer_3_0[2711:2704]} - {1'b0, layer_2_0[2711:2704]};
      btm_1[0] = {1'b0,layer_3_1[2695:2688]} - {1'b0, layer_2_1[2695:2688]};
      btm_1[1] = {1'b0,layer_3_1[2703:2696]} - {1'b0, layer_2_1[2703:2696]};
      btm_1[2] = {1'b0,layer_3_1[2711:2704]} - {1'b0, layer_2_1[2711:2704]};
      btm_2[0] = {1'b0,layer_3_2[2695:2688]} - {1'b0, layer_2_2[2695:2688]};
      btm_2[1] = {1'b0,layer_3_2[2703:2696]} - {1'b0, layer_2_2[2703:2696]};
      btm_2[2] = {1'b0,layer_3_2[2711:2704]} - {1'b0, layer_2_2[2711:2704]};
    end
    'd338: begin
      top_0[0] = {1'b0,layer_1_0[2703:2696]} - {1'b0, layer_0_0[2703:2696]};
      top_0[1] = {1'b0,layer_1_0[2711:2704]} - {1'b0, layer_0_0[2711:2704]};
      top_0[2] = {1'b0,layer_1_0[2719:2712]} - {1'b0, layer_0_0[2719:2712]};
      top_1[0] = {1'b0,layer_1_1[2703:2696]} - {1'b0, layer_0_1[2703:2696]};
      top_1[1] = {1'b0,layer_1_1[2711:2704]} - {1'b0, layer_0_1[2711:2704]};
      top_1[2] = {1'b0,layer_1_1[2719:2712]} - {1'b0, layer_0_1[2719:2712]};
      top_2[0] = {1'b0,layer_1_2[2703:2696]} - {1'b0, layer_0_2[2703:2696]};
      top_2[1] = {1'b0,layer_1_2[2711:2704]} - {1'b0, layer_0_2[2711:2704]};
      top_2[2] = {1'b0,layer_1_2[2719:2712]} - {1'b0, layer_0_2[2719:2712]};
      mid_0[0] = {1'b0,layer_2_0[2703:2696]} - {1'b0, layer_1_0[2703:2696]};
      mid_0[1] = {1'b0,layer_2_0[2711:2704]} - {1'b0, layer_1_0[2711:2704]};
      mid_0[2] = {1'b0,layer_2_0[2719:2712]} - {1'b0, layer_1_0[2719:2712]};
      mid_1[0] = {1'b0,layer_2_1[2703:2696]} - {1'b0, layer_1_1[2703:2696]};
      mid_1[1] = {1'b0,layer_2_1[2711:2704]} - {1'b0, layer_1_1[2711:2704]};
      mid_1[2] = {1'b0,layer_2_1[2719:2712]} - {1'b0, layer_1_1[2719:2712]};
      mid_2[0] = {1'b0,layer_2_2[2703:2696]} - {1'b0, layer_1_2[2703:2696]};
      mid_2[1] = {1'b0,layer_2_2[2711:2704]} - {1'b0, layer_1_2[2711:2704]};
      mid_2[2] = {1'b0,layer_2_2[2719:2712]} - {1'b0, layer_1_2[2719:2712]};
      btm_0[0] = {1'b0,layer_3_0[2703:2696]} - {1'b0, layer_2_0[2703:2696]};
      btm_0[1] = {1'b0,layer_3_0[2711:2704]} - {1'b0, layer_2_0[2711:2704]};
      btm_0[2] = {1'b0,layer_3_0[2719:2712]} - {1'b0, layer_2_0[2719:2712]};
      btm_1[0] = {1'b0,layer_3_1[2703:2696]} - {1'b0, layer_2_1[2703:2696]};
      btm_1[1] = {1'b0,layer_3_1[2711:2704]} - {1'b0, layer_2_1[2711:2704]};
      btm_1[2] = {1'b0,layer_3_1[2719:2712]} - {1'b0, layer_2_1[2719:2712]};
      btm_2[0] = {1'b0,layer_3_2[2703:2696]} - {1'b0, layer_2_2[2703:2696]};
      btm_2[1] = {1'b0,layer_3_2[2711:2704]} - {1'b0, layer_2_2[2711:2704]};
      btm_2[2] = {1'b0,layer_3_2[2719:2712]} - {1'b0, layer_2_2[2719:2712]};
    end
    'd339: begin
      top_0[0] = {1'b0,layer_1_0[2711:2704]} - {1'b0, layer_0_0[2711:2704]};
      top_0[1] = {1'b0,layer_1_0[2719:2712]} - {1'b0, layer_0_0[2719:2712]};
      top_0[2] = {1'b0,layer_1_0[2727:2720]} - {1'b0, layer_0_0[2727:2720]};
      top_1[0] = {1'b0,layer_1_1[2711:2704]} - {1'b0, layer_0_1[2711:2704]};
      top_1[1] = {1'b0,layer_1_1[2719:2712]} - {1'b0, layer_0_1[2719:2712]};
      top_1[2] = {1'b0,layer_1_1[2727:2720]} - {1'b0, layer_0_1[2727:2720]};
      top_2[0] = {1'b0,layer_1_2[2711:2704]} - {1'b0, layer_0_2[2711:2704]};
      top_2[1] = {1'b0,layer_1_2[2719:2712]} - {1'b0, layer_0_2[2719:2712]};
      top_2[2] = {1'b0,layer_1_2[2727:2720]} - {1'b0, layer_0_2[2727:2720]};
      mid_0[0] = {1'b0,layer_2_0[2711:2704]} - {1'b0, layer_1_0[2711:2704]};
      mid_0[1] = {1'b0,layer_2_0[2719:2712]} - {1'b0, layer_1_0[2719:2712]};
      mid_0[2] = {1'b0,layer_2_0[2727:2720]} - {1'b0, layer_1_0[2727:2720]};
      mid_1[0] = {1'b0,layer_2_1[2711:2704]} - {1'b0, layer_1_1[2711:2704]};
      mid_1[1] = {1'b0,layer_2_1[2719:2712]} - {1'b0, layer_1_1[2719:2712]};
      mid_1[2] = {1'b0,layer_2_1[2727:2720]} - {1'b0, layer_1_1[2727:2720]};
      mid_2[0] = {1'b0,layer_2_2[2711:2704]} - {1'b0, layer_1_2[2711:2704]};
      mid_2[1] = {1'b0,layer_2_2[2719:2712]} - {1'b0, layer_1_2[2719:2712]};
      mid_2[2] = {1'b0,layer_2_2[2727:2720]} - {1'b0, layer_1_2[2727:2720]};
      btm_0[0] = {1'b0,layer_3_0[2711:2704]} - {1'b0, layer_2_0[2711:2704]};
      btm_0[1] = {1'b0,layer_3_0[2719:2712]} - {1'b0, layer_2_0[2719:2712]};
      btm_0[2] = {1'b0,layer_3_0[2727:2720]} - {1'b0, layer_2_0[2727:2720]};
      btm_1[0] = {1'b0,layer_3_1[2711:2704]} - {1'b0, layer_2_1[2711:2704]};
      btm_1[1] = {1'b0,layer_3_1[2719:2712]} - {1'b0, layer_2_1[2719:2712]};
      btm_1[2] = {1'b0,layer_3_1[2727:2720]} - {1'b0, layer_2_1[2727:2720]};
      btm_2[0] = {1'b0,layer_3_2[2711:2704]} - {1'b0, layer_2_2[2711:2704]};
      btm_2[1] = {1'b0,layer_3_2[2719:2712]} - {1'b0, layer_2_2[2719:2712]};
      btm_2[2] = {1'b0,layer_3_2[2727:2720]} - {1'b0, layer_2_2[2727:2720]};
    end
    'd340: begin
      top_0[0] = {1'b0,layer_1_0[2719:2712]} - {1'b0, layer_0_0[2719:2712]};
      top_0[1] = {1'b0,layer_1_0[2727:2720]} - {1'b0, layer_0_0[2727:2720]};
      top_0[2] = {1'b0,layer_1_0[2735:2728]} - {1'b0, layer_0_0[2735:2728]};
      top_1[0] = {1'b0,layer_1_1[2719:2712]} - {1'b0, layer_0_1[2719:2712]};
      top_1[1] = {1'b0,layer_1_1[2727:2720]} - {1'b0, layer_0_1[2727:2720]};
      top_1[2] = {1'b0,layer_1_1[2735:2728]} - {1'b0, layer_0_1[2735:2728]};
      top_2[0] = {1'b0,layer_1_2[2719:2712]} - {1'b0, layer_0_2[2719:2712]};
      top_2[1] = {1'b0,layer_1_2[2727:2720]} - {1'b0, layer_0_2[2727:2720]};
      top_2[2] = {1'b0,layer_1_2[2735:2728]} - {1'b0, layer_0_2[2735:2728]};
      mid_0[0] = {1'b0,layer_2_0[2719:2712]} - {1'b0, layer_1_0[2719:2712]};
      mid_0[1] = {1'b0,layer_2_0[2727:2720]} - {1'b0, layer_1_0[2727:2720]};
      mid_0[2] = {1'b0,layer_2_0[2735:2728]} - {1'b0, layer_1_0[2735:2728]};
      mid_1[0] = {1'b0,layer_2_1[2719:2712]} - {1'b0, layer_1_1[2719:2712]};
      mid_1[1] = {1'b0,layer_2_1[2727:2720]} - {1'b0, layer_1_1[2727:2720]};
      mid_1[2] = {1'b0,layer_2_1[2735:2728]} - {1'b0, layer_1_1[2735:2728]};
      mid_2[0] = {1'b0,layer_2_2[2719:2712]} - {1'b0, layer_1_2[2719:2712]};
      mid_2[1] = {1'b0,layer_2_2[2727:2720]} - {1'b0, layer_1_2[2727:2720]};
      mid_2[2] = {1'b0,layer_2_2[2735:2728]} - {1'b0, layer_1_2[2735:2728]};
      btm_0[0] = {1'b0,layer_3_0[2719:2712]} - {1'b0, layer_2_0[2719:2712]};
      btm_0[1] = {1'b0,layer_3_0[2727:2720]} - {1'b0, layer_2_0[2727:2720]};
      btm_0[2] = {1'b0,layer_3_0[2735:2728]} - {1'b0, layer_2_0[2735:2728]};
      btm_1[0] = {1'b0,layer_3_1[2719:2712]} - {1'b0, layer_2_1[2719:2712]};
      btm_1[1] = {1'b0,layer_3_1[2727:2720]} - {1'b0, layer_2_1[2727:2720]};
      btm_1[2] = {1'b0,layer_3_1[2735:2728]} - {1'b0, layer_2_1[2735:2728]};
      btm_2[0] = {1'b0,layer_3_2[2719:2712]} - {1'b0, layer_2_2[2719:2712]};
      btm_2[1] = {1'b0,layer_3_2[2727:2720]} - {1'b0, layer_2_2[2727:2720]};
      btm_2[2] = {1'b0,layer_3_2[2735:2728]} - {1'b0, layer_2_2[2735:2728]};
    end
    'd341: begin
      top_0[0] = {1'b0,layer_1_0[2727:2720]} - {1'b0, layer_0_0[2727:2720]};
      top_0[1] = {1'b0,layer_1_0[2735:2728]} - {1'b0, layer_0_0[2735:2728]};
      top_0[2] = {1'b0,layer_1_0[2743:2736]} - {1'b0, layer_0_0[2743:2736]};
      top_1[0] = {1'b0,layer_1_1[2727:2720]} - {1'b0, layer_0_1[2727:2720]};
      top_1[1] = {1'b0,layer_1_1[2735:2728]} - {1'b0, layer_0_1[2735:2728]};
      top_1[2] = {1'b0,layer_1_1[2743:2736]} - {1'b0, layer_0_1[2743:2736]};
      top_2[0] = {1'b0,layer_1_2[2727:2720]} - {1'b0, layer_0_2[2727:2720]};
      top_2[1] = {1'b0,layer_1_2[2735:2728]} - {1'b0, layer_0_2[2735:2728]};
      top_2[2] = {1'b0,layer_1_2[2743:2736]} - {1'b0, layer_0_2[2743:2736]};
      mid_0[0] = {1'b0,layer_2_0[2727:2720]} - {1'b0, layer_1_0[2727:2720]};
      mid_0[1] = {1'b0,layer_2_0[2735:2728]} - {1'b0, layer_1_0[2735:2728]};
      mid_0[2] = {1'b0,layer_2_0[2743:2736]} - {1'b0, layer_1_0[2743:2736]};
      mid_1[0] = {1'b0,layer_2_1[2727:2720]} - {1'b0, layer_1_1[2727:2720]};
      mid_1[1] = {1'b0,layer_2_1[2735:2728]} - {1'b0, layer_1_1[2735:2728]};
      mid_1[2] = {1'b0,layer_2_1[2743:2736]} - {1'b0, layer_1_1[2743:2736]};
      mid_2[0] = {1'b0,layer_2_2[2727:2720]} - {1'b0, layer_1_2[2727:2720]};
      mid_2[1] = {1'b0,layer_2_2[2735:2728]} - {1'b0, layer_1_2[2735:2728]};
      mid_2[2] = {1'b0,layer_2_2[2743:2736]} - {1'b0, layer_1_2[2743:2736]};
      btm_0[0] = {1'b0,layer_3_0[2727:2720]} - {1'b0, layer_2_0[2727:2720]};
      btm_0[1] = {1'b0,layer_3_0[2735:2728]} - {1'b0, layer_2_0[2735:2728]};
      btm_0[2] = {1'b0,layer_3_0[2743:2736]} - {1'b0, layer_2_0[2743:2736]};
      btm_1[0] = {1'b0,layer_3_1[2727:2720]} - {1'b0, layer_2_1[2727:2720]};
      btm_1[1] = {1'b0,layer_3_1[2735:2728]} - {1'b0, layer_2_1[2735:2728]};
      btm_1[2] = {1'b0,layer_3_1[2743:2736]} - {1'b0, layer_2_1[2743:2736]};
      btm_2[0] = {1'b0,layer_3_2[2727:2720]} - {1'b0, layer_2_2[2727:2720]};
      btm_2[1] = {1'b0,layer_3_2[2735:2728]} - {1'b0, layer_2_2[2735:2728]};
      btm_2[2] = {1'b0,layer_3_2[2743:2736]} - {1'b0, layer_2_2[2743:2736]};
    end
    'd342: begin
      top_0[0] = {1'b0,layer_1_0[2735:2728]} - {1'b0, layer_0_0[2735:2728]};
      top_0[1] = {1'b0,layer_1_0[2743:2736]} - {1'b0, layer_0_0[2743:2736]};
      top_0[2] = {1'b0,layer_1_0[2751:2744]} - {1'b0, layer_0_0[2751:2744]};
      top_1[0] = {1'b0,layer_1_1[2735:2728]} - {1'b0, layer_0_1[2735:2728]};
      top_1[1] = {1'b0,layer_1_1[2743:2736]} - {1'b0, layer_0_1[2743:2736]};
      top_1[2] = {1'b0,layer_1_1[2751:2744]} - {1'b0, layer_0_1[2751:2744]};
      top_2[0] = {1'b0,layer_1_2[2735:2728]} - {1'b0, layer_0_2[2735:2728]};
      top_2[1] = {1'b0,layer_1_2[2743:2736]} - {1'b0, layer_0_2[2743:2736]};
      top_2[2] = {1'b0,layer_1_2[2751:2744]} - {1'b0, layer_0_2[2751:2744]};
      mid_0[0] = {1'b0,layer_2_0[2735:2728]} - {1'b0, layer_1_0[2735:2728]};
      mid_0[1] = {1'b0,layer_2_0[2743:2736]} - {1'b0, layer_1_0[2743:2736]};
      mid_0[2] = {1'b0,layer_2_0[2751:2744]} - {1'b0, layer_1_0[2751:2744]};
      mid_1[0] = {1'b0,layer_2_1[2735:2728]} - {1'b0, layer_1_1[2735:2728]};
      mid_1[1] = {1'b0,layer_2_1[2743:2736]} - {1'b0, layer_1_1[2743:2736]};
      mid_1[2] = {1'b0,layer_2_1[2751:2744]} - {1'b0, layer_1_1[2751:2744]};
      mid_2[0] = {1'b0,layer_2_2[2735:2728]} - {1'b0, layer_1_2[2735:2728]};
      mid_2[1] = {1'b0,layer_2_2[2743:2736]} - {1'b0, layer_1_2[2743:2736]};
      mid_2[2] = {1'b0,layer_2_2[2751:2744]} - {1'b0, layer_1_2[2751:2744]};
      btm_0[0] = {1'b0,layer_3_0[2735:2728]} - {1'b0, layer_2_0[2735:2728]};
      btm_0[1] = {1'b0,layer_3_0[2743:2736]} - {1'b0, layer_2_0[2743:2736]};
      btm_0[2] = {1'b0,layer_3_0[2751:2744]} - {1'b0, layer_2_0[2751:2744]};
      btm_1[0] = {1'b0,layer_3_1[2735:2728]} - {1'b0, layer_2_1[2735:2728]};
      btm_1[1] = {1'b0,layer_3_1[2743:2736]} - {1'b0, layer_2_1[2743:2736]};
      btm_1[2] = {1'b0,layer_3_1[2751:2744]} - {1'b0, layer_2_1[2751:2744]};
      btm_2[0] = {1'b0,layer_3_2[2735:2728]} - {1'b0, layer_2_2[2735:2728]};
      btm_2[1] = {1'b0,layer_3_2[2743:2736]} - {1'b0, layer_2_2[2743:2736]};
      btm_2[2] = {1'b0,layer_3_2[2751:2744]} - {1'b0, layer_2_2[2751:2744]};
    end
    'd343: begin
      top_0[0] = {1'b0,layer_1_0[2743:2736]} - {1'b0, layer_0_0[2743:2736]};
      top_0[1] = {1'b0,layer_1_0[2751:2744]} - {1'b0, layer_0_0[2751:2744]};
      top_0[2] = {1'b0,layer_1_0[2759:2752]} - {1'b0, layer_0_0[2759:2752]};
      top_1[0] = {1'b0,layer_1_1[2743:2736]} - {1'b0, layer_0_1[2743:2736]};
      top_1[1] = {1'b0,layer_1_1[2751:2744]} - {1'b0, layer_0_1[2751:2744]};
      top_1[2] = {1'b0,layer_1_1[2759:2752]} - {1'b0, layer_0_1[2759:2752]};
      top_2[0] = {1'b0,layer_1_2[2743:2736]} - {1'b0, layer_0_2[2743:2736]};
      top_2[1] = {1'b0,layer_1_2[2751:2744]} - {1'b0, layer_0_2[2751:2744]};
      top_2[2] = {1'b0,layer_1_2[2759:2752]} - {1'b0, layer_0_2[2759:2752]};
      mid_0[0] = {1'b0,layer_2_0[2743:2736]} - {1'b0, layer_1_0[2743:2736]};
      mid_0[1] = {1'b0,layer_2_0[2751:2744]} - {1'b0, layer_1_0[2751:2744]};
      mid_0[2] = {1'b0,layer_2_0[2759:2752]} - {1'b0, layer_1_0[2759:2752]};
      mid_1[0] = {1'b0,layer_2_1[2743:2736]} - {1'b0, layer_1_1[2743:2736]};
      mid_1[1] = {1'b0,layer_2_1[2751:2744]} - {1'b0, layer_1_1[2751:2744]};
      mid_1[2] = {1'b0,layer_2_1[2759:2752]} - {1'b0, layer_1_1[2759:2752]};
      mid_2[0] = {1'b0,layer_2_2[2743:2736]} - {1'b0, layer_1_2[2743:2736]};
      mid_2[1] = {1'b0,layer_2_2[2751:2744]} - {1'b0, layer_1_2[2751:2744]};
      mid_2[2] = {1'b0,layer_2_2[2759:2752]} - {1'b0, layer_1_2[2759:2752]};
      btm_0[0] = {1'b0,layer_3_0[2743:2736]} - {1'b0, layer_2_0[2743:2736]};
      btm_0[1] = {1'b0,layer_3_0[2751:2744]} - {1'b0, layer_2_0[2751:2744]};
      btm_0[2] = {1'b0,layer_3_0[2759:2752]} - {1'b0, layer_2_0[2759:2752]};
      btm_1[0] = {1'b0,layer_3_1[2743:2736]} - {1'b0, layer_2_1[2743:2736]};
      btm_1[1] = {1'b0,layer_3_1[2751:2744]} - {1'b0, layer_2_1[2751:2744]};
      btm_1[2] = {1'b0,layer_3_1[2759:2752]} - {1'b0, layer_2_1[2759:2752]};
      btm_2[0] = {1'b0,layer_3_2[2743:2736]} - {1'b0, layer_2_2[2743:2736]};
      btm_2[1] = {1'b0,layer_3_2[2751:2744]} - {1'b0, layer_2_2[2751:2744]};
      btm_2[2] = {1'b0,layer_3_2[2759:2752]} - {1'b0, layer_2_2[2759:2752]};
    end
    'd344: begin
      top_0[0] = {1'b0,layer_1_0[2751:2744]} - {1'b0, layer_0_0[2751:2744]};
      top_0[1] = {1'b0,layer_1_0[2759:2752]} - {1'b0, layer_0_0[2759:2752]};
      top_0[2] = {1'b0,layer_1_0[2767:2760]} - {1'b0, layer_0_0[2767:2760]};
      top_1[0] = {1'b0,layer_1_1[2751:2744]} - {1'b0, layer_0_1[2751:2744]};
      top_1[1] = {1'b0,layer_1_1[2759:2752]} - {1'b0, layer_0_1[2759:2752]};
      top_1[2] = {1'b0,layer_1_1[2767:2760]} - {1'b0, layer_0_1[2767:2760]};
      top_2[0] = {1'b0,layer_1_2[2751:2744]} - {1'b0, layer_0_2[2751:2744]};
      top_2[1] = {1'b0,layer_1_2[2759:2752]} - {1'b0, layer_0_2[2759:2752]};
      top_2[2] = {1'b0,layer_1_2[2767:2760]} - {1'b0, layer_0_2[2767:2760]};
      mid_0[0] = {1'b0,layer_2_0[2751:2744]} - {1'b0, layer_1_0[2751:2744]};
      mid_0[1] = {1'b0,layer_2_0[2759:2752]} - {1'b0, layer_1_0[2759:2752]};
      mid_0[2] = {1'b0,layer_2_0[2767:2760]} - {1'b0, layer_1_0[2767:2760]};
      mid_1[0] = {1'b0,layer_2_1[2751:2744]} - {1'b0, layer_1_1[2751:2744]};
      mid_1[1] = {1'b0,layer_2_1[2759:2752]} - {1'b0, layer_1_1[2759:2752]};
      mid_1[2] = {1'b0,layer_2_1[2767:2760]} - {1'b0, layer_1_1[2767:2760]};
      mid_2[0] = {1'b0,layer_2_2[2751:2744]} - {1'b0, layer_1_2[2751:2744]};
      mid_2[1] = {1'b0,layer_2_2[2759:2752]} - {1'b0, layer_1_2[2759:2752]};
      mid_2[2] = {1'b0,layer_2_2[2767:2760]} - {1'b0, layer_1_2[2767:2760]};
      btm_0[0] = {1'b0,layer_3_0[2751:2744]} - {1'b0, layer_2_0[2751:2744]};
      btm_0[1] = {1'b0,layer_3_0[2759:2752]} - {1'b0, layer_2_0[2759:2752]};
      btm_0[2] = {1'b0,layer_3_0[2767:2760]} - {1'b0, layer_2_0[2767:2760]};
      btm_1[0] = {1'b0,layer_3_1[2751:2744]} - {1'b0, layer_2_1[2751:2744]};
      btm_1[1] = {1'b0,layer_3_1[2759:2752]} - {1'b0, layer_2_1[2759:2752]};
      btm_1[2] = {1'b0,layer_3_1[2767:2760]} - {1'b0, layer_2_1[2767:2760]};
      btm_2[0] = {1'b0,layer_3_2[2751:2744]} - {1'b0, layer_2_2[2751:2744]};
      btm_2[1] = {1'b0,layer_3_2[2759:2752]} - {1'b0, layer_2_2[2759:2752]};
      btm_2[2] = {1'b0,layer_3_2[2767:2760]} - {1'b0, layer_2_2[2767:2760]};
    end
    'd345: begin
      top_0[0] = {1'b0,layer_1_0[2759:2752]} - {1'b0, layer_0_0[2759:2752]};
      top_0[1] = {1'b0,layer_1_0[2767:2760]} - {1'b0, layer_0_0[2767:2760]};
      top_0[2] = {1'b0,layer_1_0[2775:2768]} - {1'b0, layer_0_0[2775:2768]};
      top_1[0] = {1'b0,layer_1_1[2759:2752]} - {1'b0, layer_0_1[2759:2752]};
      top_1[1] = {1'b0,layer_1_1[2767:2760]} - {1'b0, layer_0_1[2767:2760]};
      top_1[2] = {1'b0,layer_1_1[2775:2768]} - {1'b0, layer_0_1[2775:2768]};
      top_2[0] = {1'b0,layer_1_2[2759:2752]} - {1'b0, layer_0_2[2759:2752]};
      top_2[1] = {1'b0,layer_1_2[2767:2760]} - {1'b0, layer_0_2[2767:2760]};
      top_2[2] = {1'b0,layer_1_2[2775:2768]} - {1'b0, layer_0_2[2775:2768]};
      mid_0[0] = {1'b0,layer_2_0[2759:2752]} - {1'b0, layer_1_0[2759:2752]};
      mid_0[1] = {1'b0,layer_2_0[2767:2760]} - {1'b0, layer_1_0[2767:2760]};
      mid_0[2] = {1'b0,layer_2_0[2775:2768]} - {1'b0, layer_1_0[2775:2768]};
      mid_1[0] = {1'b0,layer_2_1[2759:2752]} - {1'b0, layer_1_1[2759:2752]};
      mid_1[1] = {1'b0,layer_2_1[2767:2760]} - {1'b0, layer_1_1[2767:2760]};
      mid_1[2] = {1'b0,layer_2_1[2775:2768]} - {1'b0, layer_1_1[2775:2768]};
      mid_2[0] = {1'b0,layer_2_2[2759:2752]} - {1'b0, layer_1_2[2759:2752]};
      mid_2[1] = {1'b0,layer_2_2[2767:2760]} - {1'b0, layer_1_2[2767:2760]};
      mid_2[2] = {1'b0,layer_2_2[2775:2768]} - {1'b0, layer_1_2[2775:2768]};
      btm_0[0] = {1'b0,layer_3_0[2759:2752]} - {1'b0, layer_2_0[2759:2752]};
      btm_0[1] = {1'b0,layer_3_0[2767:2760]} - {1'b0, layer_2_0[2767:2760]};
      btm_0[2] = {1'b0,layer_3_0[2775:2768]} - {1'b0, layer_2_0[2775:2768]};
      btm_1[0] = {1'b0,layer_3_1[2759:2752]} - {1'b0, layer_2_1[2759:2752]};
      btm_1[1] = {1'b0,layer_3_1[2767:2760]} - {1'b0, layer_2_1[2767:2760]};
      btm_1[2] = {1'b0,layer_3_1[2775:2768]} - {1'b0, layer_2_1[2775:2768]};
      btm_2[0] = {1'b0,layer_3_2[2759:2752]} - {1'b0, layer_2_2[2759:2752]};
      btm_2[1] = {1'b0,layer_3_2[2767:2760]} - {1'b0, layer_2_2[2767:2760]};
      btm_2[2] = {1'b0,layer_3_2[2775:2768]} - {1'b0, layer_2_2[2775:2768]};
    end
    'd346: begin
      top_0[0] = {1'b0,layer_1_0[2767:2760]} - {1'b0, layer_0_0[2767:2760]};
      top_0[1] = {1'b0,layer_1_0[2775:2768]} - {1'b0, layer_0_0[2775:2768]};
      top_0[2] = {1'b0,layer_1_0[2783:2776]} - {1'b0, layer_0_0[2783:2776]};
      top_1[0] = {1'b0,layer_1_1[2767:2760]} - {1'b0, layer_0_1[2767:2760]};
      top_1[1] = {1'b0,layer_1_1[2775:2768]} - {1'b0, layer_0_1[2775:2768]};
      top_1[2] = {1'b0,layer_1_1[2783:2776]} - {1'b0, layer_0_1[2783:2776]};
      top_2[0] = {1'b0,layer_1_2[2767:2760]} - {1'b0, layer_0_2[2767:2760]};
      top_2[1] = {1'b0,layer_1_2[2775:2768]} - {1'b0, layer_0_2[2775:2768]};
      top_2[2] = {1'b0,layer_1_2[2783:2776]} - {1'b0, layer_0_2[2783:2776]};
      mid_0[0] = {1'b0,layer_2_0[2767:2760]} - {1'b0, layer_1_0[2767:2760]};
      mid_0[1] = {1'b0,layer_2_0[2775:2768]} - {1'b0, layer_1_0[2775:2768]};
      mid_0[2] = {1'b0,layer_2_0[2783:2776]} - {1'b0, layer_1_0[2783:2776]};
      mid_1[0] = {1'b0,layer_2_1[2767:2760]} - {1'b0, layer_1_1[2767:2760]};
      mid_1[1] = {1'b0,layer_2_1[2775:2768]} - {1'b0, layer_1_1[2775:2768]};
      mid_1[2] = {1'b0,layer_2_1[2783:2776]} - {1'b0, layer_1_1[2783:2776]};
      mid_2[0] = {1'b0,layer_2_2[2767:2760]} - {1'b0, layer_1_2[2767:2760]};
      mid_2[1] = {1'b0,layer_2_2[2775:2768]} - {1'b0, layer_1_2[2775:2768]};
      mid_2[2] = {1'b0,layer_2_2[2783:2776]} - {1'b0, layer_1_2[2783:2776]};
      btm_0[0] = {1'b0,layer_3_0[2767:2760]} - {1'b0, layer_2_0[2767:2760]};
      btm_0[1] = {1'b0,layer_3_0[2775:2768]} - {1'b0, layer_2_0[2775:2768]};
      btm_0[2] = {1'b0,layer_3_0[2783:2776]} - {1'b0, layer_2_0[2783:2776]};
      btm_1[0] = {1'b0,layer_3_1[2767:2760]} - {1'b0, layer_2_1[2767:2760]};
      btm_1[1] = {1'b0,layer_3_1[2775:2768]} - {1'b0, layer_2_1[2775:2768]};
      btm_1[2] = {1'b0,layer_3_1[2783:2776]} - {1'b0, layer_2_1[2783:2776]};
      btm_2[0] = {1'b0,layer_3_2[2767:2760]} - {1'b0, layer_2_2[2767:2760]};
      btm_2[1] = {1'b0,layer_3_2[2775:2768]} - {1'b0, layer_2_2[2775:2768]};
      btm_2[2] = {1'b0,layer_3_2[2783:2776]} - {1'b0, layer_2_2[2783:2776]};
    end
    'd347: begin
      top_0[0] = {1'b0,layer_1_0[2775:2768]} - {1'b0, layer_0_0[2775:2768]};
      top_0[1] = {1'b0,layer_1_0[2783:2776]} - {1'b0, layer_0_0[2783:2776]};
      top_0[2] = {1'b0,layer_1_0[2791:2784]} - {1'b0, layer_0_0[2791:2784]};
      top_1[0] = {1'b0,layer_1_1[2775:2768]} - {1'b0, layer_0_1[2775:2768]};
      top_1[1] = {1'b0,layer_1_1[2783:2776]} - {1'b0, layer_0_1[2783:2776]};
      top_1[2] = {1'b0,layer_1_1[2791:2784]} - {1'b0, layer_0_1[2791:2784]};
      top_2[0] = {1'b0,layer_1_2[2775:2768]} - {1'b0, layer_0_2[2775:2768]};
      top_2[1] = {1'b0,layer_1_2[2783:2776]} - {1'b0, layer_0_2[2783:2776]};
      top_2[2] = {1'b0,layer_1_2[2791:2784]} - {1'b0, layer_0_2[2791:2784]};
      mid_0[0] = {1'b0,layer_2_0[2775:2768]} - {1'b0, layer_1_0[2775:2768]};
      mid_0[1] = {1'b0,layer_2_0[2783:2776]} - {1'b0, layer_1_0[2783:2776]};
      mid_0[2] = {1'b0,layer_2_0[2791:2784]} - {1'b0, layer_1_0[2791:2784]};
      mid_1[0] = {1'b0,layer_2_1[2775:2768]} - {1'b0, layer_1_1[2775:2768]};
      mid_1[1] = {1'b0,layer_2_1[2783:2776]} - {1'b0, layer_1_1[2783:2776]};
      mid_1[2] = {1'b0,layer_2_1[2791:2784]} - {1'b0, layer_1_1[2791:2784]};
      mid_2[0] = {1'b0,layer_2_2[2775:2768]} - {1'b0, layer_1_2[2775:2768]};
      mid_2[1] = {1'b0,layer_2_2[2783:2776]} - {1'b0, layer_1_2[2783:2776]};
      mid_2[2] = {1'b0,layer_2_2[2791:2784]} - {1'b0, layer_1_2[2791:2784]};
      btm_0[0] = {1'b0,layer_3_0[2775:2768]} - {1'b0, layer_2_0[2775:2768]};
      btm_0[1] = {1'b0,layer_3_0[2783:2776]} - {1'b0, layer_2_0[2783:2776]};
      btm_0[2] = {1'b0,layer_3_0[2791:2784]} - {1'b0, layer_2_0[2791:2784]};
      btm_1[0] = {1'b0,layer_3_1[2775:2768]} - {1'b0, layer_2_1[2775:2768]};
      btm_1[1] = {1'b0,layer_3_1[2783:2776]} - {1'b0, layer_2_1[2783:2776]};
      btm_1[2] = {1'b0,layer_3_1[2791:2784]} - {1'b0, layer_2_1[2791:2784]};
      btm_2[0] = {1'b0,layer_3_2[2775:2768]} - {1'b0, layer_2_2[2775:2768]};
      btm_2[1] = {1'b0,layer_3_2[2783:2776]} - {1'b0, layer_2_2[2783:2776]};
      btm_2[2] = {1'b0,layer_3_2[2791:2784]} - {1'b0, layer_2_2[2791:2784]};
    end
    'd348: begin
      top_0[0] = {1'b0,layer_1_0[2783:2776]} - {1'b0, layer_0_0[2783:2776]};
      top_0[1] = {1'b0,layer_1_0[2791:2784]} - {1'b0, layer_0_0[2791:2784]};
      top_0[2] = {1'b0,layer_1_0[2799:2792]} - {1'b0, layer_0_0[2799:2792]};
      top_1[0] = {1'b0,layer_1_1[2783:2776]} - {1'b0, layer_0_1[2783:2776]};
      top_1[1] = {1'b0,layer_1_1[2791:2784]} - {1'b0, layer_0_1[2791:2784]};
      top_1[2] = {1'b0,layer_1_1[2799:2792]} - {1'b0, layer_0_1[2799:2792]};
      top_2[0] = {1'b0,layer_1_2[2783:2776]} - {1'b0, layer_0_2[2783:2776]};
      top_2[1] = {1'b0,layer_1_2[2791:2784]} - {1'b0, layer_0_2[2791:2784]};
      top_2[2] = {1'b0,layer_1_2[2799:2792]} - {1'b0, layer_0_2[2799:2792]};
      mid_0[0] = {1'b0,layer_2_0[2783:2776]} - {1'b0, layer_1_0[2783:2776]};
      mid_0[1] = {1'b0,layer_2_0[2791:2784]} - {1'b0, layer_1_0[2791:2784]};
      mid_0[2] = {1'b0,layer_2_0[2799:2792]} - {1'b0, layer_1_0[2799:2792]};
      mid_1[0] = {1'b0,layer_2_1[2783:2776]} - {1'b0, layer_1_1[2783:2776]};
      mid_1[1] = {1'b0,layer_2_1[2791:2784]} - {1'b0, layer_1_1[2791:2784]};
      mid_1[2] = {1'b0,layer_2_1[2799:2792]} - {1'b0, layer_1_1[2799:2792]};
      mid_2[0] = {1'b0,layer_2_2[2783:2776]} - {1'b0, layer_1_2[2783:2776]};
      mid_2[1] = {1'b0,layer_2_2[2791:2784]} - {1'b0, layer_1_2[2791:2784]};
      mid_2[2] = {1'b0,layer_2_2[2799:2792]} - {1'b0, layer_1_2[2799:2792]};
      btm_0[0] = {1'b0,layer_3_0[2783:2776]} - {1'b0, layer_2_0[2783:2776]};
      btm_0[1] = {1'b0,layer_3_0[2791:2784]} - {1'b0, layer_2_0[2791:2784]};
      btm_0[2] = {1'b0,layer_3_0[2799:2792]} - {1'b0, layer_2_0[2799:2792]};
      btm_1[0] = {1'b0,layer_3_1[2783:2776]} - {1'b0, layer_2_1[2783:2776]};
      btm_1[1] = {1'b0,layer_3_1[2791:2784]} - {1'b0, layer_2_1[2791:2784]};
      btm_1[2] = {1'b0,layer_3_1[2799:2792]} - {1'b0, layer_2_1[2799:2792]};
      btm_2[0] = {1'b0,layer_3_2[2783:2776]} - {1'b0, layer_2_2[2783:2776]};
      btm_2[1] = {1'b0,layer_3_2[2791:2784]} - {1'b0, layer_2_2[2791:2784]};
      btm_2[2] = {1'b0,layer_3_2[2799:2792]} - {1'b0, layer_2_2[2799:2792]};
    end
    'd349: begin
      top_0[0] = {1'b0,layer_1_0[2791:2784]} - {1'b0, layer_0_0[2791:2784]};
      top_0[1] = {1'b0,layer_1_0[2799:2792]} - {1'b0, layer_0_0[2799:2792]};
      top_0[2] = {1'b0,layer_1_0[2807:2800]} - {1'b0, layer_0_0[2807:2800]};
      top_1[0] = {1'b0,layer_1_1[2791:2784]} - {1'b0, layer_0_1[2791:2784]};
      top_1[1] = {1'b0,layer_1_1[2799:2792]} - {1'b0, layer_0_1[2799:2792]};
      top_1[2] = {1'b0,layer_1_1[2807:2800]} - {1'b0, layer_0_1[2807:2800]};
      top_2[0] = {1'b0,layer_1_2[2791:2784]} - {1'b0, layer_0_2[2791:2784]};
      top_2[1] = {1'b0,layer_1_2[2799:2792]} - {1'b0, layer_0_2[2799:2792]};
      top_2[2] = {1'b0,layer_1_2[2807:2800]} - {1'b0, layer_0_2[2807:2800]};
      mid_0[0] = {1'b0,layer_2_0[2791:2784]} - {1'b0, layer_1_0[2791:2784]};
      mid_0[1] = {1'b0,layer_2_0[2799:2792]} - {1'b0, layer_1_0[2799:2792]};
      mid_0[2] = {1'b0,layer_2_0[2807:2800]} - {1'b0, layer_1_0[2807:2800]};
      mid_1[0] = {1'b0,layer_2_1[2791:2784]} - {1'b0, layer_1_1[2791:2784]};
      mid_1[1] = {1'b0,layer_2_1[2799:2792]} - {1'b0, layer_1_1[2799:2792]};
      mid_1[2] = {1'b0,layer_2_1[2807:2800]} - {1'b0, layer_1_1[2807:2800]};
      mid_2[0] = {1'b0,layer_2_2[2791:2784]} - {1'b0, layer_1_2[2791:2784]};
      mid_2[1] = {1'b0,layer_2_2[2799:2792]} - {1'b0, layer_1_2[2799:2792]};
      mid_2[2] = {1'b0,layer_2_2[2807:2800]} - {1'b0, layer_1_2[2807:2800]};
      btm_0[0] = {1'b0,layer_3_0[2791:2784]} - {1'b0, layer_2_0[2791:2784]};
      btm_0[1] = {1'b0,layer_3_0[2799:2792]} - {1'b0, layer_2_0[2799:2792]};
      btm_0[2] = {1'b0,layer_3_0[2807:2800]} - {1'b0, layer_2_0[2807:2800]};
      btm_1[0] = {1'b0,layer_3_1[2791:2784]} - {1'b0, layer_2_1[2791:2784]};
      btm_1[1] = {1'b0,layer_3_1[2799:2792]} - {1'b0, layer_2_1[2799:2792]};
      btm_1[2] = {1'b0,layer_3_1[2807:2800]} - {1'b0, layer_2_1[2807:2800]};
      btm_2[0] = {1'b0,layer_3_2[2791:2784]} - {1'b0, layer_2_2[2791:2784]};
      btm_2[1] = {1'b0,layer_3_2[2799:2792]} - {1'b0, layer_2_2[2799:2792]};
      btm_2[2] = {1'b0,layer_3_2[2807:2800]} - {1'b0, layer_2_2[2807:2800]};
    end
    'd350: begin
      top_0[0] = {1'b0,layer_1_0[2799:2792]} - {1'b0, layer_0_0[2799:2792]};
      top_0[1] = {1'b0,layer_1_0[2807:2800]} - {1'b0, layer_0_0[2807:2800]};
      top_0[2] = {1'b0,layer_1_0[2815:2808]} - {1'b0, layer_0_0[2815:2808]};
      top_1[0] = {1'b0,layer_1_1[2799:2792]} - {1'b0, layer_0_1[2799:2792]};
      top_1[1] = {1'b0,layer_1_1[2807:2800]} - {1'b0, layer_0_1[2807:2800]};
      top_1[2] = {1'b0,layer_1_1[2815:2808]} - {1'b0, layer_0_1[2815:2808]};
      top_2[0] = {1'b0,layer_1_2[2799:2792]} - {1'b0, layer_0_2[2799:2792]};
      top_2[1] = {1'b0,layer_1_2[2807:2800]} - {1'b0, layer_0_2[2807:2800]};
      top_2[2] = {1'b0,layer_1_2[2815:2808]} - {1'b0, layer_0_2[2815:2808]};
      mid_0[0] = {1'b0,layer_2_0[2799:2792]} - {1'b0, layer_1_0[2799:2792]};
      mid_0[1] = {1'b0,layer_2_0[2807:2800]} - {1'b0, layer_1_0[2807:2800]};
      mid_0[2] = {1'b0,layer_2_0[2815:2808]} - {1'b0, layer_1_0[2815:2808]};
      mid_1[0] = {1'b0,layer_2_1[2799:2792]} - {1'b0, layer_1_1[2799:2792]};
      mid_1[1] = {1'b0,layer_2_1[2807:2800]} - {1'b0, layer_1_1[2807:2800]};
      mid_1[2] = {1'b0,layer_2_1[2815:2808]} - {1'b0, layer_1_1[2815:2808]};
      mid_2[0] = {1'b0,layer_2_2[2799:2792]} - {1'b0, layer_1_2[2799:2792]};
      mid_2[1] = {1'b0,layer_2_2[2807:2800]} - {1'b0, layer_1_2[2807:2800]};
      mid_2[2] = {1'b0,layer_2_2[2815:2808]} - {1'b0, layer_1_2[2815:2808]};
      btm_0[0] = {1'b0,layer_3_0[2799:2792]} - {1'b0, layer_2_0[2799:2792]};
      btm_0[1] = {1'b0,layer_3_0[2807:2800]} - {1'b0, layer_2_0[2807:2800]};
      btm_0[2] = {1'b0,layer_3_0[2815:2808]} - {1'b0, layer_2_0[2815:2808]};
      btm_1[0] = {1'b0,layer_3_1[2799:2792]} - {1'b0, layer_2_1[2799:2792]};
      btm_1[1] = {1'b0,layer_3_1[2807:2800]} - {1'b0, layer_2_1[2807:2800]};
      btm_1[2] = {1'b0,layer_3_1[2815:2808]} - {1'b0, layer_2_1[2815:2808]};
      btm_2[0] = {1'b0,layer_3_2[2799:2792]} - {1'b0, layer_2_2[2799:2792]};
      btm_2[1] = {1'b0,layer_3_2[2807:2800]} - {1'b0, layer_2_2[2807:2800]};
      btm_2[2] = {1'b0,layer_3_2[2815:2808]} - {1'b0, layer_2_2[2815:2808]};
    end
    'd351: begin
      top_0[0] = {1'b0,layer_1_0[2807:2800]} - {1'b0, layer_0_0[2807:2800]};
      top_0[1] = {1'b0,layer_1_0[2815:2808]} - {1'b0, layer_0_0[2815:2808]};
      top_0[2] = {1'b0,layer_1_0[2823:2816]} - {1'b0, layer_0_0[2823:2816]};
      top_1[0] = {1'b0,layer_1_1[2807:2800]} - {1'b0, layer_0_1[2807:2800]};
      top_1[1] = {1'b0,layer_1_1[2815:2808]} - {1'b0, layer_0_1[2815:2808]};
      top_1[2] = {1'b0,layer_1_1[2823:2816]} - {1'b0, layer_0_1[2823:2816]};
      top_2[0] = {1'b0,layer_1_2[2807:2800]} - {1'b0, layer_0_2[2807:2800]};
      top_2[1] = {1'b0,layer_1_2[2815:2808]} - {1'b0, layer_0_2[2815:2808]};
      top_2[2] = {1'b0,layer_1_2[2823:2816]} - {1'b0, layer_0_2[2823:2816]};
      mid_0[0] = {1'b0,layer_2_0[2807:2800]} - {1'b0, layer_1_0[2807:2800]};
      mid_0[1] = {1'b0,layer_2_0[2815:2808]} - {1'b0, layer_1_0[2815:2808]};
      mid_0[2] = {1'b0,layer_2_0[2823:2816]} - {1'b0, layer_1_0[2823:2816]};
      mid_1[0] = {1'b0,layer_2_1[2807:2800]} - {1'b0, layer_1_1[2807:2800]};
      mid_1[1] = {1'b0,layer_2_1[2815:2808]} - {1'b0, layer_1_1[2815:2808]};
      mid_1[2] = {1'b0,layer_2_1[2823:2816]} - {1'b0, layer_1_1[2823:2816]};
      mid_2[0] = {1'b0,layer_2_2[2807:2800]} - {1'b0, layer_1_2[2807:2800]};
      mid_2[1] = {1'b0,layer_2_2[2815:2808]} - {1'b0, layer_1_2[2815:2808]};
      mid_2[2] = {1'b0,layer_2_2[2823:2816]} - {1'b0, layer_1_2[2823:2816]};
      btm_0[0] = {1'b0,layer_3_0[2807:2800]} - {1'b0, layer_2_0[2807:2800]};
      btm_0[1] = {1'b0,layer_3_0[2815:2808]} - {1'b0, layer_2_0[2815:2808]};
      btm_0[2] = {1'b0,layer_3_0[2823:2816]} - {1'b0, layer_2_0[2823:2816]};
      btm_1[0] = {1'b0,layer_3_1[2807:2800]} - {1'b0, layer_2_1[2807:2800]};
      btm_1[1] = {1'b0,layer_3_1[2815:2808]} - {1'b0, layer_2_1[2815:2808]};
      btm_1[2] = {1'b0,layer_3_1[2823:2816]} - {1'b0, layer_2_1[2823:2816]};
      btm_2[0] = {1'b0,layer_3_2[2807:2800]} - {1'b0, layer_2_2[2807:2800]};
      btm_2[1] = {1'b0,layer_3_2[2815:2808]} - {1'b0, layer_2_2[2815:2808]};
      btm_2[2] = {1'b0,layer_3_2[2823:2816]} - {1'b0, layer_2_2[2823:2816]};
    end
    'd352: begin
      top_0[0] = {1'b0,layer_1_0[2815:2808]} - {1'b0, layer_0_0[2815:2808]};
      top_0[1] = {1'b0,layer_1_0[2823:2816]} - {1'b0, layer_0_0[2823:2816]};
      top_0[2] = {1'b0,layer_1_0[2831:2824]} - {1'b0, layer_0_0[2831:2824]};
      top_1[0] = {1'b0,layer_1_1[2815:2808]} - {1'b0, layer_0_1[2815:2808]};
      top_1[1] = {1'b0,layer_1_1[2823:2816]} - {1'b0, layer_0_1[2823:2816]};
      top_1[2] = {1'b0,layer_1_1[2831:2824]} - {1'b0, layer_0_1[2831:2824]};
      top_2[0] = {1'b0,layer_1_2[2815:2808]} - {1'b0, layer_0_2[2815:2808]};
      top_2[1] = {1'b0,layer_1_2[2823:2816]} - {1'b0, layer_0_2[2823:2816]};
      top_2[2] = {1'b0,layer_1_2[2831:2824]} - {1'b0, layer_0_2[2831:2824]};
      mid_0[0] = {1'b0,layer_2_0[2815:2808]} - {1'b0, layer_1_0[2815:2808]};
      mid_0[1] = {1'b0,layer_2_0[2823:2816]} - {1'b0, layer_1_0[2823:2816]};
      mid_0[2] = {1'b0,layer_2_0[2831:2824]} - {1'b0, layer_1_0[2831:2824]};
      mid_1[0] = {1'b0,layer_2_1[2815:2808]} - {1'b0, layer_1_1[2815:2808]};
      mid_1[1] = {1'b0,layer_2_1[2823:2816]} - {1'b0, layer_1_1[2823:2816]};
      mid_1[2] = {1'b0,layer_2_1[2831:2824]} - {1'b0, layer_1_1[2831:2824]};
      mid_2[0] = {1'b0,layer_2_2[2815:2808]} - {1'b0, layer_1_2[2815:2808]};
      mid_2[1] = {1'b0,layer_2_2[2823:2816]} - {1'b0, layer_1_2[2823:2816]};
      mid_2[2] = {1'b0,layer_2_2[2831:2824]} - {1'b0, layer_1_2[2831:2824]};
      btm_0[0] = {1'b0,layer_3_0[2815:2808]} - {1'b0, layer_2_0[2815:2808]};
      btm_0[1] = {1'b0,layer_3_0[2823:2816]} - {1'b0, layer_2_0[2823:2816]};
      btm_0[2] = {1'b0,layer_3_0[2831:2824]} - {1'b0, layer_2_0[2831:2824]};
      btm_1[0] = {1'b0,layer_3_1[2815:2808]} - {1'b0, layer_2_1[2815:2808]};
      btm_1[1] = {1'b0,layer_3_1[2823:2816]} - {1'b0, layer_2_1[2823:2816]};
      btm_1[2] = {1'b0,layer_3_1[2831:2824]} - {1'b0, layer_2_1[2831:2824]};
      btm_2[0] = {1'b0,layer_3_2[2815:2808]} - {1'b0, layer_2_2[2815:2808]};
      btm_2[1] = {1'b0,layer_3_2[2823:2816]} - {1'b0, layer_2_2[2823:2816]};
      btm_2[2] = {1'b0,layer_3_2[2831:2824]} - {1'b0, layer_2_2[2831:2824]};
    end
    'd353: begin
      top_0[0] = {1'b0,layer_1_0[2823:2816]} - {1'b0, layer_0_0[2823:2816]};
      top_0[1] = {1'b0,layer_1_0[2831:2824]} - {1'b0, layer_0_0[2831:2824]};
      top_0[2] = {1'b0,layer_1_0[2839:2832]} - {1'b0, layer_0_0[2839:2832]};
      top_1[0] = {1'b0,layer_1_1[2823:2816]} - {1'b0, layer_0_1[2823:2816]};
      top_1[1] = {1'b0,layer_1_1[2831:2824]} - {1'b0, layer_0_1[2831:2824]};
      top_1[2] = {1'b0,layer_1_1[2839:2832]} - {1'b0, layer_0_1[2839:2832]};
      top_2[0] = {1'b0,layer_1_2[2823:2816]} - {1'b0, layer_0_2[2823:2816]};
      top_2[1] = {1'b0,layer_1_2[2831:2824]} - {1'b0, layer_0_2[2831:2824]};
      top_2[2] = {1'b0,layer_1_2[2839:2832]} - {1'b0, layer_0_2[2839:2832]};
      mid_0[0] = {1'b0,layer_2_0[2823:2816]} - {1'b0, layer_1_0[2823:2816]};
      mid_0[1] = {1'b0,layer_2_0[2831:2824]} - {1'b0, layer_1_0[2831:2824]};
      mid_0[2] = {1'b0,layer_2_0[2839:2832]} - {1'b0, layer_1_0[2839:2832]};
      mid_1[0] = {1'b0,layer_2_1[2823:2816]} - {1'b0, layer_1_1[2823:2816]};
      mid_1[1] = {1'b0,layer_2_1[2831:2824]} - {1'b0, layer_1_1[2831:2824]};
      mid_1[2] = {1'b0,layer_2_1[2839:2832]} - {1'b0, layer_1_1[2839:2832]};
      mid_2[0] = {1'b0,layer_2_2[2823:2816]} - {1'b0, layer_1_2[2823:2816]};
      mid_2[1] = {1'b0,layer_2_2[2831:2824]} - {1'b0, layer_1_2[2831:2824]};
      mid_2[2] = {1'b0,layer_2_2[2839:2832]} - {1'b0, layer_1_2[2839:2832]};
      btm_0[0] = {1'b0,layer_3_0[2823:2816]} - {1'b0, layer_2_0[2823:2816]};
      btm_0[1] = {1'b0,layer_3_0[2831:2824]} - {1'b0, layer_2_0[2831:2824]};
      btm_0[2] = {1'b0,layer_3_0[2839:2832]} - {1'b0, layer_2_0[2839:2832]};
      btm_1[0] = {1'b0,layer_3_1[2823:2816]} - {1'b0, layer_2_1[2823:2816]};
      btm_1[1] = {1'b0,layer_3_1[2831:2824]} - {1'b0, layer_2_1[2831:2824]};
      btm_1[2] = {1'b0,layer_3_1[2839:2832]} - {1'b0, layer_2_1[2839:2832]};
      btm_2[0] = {1'b0,layer_3_2[2823:2816]} - {1'b0, layer_2_2[2823:2816]};
      btm_2[1] = {1'b0,layer_3_2[2831:2824]} - {1'b0, layer_2_2[2831:2824]};
      btm_2[2] = {1'b0,layer_3_2[2839:2832]} - {1'b0, layer_2_2[2839:2832]};
    end
    'd354: begin
      top_0[0] = {1'b0,layer_1_0[2831:2824]} - {1'b0, layer_0_0[2831:2824]};
      top_0[1] = {1'b0,layer_1_0[2839:2832]} - {1'b0, layer_0_0[2839:2832]};
      top_0[2] = {1'b0,layer_1_0[2847:2840]} - {1'b0, layer_0_0[2847:2840]};
      top_1[0] = {1'b0,layer_1_1[2831:2824]} - {1'b0, layer_0_1[2831:2824]};
      top_1[1] = {1'b0,layer_1_1[2839:2832]} - {1'b0, layer_0_1[2839:2832]};
      top_1[2] = {1'b0,layer_1_1[2847:2840]} - {1'b0, layer_0_1[2847:2840]};
      top_2[0] = {1'b0,layer_1_2[2831:2824]} - {1'b0, layer_0_2[2831:2824]};
      top_2[1] = {1'b0,layer_1_2[2839:2832]} - {1'b0, layer_0_2[2839:2832]};
      top_2[2] = {1'b0,layer_1_2[2847:2840]} - {1'b0, layer_0_2[2847:2840]};
      mid_0[0] = {1'b0,layer_2_0[2831:2824]} - {1'b0, layer_1_0[2831:2824]};
      mid_0[1] = {1'b0,layer_2_0[2839:2832]} - {1'b0, layer_1_0[2839:2832]};
      mid_0[2] = {1'b0,layer_2_0[2847:2840]} - {1'b0, layer_1_0[2847:2840]};
      mid_1[0] = {1'b0,layer_2_1[2831:2824]} - {1'b0, layer_1_1[2831:2824]};
      mid_1[1] = {1'b0,layer_2_1[2839:2832]} - {1'b0, layer_1_1[2839:2832]};
      mid_1[2] = {1'b0,layer_2_1[2847:2840]} - {1'b0, layer_1_1[2847:2840]};
      mid_2[0] = {1'b0,layer_2_2[2831:2824]} - {1'b0, layer_1_2[2831:2824]};
      mid_2[1] = {1'b0,layer_2_2[2839:2832]} - {1'b0, layer_1_2[2839:2832]};
      mid_2[2] = {1'b0,layer_2_2[2847:2840]} - {1'b0, layer_1_2[2847:2840]};
      btm_0[0] = {1'b0,layer_3_0[2831:2824]} - {1'b0, layer_2_0[2831:2824]};
      btm_0[1] = {1'b0,layer_3_0[2839:2832]} - {1'b0, layer_2_0[2839:2832]};
      btm_0[2] = {1'b0,layer_3_0[2847:2840]} - {1'b0, layer_2_0[2847:2840]};
      btm_1[0] = {1'b0,layer_3_1[2831:2824]} - {1'b0, layer_2_1[2831:2824]};
      btm_1[1] = {1'b0,layer_3_1[2839:2832]} - {1'b0, layer_2_1[2839:2832]};
      btm_1[2] = {1'b0,layer_3_1[2847:2840]} - {1'b0, layer_2_1[2847:2840]};
      btm_2[0] = {1'b0,layer_3_2[2831:2824]} - {1'b0, layer_2_2[2831:2824]};
      btm_2[1] = {1'b0,layer_3_2[2839:2832]} - {1'b0, layer_2_2[2839:2832]};
      btm_2[2] = {1'b0,layer_3_2[2847:2840]} - {1'b0, layer_2_2[2847:2840]};
    end
    'd355: begin
      top_0[0] = {1'b0,layer_1_0[2839:2832]} - {1'b0, layer_0_0[2839:2832]};
      top_0[1] = {1'b0,layer_1_0[2847:2840]} - {1'b0, layer_0_0[2847:2840]};
      top_0[2] = {1'b0,layer_1_0[2855:2848]} - {1'b0, layer_0_0[2855:2848]};
      top_1[0] = {1'b0,layer_1_1[2839:2832]} - {1'b0, layer_0_1[2839:2832]};
      top_1[1] = {1'b0,layer_1_1[2847:2840]} - {1'b0, layer_0_1[2847:2840]};
      top_1[2] = {1'b0,layer_1_1[2855:2848]} - {1'b0, layer_0_1[2855:2848]};
      top_2[0] = {1'b0,layer_1_2[2839:2832]} - {1'b0, layer_0_2[2839:2832]};
      top_2[1] = {1'b0,layer_1_2[2847:2840]} - {1'b0, layer_0_2[2847:2840]};
      top_2[2] = {1'b0,layer_1_2[2855:2848]} - {1'b0, layer_0_2[2855:2848]};
      mid_0[0] = {1'b0,layer_2_0[2839:2832]} - {1'b0, layer_1_0[2839:2832]};
      mid_0[1] = {1'b0,layer_2_0[2847:2840]} - {1'b0, layer_1_0[2847:2840]};
      mid_0[2] = {1'b0,layer_2_0[2855:2848]} - {1'b0, layer_1_0[2855:2848]};
      mid_1[0] = {1'b0,layer_2_1[2839:2832]} - {1'b0, layer_1_1[2839:2832]};
      mid_1[1] = {1'b0,layer_2_1[2847:2840]} - {1'b0, layer_1_1[2847:2840]};
      mid_1[2] = {1'b0,layer_2_1[2855:2848]} - {1'b0, layer_1_1[2855:2848]};
      mid_2[0] = {1'b0,layer_2_2[2839:2832]} - {1'b0, layer_1_2[2839:2832]};
      mid_2[1] = {1'b0,layer_2_2[2847:2840]} - {1'b0, layer_1_2[2847:2840]};
      mid_2[2] = {1'b0,layer_2_2[2855:2848]} - {1'b0, layer_1_2[2855:2848]};
      btm_0[0] = {1'b0,layer_3_0[2839:2832]} - {1'b0, layer_2_0[2839:2832]};
      btm_0[1] = {1'b0,layer_3_0[2847:2840]} - {1'b0, layer_2_0[2847:2840]};
      btm_0[2] = {1'b0,layer_3_0[2855:2848]} - {1'b0, layer_2_0[2855:2848]};
      btm_1[0] = {1'b0,layer_3_1[2839:2832]} - {1'b0, layer_2_1[2839:2832]};
      btm_1[1] = {1'b0,layer_3_1[2847:2840]} - {1'b0, layer_2_1[2847:2840]};
      btm_1[2] = {1'b0,layer_3_1[2855:2848]} - {1'b0, layer_2_1[2855:2848]};
      btm_2[0] = {1'b0,layer_3_2[2839:2832]} - {1'b0, layer_2_2[2839:2832]};
      btm_2[1] = {1'b0,layer_3_2[2847:2840]} - {1'b0, layer_2_2[2847:2840]};
      btm_2[2] = {1'b0,layer_3_2[2855:2848]} - {1'b0, layer_2_2[2855:2848]};
    end
    'd356: begin
      top_0[0] = {1'b0,layer_1_0[2847:2840]} - {1'b0, layer_0_0[2847:2840]};
      top_0[1] = {1'b0,layer_1_0[2855:2848]} - {1'b0, layer_0_0[2855:2848]};
      top_0[2] = {1'b0,layer_1_0[2863:2856]} - {1'b0, layer_0_0[2863:2856]};
      top_1[0] = {1'b0,layer_1_1[2847:2840]} - {1'b0, layer_0_1[2847:2840]};
      top_1[1] = {1'b0,layer_1_1[2855:2848]} - {1'b0, layer_0_1[2855:2848]};
      top_1[2] = {1'b0,layer_1_1[2863:2856]} - {1'b0, layer_0_1[2863:2856]};
      top_2[0] = {1'b0,layer_1_2[2847:2840]} - {1'b0, layer_0_2[2847:2840]};
      top_2[1] = {1'b0,layer_1_2[2855:2848]} - {1'b0, layer_0_2[2855:2848]};
      top_2[2] = {1'b0,layer_1_2[2863:2856]} - {1'b0, layer_0_2[2863:2856]};
      mid_0[0] = {1'b0,layer_2_0[2847:2840]} - {1'b0, layer_1_0[2847:2840]};
      mid_0[1] = {1'b0,layer_2_0[2855:2848]} - {1'b0, layer_1_0[2855:2848]};
      mid_0[2] = {1'b0,layer_2_0[2863:2856]} - {1'b0, layer_1_0[2863:2856]};
      mid_1[0] = {1'b0,layer_2_1[2847:2840]} - {1'b0, layer_1_1[2847:2840]};
      mid_1[1] = {1'b0,layer_2_1[2855:2848]} - {1'b0, layer_1_1[2855:2848]};
      mid_1[2] = {1'b0,layer_2_1[2863:2856]} - {1'b0, layer_1_1[2863:2856]};
      mid_2[0] = {1'b0,layer_2_2[2847:2840]} - {1'b0, layer_1_2[2847:2840]};
      mid_2[1] = {1'b0,layer_2_2[2855:2848]} - {1'b0, layer_1_2[2855:2848]};
      mid_2[2] = {1'b0,layer_2_2[2863:2856]} - {1'b0, layer_1_2[2863:2856]};
      btm_0[0] = {1'b0,layer_3_0[2847:2840]} - {1'b0, layer_2_0[2847:2840]};
      btm_0[1] = {1'b0,layer_3_0[2855:2848]} - {1'b0, layer_2_0[2855:2848]};
      btm_0[2] = {1'b0,layer_3_0[2863:2856]} - {1'b0, layer_2_0[2863:2856]};
      btm_1[0] = {1'b0,layer_3_1[2847:2840]} - {1'b0, layer_2_1[2847:2840]};
      btm_1[1] = {1'b0,layer_3_1[2855:2848]} - {1'b0, layer_2_1[2855:2848]};
      btm_1[2] = {1'b0,layer_3_1[2863:2856]} - {1'b0, layer_2_1[2863:2856]};
      btm_2[0] = {1'b0,layer_3_2[2847:2840]} - {1'b0, layer_2_2[2847:2840]};
      btm_2[1] = {1'b0,layer_3_2[2855:2848]} - {1'b0, layer_2_2[2855:2848]};
      btm_2[2] = {1'b0,layer_3_2[2863:2856]} - {1'b0, layer_2_2[2863:2856]};
    end
    'd357: begin
      top_0[0] = {1'b0,layer_1_0[2855:2848]} - {1'b0, layer_0_0[2855:2848]};
      top_0[1] = {1'b0,layer_1_0[2863:2856]} - {1'b0, layer_0_0[2863:2856]};
      top_0[2] = {1'b0,layer_1_0[2871:2864]} - {1'b0, layer_0_0[2871:2864]};
      top_1[0] = {1'b0,layer_1_1[2855:2848]} - {1'b0, layer_0_1[2855:2848]};
      top_1[1] = {1'b0,layer_1_1[2863:2856]} - {1'b0, layer_0_1[2863:2856]};
      top_1[2] = {1'b0,layer_1_1[2871:2864]} - {1'b0, layer_0_1[2871:2864]};
      top_2[0] = {1'b0,layer_1_2[2855:2848]} - {1'b0, layer_0_2[2855:2848]};
      top_2[1] = {1'b0,layer_1_2[2863:2856]} - {1'b0, layer_0_2[2863:2856]};
      top_2[2] = {1'b0,layer_1_2[2871:2864]} - {1'b0, layer_0_2[2871:2864]};
      mid_0[0] = {1'b0,layer_2_0[2855:2848]} - {1'b0, layer_1_0[2855:2848]};
      mid_0[1] = {1'b0,layer_2_0[2863:2856]} - {1'b0, layer_1_0[2863:2856]};
      mid_0[2] = {1'b0,layer_2_0[2871:2864]} - {1'b0, layer_1_0[2871:2864]};
      mid_1[0] = {1'b0,layer_2_1[2855:2848]} - {1'b0, layer_1_1[2855:2848]};
      mid_1[1] = {1'b0,layer_2_1[2863:2856]} - {1'b0, layer_1_1[2863:2856]};
      mid_1[2] = {1'b0,layer_2_1[2871:2864]} - {1'b0, layer_1_1[2871:2864]};
      mid_2[0] = {1'b0,layer_2_2[2855:2848]} - {1'b0, layer_1_2[2855:2848]};
      mid_2[1] = {1'b0,layer_2_2[2863:2856]} - {1'b0, layer_1_2[2863:2856]};
      mid_2[2] = {1'b0,layer_2_2[2871:2864]} - {1'b0, layer_1_2[2871:2864]};
      btm_0[0] = {1'b0,layer_3_0[2855:2848]} - {1'b0, layer_2_0[2855:2848]};
      btm_0[1] = {1'b0,layer_3_0[2863:2856]} - {1'b0, layer_2_0[2863:2856]};
      btm_0[2] = {1'b0,layer_3_0[2871:2864]} - {1'b0, layer_2_0[2871:2864]};
      btm_1[0] = {1'b0,layer_3_1[2855:2848]} - {1'b0, layer_2_1[2855:2848]};
      btm_1[1] = {1'b0,layer_3_1[2863:2856]} - {1'b0, layer_2_1[2863:2856]};
      btm_1[2] = {1'b0,layer_3_1[2871:2864]} - {1'b0, layer_2_1[2871:2864]};
      btm_2[0] = {1'b0,layer_3_2[2855:2848]} - {1'b0, layer_2_2[2855:2848]};
      btm_2[1] = {1'b0,layer_3_2[2863:2856]} - {1'b0, layer_2_2[2863:2856]};
      btm_2[2] = {1'b0,layer_3_2[2871:2864]} - {1'b0, layer_2_2[2871:2864]};
    end
    'd358: begin
      top_0[0] = {1'b0,layer_1_0[2863:2856]} - {1'b0, layer_0_0[2863:2856]};
      top_0[1] = {1'b0,layer_1_0[2871:2864]} - {1'b0, layer_0_0[2871:2864]};
      top_0[2] = {1'b0,layer_1_0[2879:2872]} - {1'b0, layer_0_0[2879:2872]};
      top_1[0] = {1'b0,layer_1_1[2863:2856]} - {1'b0, layer_0_1[2863:2856]};
      top_1[1] = {1'b0,layer_1_1[2871:2864]} - {1'b0, layer_0_1[2871:2864]};
      top_1[2] = {1'b0,layer_1_1[2879:2872]} - {1'b0, layer_0_1[2879:2872]};
      top_2[0] = {1'b0,layer_1_2[2863:2856]} - {1'b0, layer_0_2[2863:2856]};
      top_2[1] = {1'b0,layer_1_2[2871:2864]} - {1'b0, layer_0_2[2871:2864]};
      top_2[2] = {1'b0,layer_1_2[2879:2872]} - {1'b0, layer_0_2[2879:2872]};
      mid_0[0] = {1'b0,layer_2_0[2863:2856]} - {1'b0, layer_1_0[2863:2856]};
      mid_0[1] = {1'b0,layer_2_0[2871:2864]} - {1'b0, layer_1_0[2871:2864]};
      mid_0[2] = {1'b0,layer_2_0[2879:2872]} - {1'b0, layer_1_0[2879:2872]};
      mid_1[0] = {1'b0,layer_2_1[2863:2856]} - {1'b0, layer_1_1[2863:2856]};
      mid_1[1] = {1'b0,layer_2_1[2871:2864]} - {1'b0, layer_1_1[2871:2864]};
      mid_1[2] = {1'b0,layer_2_1[2879:2872]} - {1'b0, layer_1_1[2879:2872]};
      mid_2[0] = {1'b0,layer_2_2[2863:2856]} - {1'b0, layer_1_2[2863:2856]};
      mid_2[1] = {1'b0,layer_2_2[2871:2864]} - {1'b0, layer_1_2[2871:2864]};
      mid_2[2] = {1'b0,layer_2_2[2879:2872]} - {1'b0, layer_1_2[2879:2872]};
      btm_0[0] = {1'b0,layer_3_0[2863:2856]} - {1'b0, layer_2_0[2863:2856]};
      btm_0[1] = {1'b0,layer_3_0[2871:2864]} - {1'b0, layer_2_0[2871:2864]};
      btm_0[2] = {1'b0,layer_3_0[2879:2872]} - {1'b0, layer_2_0[2879:2872]};
      btm_1[0] = {1'b0,layer_3_1[2863:2856]} - {1'b0, layer_2_1[2863:2856]};
      btm_1[1] = {1'b0,layer_3_1[2871:2864]} - {1'b0, layer_2_1[2871:2864]};
      btm_1[2] = {1'b0,layer_3_1[2879:2872]} - {1'b0, layer_2_1[2879:2872]};
      btm_2[0] = {1'b0,layer_3_2[2863:2856]} - {1'b0, layer_2_2[2863:2856]};
      btm_2[1] = {1'b0,layer_3_2[2871:2864]} - {1'b0, layer_2_2[2871:2864]};
      btm_2[2] = {1'b0,layer_3_2[2879:2872]} - {1'b0, layer_2_2[2879:2872]};
    end
    'd359: begin
      top_0[0] = {1'b0,layer_1_0[2871:2864]} - {1'b0, layer_0_0[2871:2864]};
      top_0[1] = {1'b0,layer_1_0[2879:2872]} - {1'b0, layer_0_0[2879:2872]};
      top_0[2] = {1'b0,layer_1_0[2887:2880]} - {1'b0, layer_0_0[2887:2880]};
      top_1[0] = {1'b0,layer_1_1[2871:2864]} - {1'b0, layer_0_1[2871:2864]};
      top_1[1] = {1'b0,layer_1_1[2879:2872]} - {1'b0, layer_0_1[2879:2872]};
      top_1[2] = {1'b0,layer_1_1[2887:2880]} - {1'b0, layer_0_1[2887:2880]};
      top_2[0] = {1'b0,layer_1_2[2871:2864]} - {1'b0, layer_0_2[2871:2864]};
      top_2[1] = {1'b0,layer_1_2[2879:2872]} - {1'b0, layer_0_2[2879:2872]};
      top_2[2] = {1'b0,layer_1_2[2887:2880]} - {1'b0, layer_0_2[2887:2880]};
      mid_0[0] = {1'b0,layer_2_0[2871:2864]} - {1'b0, layer_1_0[2871:2864]};
      mid_0[1] = {1'b0,layer_2_0[2879:2872]} - {1'b0, layer_1_0[2879:2872]};
      mid_0[2] = {1'b0,layer_2_0[2887:2880]} - {1'b0, layer_1_0[2887:2880]};
      mid_1[0] = {1'b0,layer_2_1[2871:2864]} - {1'b0, layer_1_1[2871:2864]};
      mid_1[1] = {1'b0,layer_2_1[2879:2872]} - {1'b0, layer_1_1[2879:2872]};
      mid_1[2] = {1'b0,layer_2_1[2887:2880]} - {1'b0, layer_1_1[2887:2880]};
      mid_2[0] = {1'b0,layer_2_2[2871:2864]} - {1'b0, layer_1_2[2871:2864]};
      mid_2[1] = {1'b0,layer_2_2[2879:2872]} - {1'b0, layer_1_2[2879:2872]};
      mid_2[2] = {1'b0,layer_2_2[2887:2880]} - {1'b0, layer_1_2[2887:2880]};
      btm_0[0] = {1'b0,layer_3_0[2871:2864]} - {1'b0, layer_2_0[2871:2864]};
      btm_0[1] = {1'b0,layer_3_0[2879:2872]} - {1'b0, layer_2_0[2879:2872]};
      btm_0[2] = {1'b0,layer_3_0[2887:2880]} - {1'b0, layer_2_0[2887:2880]};
      btm_1[0] = {1'b0,layer_3_1[2871:2864]} - {1'b0, layer_2_1[2871:2864]};
      btm_1[1] = {1'b0,layer_3_1[2879:2872]} - {1'b0, layer_2_1[2879:2872]};
      btm_1[2] = {1'b0,layer_3_1[2887:2880]} - {1'b0, layer_2_1[2887:2880]};
      btm_2[0] = {1'b0,layer_3_2[2871:2864]} - {1'b0, layer_2_2[2871:2864]};
      btm_2[1] = {1'b0,layer_3_2[2879:2872]} - {1'b0, layer_2_2[2879:2872]};
      btm_2[2] = {1'b0,layer_3_2[2887:2880]} - {1'b0, layer_2_2[2887:2880]};
    end
    'd360: begin
      top_0[0] = {1'b0,layer_1_0[2879:2872]} - {1'b0, layer_0_0[2879:2872]};
      top_0[1] = {1'b0,layer_1_0[2887:2880]} - {1'b0, layer_0_0[2887:2880]};
      top_0[2] = {1'b0,layer_1_0[2895:2888]} - {1'b0, layer_0_0[2895:2888]};
      top_1[0] = {1'b0,layer_1_1[2879:2872]} - {1'b0, layer_0_1[2879:2872]};
      top_1[1] = {1'b0,layer_1_1[2887:2880]} - {1'b0, layer_0_1[2887:2880]};
      top_1[2] = {1'b0,layer_1_1[2895:2888]} - {1'b0, layer_0_1[2895:2888]};
      top_2[0] = {1'b0,layer_1_2[2879:2872]} - {1'b0, layer_0_2[2879:2872]};
      top_2[1] = {1'b0,layer_1_2[2887:2880]} - {1'b0, layer_0_2[2887:2880]};
      top_2[2] = {1'b0,layer_1_2[2895:2888]} - {1'b0, layer_0_2[2895:2888]};
      mid_0[0] = {1'b0,layer_2_0[2879:2872]} - {1'b0, layer_1_0[2879:2872]};
      mid_0[1] = {1'b0,layer_2_0[2887:2880]} - {1'b0, layer_1_0[2887:2880]};
      mid_0[2] = {1'b0,layer_2_0[2895:2888]} - {1'b0, layer_1_0[2895:2888]};
      mid_1[0] = {1'b0,layer_2_1[2879:2872]} - {1'b0, layer_1_1[2879:2872]};
      mid_1[1] = {1'b0,layer_2_1[2887:2880]} - {1'b0, layer_1_1[2887:2880]};
      mid_1[2] = {1'b0,layer_2_1[2895:2888]} - {1'b0, layer_1_1[2895:2888]};
      mid_2[0] = {1'b0,layer_2_2[2879:2872]} - {1'b0, layer_1_2[2879:2872]};
      mid_2[1] = {1'b0,layer_2_2[2887:2880]} - {1'b0, layer_1_2[2887:2880]};
      mid_2[2] = {1'b0,layer_2_2[2895:2888]} - {1'b0, layer_1_2[2895:2888]};
      btm_0[0] = {1'b0,layer_3_0[2879:2872]} - {1'b0, layer_2_0[2879:2872]};
      btm_0[1] = {1'b0,layer_3_0[2887:2880]} - {1'b0, layer_2_0[2887:2880]};
      btm_0[2] = {1'b0,layer_3_0[2895:2888]} - {1'b0, layer_2_0[2895:2888]};
      btm_1[0] = {1'b0,layer_3_1[2879:2872]} - {1'b0, layer_2_1[2879:2872]};
      btm_1[1] = {1'b0,layer_3_1[2887:2880]} - {1'b0, layer_2_1[2887:2880]};
      btm_1[2] = {1'b0,layer_3_1[2895:2888]} - {1'b0, layer_2_1[2895:2888]};
      btm_2[0] = {1'b0,layer_3_2[2879:2872]} - {1'b0, layer_2_2[2879:2872]};
      btm_2[1] = {1'b0,layer_3_2[2887:2880]} - {1'b0, layer_2_2[2887:2880]};
      btm_2[2] = {1'b0,layer_3_2[2895:2888]} - {1'b0, layer_2_2[2895:2888]};
    end
    'd361: begin
      top_0[0] = {1'b0,layer_1_0[2887:2880]} - {1'b0, layer_0_0[2887:2880]};
      top_0[1] = {1'b0,layer_1_0[2895:2888]} - {1'b0, layer_0_0[2895:2888]};
      top_0[2] = {1'b0,layer_1_0[2903:2896]} - {1'b0, layer_0_0[2903:2896]};
      top_1[0] = {1'b0,layer_1_1[2887:2880]} - {1'b0, layer_0_1[2887:2880]};
      top_1[1] = {1'b0,layer_1_1[2895:2888]} - {1'b0, layer_0_1[2895:2888]};
      top_1[2] = {1'b0,layer_1_1[2903:2896]} - {1'b0, layer_0_1[2903:2896]};
      top_2[0] = {1'b0,layer_1_2[2887:2880]} - {1'b0, layer_0_2[2887:2880]};
      top_2[1] = {1'b0,layer_1_2[2895:2888]} - {1'b0, layer_0_2[2895:2888]};
      top_2[2] = {1'b0,layer_1_2[2903:2896]} - {1'b0, layer_0_2[2903:2896]};
      mid_0[0] = {1'b0,layer_2_0[2887:2880]} - {1'b0, layer_1_0[2887:2880]};
      mid_0[1] = {1'b0,layer_2_0[2895:2888]} - {1'b0, layer_1_0[2895:2888]};
      mid_0[2] = {1'b0,layer_2_0[2903:2896]} - {1'b0, layer_1_0[2903:2896]};
      mid_1[0] = {1'b0,layer_2_1[2887:2880]} - {1'b0, layer_1_1[2887:2880]};
      mid_1[1] = {1'b0,layer_2_1[2895:2888]} - {1'b0, layer_1_1[2895:2888]};
      mid_1[2] = {1'b0,layer_2_1[2903:2896]} - {1'b0, layer_1_1[2903:2896]};
      mid_2[0] = {1'b0,layer_2_2[2887:2880]} - {1'b0, layer_1_2[2887:2880]};
      mid_2[1] = {1'b0,layer_2_2[2895:2888]} - {1'b0, layer_1_2[2895:2888]};
      mid_2[2] = {1'b0,layer_2_2[2903:2896]} - {1'b0, layer_1_2[2903:2896]};
      btm_0[0] = {1'b0,layer_3_0[2887:2880]} - {1'b0, layer_2_0[2887:2880]};
      btm_0[1] = {1'b0,layer_3_0[2895:2888]} - {1'b0, layer_2_0[2895:2888]};
      btm_0[2] = {1'b0,layer_3_0[2903:2896]} - {1'b0, layer_2_0[2903:2896]};
      btm_1[0] = {1'b0,layer_3_1[2887:2880]} - {1'b0, layer_2_1[2887:2880]};
      btm_1[1] = {1'b0,layer_3_1[2895:2888]} - {1'b0, layer_2_1[2895:2888]};
      btm_1[2] = {1'b0,layer_3_1[2903:2896]} - {1'b0, layer_2_1[2903:2896]};
      btm_2[0] = {1'b0,layer_3_2[2887:2880]} - {1'b0, layer_2_2[2887:2880]};
      btm_2[1] = {1'b0,layer_3_2[2895:2888]} - {1'b0, layer_2_2[2895:2888]};
      btm_2[2] = {1'b0,layer_3_2[2903:2896]} - {1'b0, layer_2_2[2903:2896]};
    end
    'd362: begin
      top_0[0] = {1'b0,layer_1_0[2895:2888]} - {1'b0, layer_0_0[2895:2888]};
      top_0[1] = {1'b0,layer_1_0[2903:2896]} - {1'b0, layer_0_0[2903:2896]};
      top_0[2] = {1'b0,layer_1_0[2911:2904]} - {1'b0, layer_0_0[2911:2904]};
      top_1[0] = {1'b0,layer_1_1[2895:2888]} - {1'b0, layer_0_1[2895:2888]};
      top_1[1] = {1'b0,layer_1_1[2903:2896]} - {1'b0, layer_0_1[2903:2896]};
      top_1[2] = {1'b0,layer_1_1[2911:2904]} - {1'b0, layer_0_1[2911:2904]};
      top_2[0] = {1'b0,layer_1_2[2895:2888]} - {1'b0, layer_0_2[2895:2888]};
      top_2[1] = {1'b0,layer_1_2[2903:2896]} - {1'b0, layer_0_2[2903:2896]};
      top_2[2] = {1'b0,layer_1_2[2911:2904]} - {1'b0, layer_0_2[2911:2904]};
      mid_0[0] = {1'b0,layer_2_0[2895:2888]} - {1'b0, layer_1_0[2895:2888]};
      mid_0[1] = {1'b0,layer_2_0[2903:2896]} - {1'b0, layer_1_0[2903:2896]};
      mid_0[2] = {1'b0,layer_2_0[2911:2904]} - {1'b0, layer_1_0[2911:2904]};
      mid_1[0] = {1'b0,layer_2_1[2895:2888]} - {1'b0, layer_1_1[2895:2888]};
      mid_1[1] = {1'b0,layer_2_1[2903:2896]} - {1'b0, layer_1_1[2903:2896]};
      mid_1[2] = {1'b0,layer_2_1[2911:2904]} - {1'b0, layer_1_1[2911:2904]};
      mid_2[0] = {1'b0,layer_2_2[2895:2888]} - {1'b0, layer_1_2[2895:2888]};
      mid_2[1] = {1'b0,layer_2_2[2903:2896]} - {1'b0, layer_1_2[2903:2896]};
      mid_2[2] = {1'b0,layer_2_2[2911:2904]} - {1'b0, layer_1_2[2911:2904]};
      btm_0[0] = {1'b0,layer_3_0[2895:2888]} - {1'b0, layer_2_0[2895:2888]};
      btm_0[1] = {1'b0,layer_3_0[2903:2896]} - {1'b0, layer_2_0[2903:2896]};
      btm_0[2] = {1'b0,layer_3_0[2911:2904]} - {1'b0, layer_2_0[2911:2904]};
      btm_1[0] = {1'b0,layer_3_1[2895:2888]} - {1'b0, layer_2_1[2895:2888]};
      btm_1[1] = {1'b0,layer_3_1[2903:2896]} - {1'b0, layer_2_1[2903:2896]};
      btm_1[2] = {1'b0,layer_3_1[2911:2904]} - {1'b0, layer_2_1[2911:2904]};
      btm_2[0] = {1'b0,layer_3_2[2895:2888]} - {1'b0, layer_2_2[2895:2888]};
      btm_2[1] = {1'b0,layer_3_2[2903:2896]} - {1'b0, layer_2_2[2903:2896]};
      btm_2[2] = {1'b0,layer_3_2[2911:2904]} - {1'b0, layer_2_2[2911:2904]};
    end
    'd363: begin
      top_0[0] = {1'b0,layer_1_0[2903:2896]} - {1'b0, layer_0_0[2903:2896]};
      top_0[1] = {1'b0,layer_1_0[2911:2904]} - {1'b0, layer_0_0[2911:2904]};
      top_0[2] = {1'b0,layer_1_0[2919:2912]} - {1'b0, layer_0_0[2919:2912]};
      top_1[0] = {1'b0,layer_1_1[2903:2896]} - {1'b0, layer_0_1[2903:2896]};
      top_1[1] = {1'b0,layer_1_1[2911:2904]} - {1'b0, layer_0_1[2911:2904]};
      top_1[2] = {1'b0,layer_1_1[2919:2912]} - {1'b0, layer_0_1[2919:2912]};
      top_2[0] = {1'b0,layer_1_2[2903:2896]} - {1'b0, layer_0_2[2903:2896]};
      top_2[1] = {1'b0,layer_1_2[2911:2904]} - {1'b0, layer_0_2[2911:2904]};
      top_2[2] = {1'b0,layer_1_2[2919:2912]} - {1'b0, layer_0_2[2919:2912]};
      mid_0[0] = {1'b0,layer_2_0[2903:2896]} - {1'b0, layer_1_0[2903:2896]};
      mid_0[1] = {1'b0,layer_2_0[2911:2904]} - {1'b0, layer_1_0[2911:2904]};
      mid_0[2] = {1'b0,layer_2_0[2919:2912]} - {1'b0, layer_1_0[2919:2912]};
      mid_1[0] = {1'b0,layer_2_1[2903:2896]} - {1'b0, layer_1_1[2903:2896]};
      mid_1[1] = {1'b0,layer_2_1[2911:2904]} - {1'b0, layer_1_1[2911:2904]};
      mid_1[2] = {1'b0,layer_2_1[2919:2912]} - {1'b0, layer_1_1[2919:2912]};
      mid_2[0] = {1'b0,layer_2_2[2903:2896]} - {1'b0, layer_1_2[2903:2896]};
      mid_2[1] = {1'b0,layer_2_2[2911:2904]} - {1'b0, layer_1_2[2911:2904]};
      mid_2[2] = {1'b0,layer_2_2[2919:2912]} - {1'b0, layer_1_2[2919:2912]};
      btm_0[0] = {1'b0,layer_3_0[2903:2896]} - {1'b0, layer_2_0[2903:2896]};
      btm_0[1] = {1'b0,layer_3_0[2911:2904]} - {1'b0, layer_2_0[2911:2904]};
      btm_0[2] = {1'b0,layer_3_0[2919:2912]} - {1'b0, layer_2_0[2919:2912]};
      btm_1[0] = {1'b0,layer_3_1[2903:2896]} - {1'b0, layer_2_1[2903:2896]};
      btm_1[1] = {1'b0,layer_3_1[2911:2904]} - {1'b0, layer_2_1[2911:2904]};
      btm_1[2] = {1'b0,layer_3_1[2919:2912]} - {1'b0, layer_2_1[2919:2912]};
      btm_2[0] = {1'b0,layer_3_2[2903:2896]} - {1'b0, layer_2_2[2903:2896]};
      btm_2[1] = {1'b0,layer_3_2[2911:2904]} - {1'b0, layer_2_2[2911:2904]};
      btm_2[2] = {1'b0,layer_3_2[2919:2912]} - {1'b0, layer_2_2[2919:2912]};
    end
    'd364: begin
      top_0[0] = {1'b0,layer_1_0[2911:2904]} - {1'b0, layer_0_0[2911:2904]};
      top_0[1] = {1'b0,layer_1_0[2919:2912]} - {1'b0, layer_0_0[2919:2912]};
      top_0[2] = {1'b0,layer_1_0[2927:2920]} - {1'b0, layer_0_0[2927:2920]};
      top_1[0] = {1'b0,layer_1_1[2911:2904]} - {1'b0, layer_0_1[2911:2904]};
      top_1[1] = {1'b0,layer_1_1[2919:2912]} - {1'b0, layer_0_1[2919:2912]};
      top_1[2] = {1'b0,layer_1_1[2927:2920]} - {1'b0, layer_0_1[2927:2920]};
      top_2[0] = {1'b0,layer_1_2[2911:2904]} - {1'b0, layer_0_2[2911:2904]};
      top_2[1] = {1'b0,layer_1_2[2919:2912]} - {1'b0, layer_0_2[2919:2912]};
      top_2[2] = {1'b0,layer_1_2[2927:2920]} - {1'b0, layer_0_2[2927:2920]};
      mid_0[0] = {1'b0,layer_2_0[2911:2904]} - {1'b0, layer_1_0[2911:2904]};
      mid_0[1] = {1'b0,layer_2_0[2919:2912]} - {1'b0, layer_1_0[2919:2912]};
      mid_0[2] = {1'b0,layer_2_0[2927:2920]} - {1'b0, layer_1_0[2927:2920]};
      mid_1[0] = {1'b0,layer_2_1[2911:2904]} - {1'b0, layer_1_1[2911:2904]};
      mid_1[1] = {1'b0,layer_2_1[2919:2912]} - {1'b0, layer_1_1[2919:2912]};
      mid_1[2] = {1'b0,layer_2_1[2927:2920]} - {1'b0, layer_1_1[2927:2920]};
      mid_2[0] = {1'b0,layer_2_2[2911:2904]} - {1'b0, layer_1_2[2911:2904]};
      mid_2[1] = {1'b0,layer_2_2[2919:2912]} - {1'b0, layer_1_2[2919:2912]};
      mid_2[2] = {1'b0,layer_2_2[2927:2920]} - {1'b0, layer_1_2[2927:2920]};
      btm_0[0] = {1'b0,layer_3_0[2911:2904]} - {1'b0, layer_2_0[2911:2904]};
      btm_0[1] = {1'b0,layer_3_0[2919:2912]} - {1'b0, layer_2_0[2919:2912]};
      btm_0[2] = {1'b0,layer_3_0[2927:2920]} - {1'b0, layer_2_0[2927:2920]};
      btm_1[0] = {1'b0,layer_3_1[2911:2904]} - {1'b0, layer_2_1[2911:2904]};
      btm_1[1] = {1'b0,layer_3_1[2919:2912]} - {1'b0, layer_2_1[2919:2912]};
      btm_1[2] = {1'b0,layer_3_1[2927:2920]} - {1'b0, layer_2_1[2927:2920]};
      btm_2[0] = {1'b0,layer_3_2[2911:2904]} - {1'b0, layer_2_2[2911:2904]};
      btm_2[1] = {1'b0,layer_3_2[2919:2912]} - {1'b0, layer_2_2[2919:2912]};
      btm_2[2] = {1'b0,layer_3_2[2927:2920]} - {1'b0, layer_2_2[2927:2920]};
    end
    'd365: begin
      top_0[0] = {1'b0,layer_1_0[2919:2912]} - {1'b0, layer_0_0[2919:2912]};
      top_0[1] = {1'b0,layer_1_0[2927:2920]} - {1'b0, layer_0_0[2927:2920]};
      top_0[2] = {1'b0,layer_1_0[2935:2928]} - {1'b0, layer_0_0[2935:2928]};
      top_1[0] = {1'b0,layer_1_1[2919:2912]} - {1'b0, layer_0_1[2919:2912]};
      top_1[1] = {1'b0,layer_1_1[2927:2920]} - {1'b0, layer_0_1[2927:2920]};
      top_1[2] = {1'b0,layer_1_1[2935:2928]} - {1'b0, layer_0_1[2935:2928]};
      top_2[0] = {1'b0,layer_1_2[2919:2912]} - {1'b0, layer_0_2[2919:2912]};
      top_2[1] = {1'b0,layer_1_2[2927:2920]} - {1'b0, layer_0_2[2927:2920]};
      top_2[2] = {1'b0,layer_1_2[2935:2928]} - {1'b0, layer_0_2[2935:2928]};
      mid_0[0] = {1'b0,layer_2_0[2919:2912]} - {1'b0, layer_1_0[2919:2912]};
      mid_0[1] = {1'b0,layer_2_0[2927:2920]} - {1'b0, layer_1_0[2927:2920]};
      mid_0[2] = {1'b0,layer_2_0[2935:2928]} - {1'b0, layer_1_0[2935:2928]};
      mid_1[0] = {1'b0,layer_2_1[2919:2912]} - {1'b0, layer_1_1[2919:2912]};
      mid_1[1] = {1'b0,layer_2_1[2927:2920]} - {1'b0, layer_1_1[2927:2920]};
      mid_1[2] = {1'b0,layer_2_1[2935:2928]} - {1'b0, layer_1_1[2935:2928]};
      mid_2[0] = {1'b0,layer_2_2[2919:2912]} - {1'b0, layer_1_2[2919:2912]};
      mid_2[1] = {1'b0,layer_2_2[2927:2920]} - {1'b0, layer_1_2[2927:2920]};
      mid_2[2] = {1'b0,layer_2_2[2935:2928]} - {1'b0, layer_1_2[2935:2928]};
      btm_0[0] = {1'b0,layer_3_0[2919:2912]} - {1'b0, layer_2_0[2919:2912]};
      btm_0[1] = {1'b0,layer_3_0[2927:2920]} - {1'b0, layer_2_0[2927:2920]};
      btm_0[2] = {1'b0,layer_3_0[2935:2928]} - {1'b0, layer_2_0[2935:2928]};
      btm_1[0] = {1'b0,layer_3_1[2919:2912]} - {1'b0, layer_2_1[2919:2912]};
      btm_1[1] = {1'b0,layer_3_1[2927:2920]} - {1'b0, layer_2_1[2927:2920]};
      btm_1[2] = {1'b0,layer_3_1[2935:2928]} - {1'b0, layer_2_1[2935:2928]};
      btm_2[0] = {1'b0,layer_3_2[2919:2912]} - {1'b0, layer_2_2[2919:2912]};
      btm_2[1] = {1'b0,layer_3_2[2927:2920]} - {1'b0, layer_2_2[2927:2920]};
      btm_2[2] = {1'b0,layer_3_2[2935:2928]} - {1'b0, layer_2_2[2935:2928]};
    end
    'd366: begin
      top_0[0] = {1'b0,layer_1_0[2927:2920]} - {1'b0, layer_0_0[2927:2920]};
      top_0[1] = {1'b0,layer_1_0[2935:2928]} - {1'b0, layer_0_0[2935:2928]};
      top_0[2] = {1'b0,layer_1_0[2943:2936]} - {1'b0, layer_0_0[2943:2936]};
      top_1[0] = {1'b0,layer_1_1[2927:2920]} - {1'b0, layer_0_1[2927:2920]};
      top_1[1] = {1'b0,layer_1_1[2935:2928]} - {1'b0, layer_0_1[2935:2928]};
      top_1[2] = {1'b0,layer_1_1[2943:2936]} - {1'b0, layer_0_1[2943:2936]};
      top_2[0] = {1'b0,layer_1_2[2927:2920]} - {1'b0, layer_0_2[2927:2920]};
      top_2[1] = {1'b0,layer_1_2[2935:2928]} - {1'b0, layer_0_2[2935:2928]};
      top_2[2] = {1'b0,layer_1_2[2943:2936]} - {1'b0, layer_0_2[2943:2936]};
      mid_0[0] = {1'b0,layer_2_0[2927:2920]} - {1'b0, layer_1_0[2927:2920]};
      mid_0[1] = {1'b0,layer_2_0[2935:2928]} - {1'b0, layer_1_0[2935:2928]};
      mid_0[2] = {1'b0,layer_2_0[2943:2936]} - {1'b0, layer_1_0[2943:2936]};
      mid_1[0] = {1'b0,layer_2_1[2927:2920]} - {1'b0, layer_1_1[2927:2920]};
      mid_1[1] = {1'b0,layer_2_1[2935:2928]} - {1'b0, layer_1_1[2935:2928]};
      mid_1[2] = {1'b0,layer_2_1[2943:2936]} - {1'b0, layer_1_1[2943:2936]};
      mid_2[0] = {1'b0,layer_2_2[2927:2920]} - {1'b0, layer_1_2[2927:2920]};
      mid_2[1] = {1'b0,layer_2_2[2935:2928]} - {1'b0, layer_1_2[2935:2928]};
      mid_2[2] = {1'b0,layer_2_2[2943:2936]} - {1'b0, layer_1_2[2943:2936]};
      btm_0[0] = {1'b0,layer_3_0[2927:2920]} - {1'b0, layer_2_0[2927:2920]};
      btm_0[1] = {1'b0,layer_3_0[2935:2928]} - {1'b0, layer_2_0[2935:2928]};
      btm_0[2] = {1'b0,layer_3_0[2943:2936]} - {1'b0, layer_2_0[2943:2936]};
      btm_1[0] = {1'b0,layer_3_1[2927:2920]} - {1'b0, layer_2_1[2927:2920]};
      btm_1[1] = {1'b0,layer_3_1[2935:2928]} - {1'b0, layer_2_1[2935:2928]};
      btm_1[2] = {1'b0,layer_3_1[2943:2936]} - {1'b0, layer_2_1[2943:2936]};
      btm_2[0] = {1'b0,layer_3_2[2927:2920]} - {1'b0, layer_2_2[2927:2920]};
      btm_2[1] = {1'b0,layer_3_2[2935:2928]} - {1'b0, layer_2_2[2935:2928]};
      btm_2[2] = {1'b0,layer_3_2[2943:2936]} - {1'b0, layer_2_2[2943:2936]};
    end
    'd367: begin
      top_0[0] = {1'b0,layer_1_0[2935:2928]} - {1'b0, layer_0_0[2935:2928]};
      top_0[1] = {1'b0,layer_1_0[2943:2936]} - {1'b0, layer_0_0[2943:2936]};
      top_0[2] = {1'b0,layer_1_0[2951:2944]} - {1'b0, layer_0_0[2951:2944]};
      top_1[0] = {1'b0,layer_1_1[2935:2928]} - {1'b0, layer_0_1[2935:2928]};
      top_1[1] = {1'b0,layer_1_1[2943:2936]} - {1'b0, layer_0_1[2943:2936]};
      top_1[2] = {1'b0,layer_1_1[2951:2944]} - {1'b0, layer_0_1[2951:2944]};
      top_2[0] = {1'b0,layer_1_2[2935:2928]} - {1'b0, layer_0_2[2935:2928]};
      top_2[1] = {1'b0,layer_1_2[2943:2936]} - {1'b0, layer_0_2[2943:2936]};
      top_2[2] = {1'b0,layer_1_2[2951:2944]} - {1'b0, layer_0_2[2951:2944]};
      mid_0[0] = {1'b0,layer_2_0[2935:2928]} - {1'b0, layer_1_0[2935:2928]};
      mid_0[1] = {1'b0,layer_2_0[2943:2936]} - {1'b0, layer_1_0[2943:2936]};
      mid_0[2] = {1'b0,layer_2_0[2951:2944]} - {1'b0, layer_1_0[2951:2944]};
      mid_1[0] = {1'b0,layer_2_1[2935:2928]} - {1'b0, layer_1_1[2935:2928]};
      mid_1[1] = {1'b0,layer_2_1[2943:2936]} - {1'b0, layer_1_1[2943:2936]};
      mid_1[2] = {1'b0,layer_2_1[2951:2944]} - {1'b0, layer_1_1[2951:2944]};
      mid_2[0] = {1'b0,layer_2_2[2935:2928]} - {1'b0, layer_1_2[2935:2928]};
      mid_2[1] = {1'b0,layer_2_2[2943:2936]} - {1'b0, layer_1_2[2943:2936]};
      mid_2[2] = {1'b0,layer_2_2[2951:2944]} - {1'b0, layer_1_2[2951:2944]};
      btm_0[0] = {1'b0,layer_3_0[2935:2928]} - {1'b0, layer_2_0[2935:2928]};
      btm_0[1] = {1'b0,layer_3_0[2943:2936]} - {1'b0, layer_2_0[2943:2936]};
      btm_0[2] = {1'b0,layer_3_0[2951:2944]} - {1'b0, layer_2_0[2951:2944]};
      btm_1[0] = {1'b0,layer_3_1[2935:2928]} - {1'b0, layer_2_1[2935:2928]};
      btm_1[1] = {1'b0,layer_3_1[2943:2936]} - {1'b0, layer_2_1[2943:2936]};
      btm_1[2] = {1'b0,layer_3_1[2951:2944]} - {1'b0, layer_2_1[2951:2944]};
      btm_2[0] = {1'b0,layer_3_2[2935:2928]} - {1'b0, layer_2_2[2935:2928]};
      btm_2[1] = {1'b0,layer_3_2[2943:2936]} - {1'b0, layer_2_2[2943:2936]};
      btm_2[2] = {1'b0,layer_3_2[2951:2944]} - {1'b0, layer_2_2[2951:2944]};
    end
    'd368: begin
      top_0[0] = {1'b0,layer_1_0[2943:2936]} - {1'b0, layer_0_0[2943:2936]};
      top_0[1] = {1'b0,layer_1_0[2951:2944]} - {1'b0, layer_0_0[2951:2944]};
      top_0[2] = {1'b0,layer_1_0[2959:2952]} - {1'b0, layer_0_0[2959:2952]};
      top_1[0] = {1'b0,layer_1_1[2943:2936]} - {1'b0, layer_0_1[2943:2936]};
      top_1[1] = {1'b0,layer_1_1[2951:2944]} - {1'b0, layer_0_1[2951:2944]};
      top_1[2] = {1'b0,layer_1_1[2959:2952]} - {1'b0, layer_0_1[2959:2952]};
      top_2[0] = {1'b0,layer_1_2[2943:2936]} - {1'b0, layer_0_2[2943:2936]};
      top_2[1] = {1'b0,layer_1_2[2951:2944]} - {1'b0, layer_0_2[2951:2944]};
      top_2[2] = {1'b0,layer_1_2[2959:2952]} - {1'b0, layer_0_2[2959:2952]};
      mid_0[0] = {1'b0,layer_2_0[2943:2936]} - {1'b0, layer_1_0[2943:2936]};
      mid_0[1] = {1'b0,layer_2_0[2951:2944]} - {1'b0, layer_1_0[2951:2944]};
      mid_0[2] = {1'b0,layer_2_0[2959:2952]} - {1'b0, layer_1_0[2959:2952]};
      mid_1[0] = {1'b0,layer_2_1[2943:2936]} - {1'b0, layer_1_1[2943:2936]};
      mid_1[1] = {1'b0,layer_2_1[2951:2944]} - {1'b0, layer_1_1[2951:2944]};
      mid_1[2] = {1'b0,layer_2_1[2959:2952]} - {1'b0, layer_1_1[2959:2952]};
      mid_2[0] = {1'b0,layer_2_2[2943:2936]} - {1'b0, layer_1_2[2943:2936]};
      mid_2[1] = {1'b0,layer_2_2[2951:2944]} - {1'b0, layer_1_2[2951:2944]};
      mid_2[2] = {1'b0,layer_2_2[2959:2952]} - {1'b0, layer_1_2[2959:2952]};
      btm_0[0] = {1'b0,layer_3_0[2943:2936]} - {1'b0, layer_2_0[2943:2936]};
      btm_0[1] = {1'b0,layer_3_0[2951:2944]} - {1'b0, layer_2_0[2951:2944]};
      btm_0[2] = {1'b0,layer_3_0[2959:2952]} - {1'b0, layer_2_0[2959:2952]};
      btm_1[0] = {1'b0,layer_3_1[2943:2936]} - {1'b0, layer_2_1[2943:2936]};
      btm_1[1] = {1'b0,layer_3_1[2951:2944]} - {1'b0, layer_2_1[2951:2944]};
      btm_1[2] = {1'b0,layer_3_1[2959:2952]} - {1'b0, layer_2_1[2959:2952]};
      btm_2[0] = {1'b0,layer_3_2[2943:2936]} - {1'b0, layer_2_2[2943:2936]};
      btm_2[1] = {1'b0,layer_3_2[2951:2944]} - {1'b0, layer_2_2[2951:2944]};
      btm_2[2] = {1'b0,layer_3_2[2959:2952]} - {1'b0, layer_2_2[2959:2952]};
    end
    'd369: begin
      top_0[0] = {1'b0,layer_1_0[2951:2944]} - {1'b0, layer_0_0[2951:2944]};
      top_0[1] = {1'b0,layer_1_0[2959:2952]} - {1'b0, layer_0_0[2959:2952]};
      top_0[2] = {1'b0,layer_1_0[2967:2960]} - {1'b0, layer_0_0[2967:2960]};
      top_1[0] = {1'b0,layer_1_1[2951:2944]} - {1'b0, layer_0_1[2951:2944]};
      top_1[1] = {1'b0,layer_1_1[2959:2952]} - {1'b0, layer_0_1[2959:2952]};
      top_1[2] = {1'b0,layer_1_1[2967:2960]} - {1'b0, layer_0_1[2967:2960]};
      top_2[0] = {1'b0,layer_1_2[2951:2944]} - {1'b0, layer_0_2[2951:2944]};
      top_2[1] = {1'b0,layer_1_2[2959:2952]} - {1'b0, layer_0_2[2959:2952]};
      top_2[2] = {1'b0,layer_1_2[2967:2960]} - {1'b0, layer_0_2[2967:2960]};
      mid_0[0] = {1'b0,layer_2_0[2951:2944]} - {1'b0, layer_1_0[2951:2944]};
      mid_0[1] = {1'b0,layer_2_0[2959:2952]} - {1'b0, layer_1_0[2959:2952]};
      mid_0[2] = {1'b0,layer_2_0[2967:2960]} - {1'b0, layer_1_0[2967:2960]};
      mid_1[0] = {1'b0,layer_2_1[2951:2944]} - {1'b0, layer_1_1[2951:2944]};
      mid_1[1] = {1'b0,layer_2_1[2959:2952]} - {1'b0, layer_1_1[2959:2952]};
      mid_1[2] = {1'b0,layer_2_1[2967:2960]} - {1'b0, layer_1_1[2967:2960]};
      mid_2[0] = {1'b0,layer_2_2[2951:2944]} - {1'b0, layer_1_2[2951:2944]};
      mid_2[1] = {1'b0,layer_2_2[2959:2952]} - {1'b0, layer_1_2[2959:2952]};
      mid_2[2] = {1'b0,layer_2_2[2967:2960]} - {1'b0, layer_1_2[2967:2960]};
      btm_0[0] = {1'b0,layer_3_0[2951:2944]} - {1'b0, layer_2_0[2951:2944]};
      btm_0[1] = {1'b0,layer_3_0[2959:2952]} - {1'b0, layer_2_0[2959:2952]};
      btm_0[2] = {1'b0,layer_3_0[2967:2960]} - {1'b0, layer_2_0[2967:2960]};
      btm_1[0] = {1'b0,layer_3_1[2951:2944]} - {1'b0, layer_2_1[2951:2944]};
      btm_1[1] = {1'b0,layer_3_1[2959:2952]} - {1'b0, layer_2_1[2959:2952]};
      btm_1[2] = {1'b0,layer_3_1[2967:2960]} - {1'b0, layer_2_1[2967:2960]};
      btm_2[0] = {1'b0,layer_3_2[2951:2944]} - {1'b0, layer_2_2[2951:2944]};
      btm_2[1] = {1'b0,layer_3_2[2959:2952]} - {1'b0, layer_2_2[2959:2952]};
      btm_2[2] = {1'b0,layer_3_2[2967:2960]} - {1'b0, layer_2_2[2967:2960]};
    end
    'd370: begin
      top_0[0] = {1'b0,layer_1_0[2959:2952]} - {1'b0, layer_0_0[2959:2952]};
      top_0[1] = {1'b0,layer_1_0[2967:2960]} - {1'b0, layer_0_0[2967:2960]};
      top_0[2] = {1'b0,layer_1_0[2975:2968]} - {1'b0, layer_0_0[2975:2968]};
      top_1[0] = {1'b0,layer_1_1[2959:2952]} - {1'b0, layer_0_1[2959:2952]};
      top_1[1] = {1'b0,layer_1_1[2967:2960]} - {1'b0, layer_0_1[2967:2960]};
      top_1[2] = {1'b0,layer_1_1[2975:2968]} - {1'b0, layer_0_1[2975:2968]};
      top_2[0] = {1'b0,layer_1_2[2959:2952]} - {1'b0, layer_0_2[2959:2952]};
      top_2[1] = {1'b0,layer_1_2[2967:2960]} - {1'b0, layer_0_2[2967:2960]};
      top_2[2] = {1'b0,layer_1_2[2975:2968]} - {1'b0, layer_0_2[2975:2968]};
      mid_0[0] = {1'b0,layer_2_0[2959:2952]} - {1'b0, layer_1_0[2959:2952]};
      mid_0[1] = {1'b0,layer_2_0[2967:2960]} - {1'b0, layer_1_0[2967:2960]};
      mid_0[2] = {1'b0,layer_2_0[2975:2968]} - {1'b0, layer_1_0[2975:2968]};
      mid_1[0] = {1'b0,layer_2_1[2959:2952]} - {1'b0, layer_1_1[2959:2952]};
      mid_1[1] = {1'b0,layer_2_1[2967:2960]} - {1'b0, layer_1_1[2967:2960]};
      mid_1[2] = {1'b0,layer_2_1[2975:2968]} - {1'b0, layer_1_1[2975:2968]};
      mid_2[0] = {1'b0,layer_2_2[2959:2952]} - {1'b0, layer_1_2[2959:2952]};
      mid_2[1] = {1'b0,layer_2_2[2967:2960]} - {1'b0, layer_1_2[2967:2960]};
      mid_2[2] = {1'b0,layer_2_2[2975:2968]} - {1'b0, layer_1_2[2975:2968]};
      btm_0[0] = {1'b0,layer_3_0[2959:2952]} - {1'b0, layer_2_0[2959:2952]};
      btm_0[1] = {1'b0,layer_3_0[2967:2960]} - {1'b0, layer_2_0[2967:2960]};
      btm_0[2] = {1'b0,layer_3_0[2975:2968]} - {1'b0, layer_2_0[2975:2968]};
      btm_1[0] = {1'b0,layer_3_1[2959:2952]} - {1'b0, layer_2_1[2959:2952]};
      btm_1[1] = {1'b0,layer_3_1[2967:2960]} - {1'b0, layer_2_1[2967:2960]};
      btm_1[2] = {1'b0,layer_3_1[2975:2968]} - {1'b0, layer_2_1[2975:2968]};
      btm_2[0] = {1'b0,layer_3_2[2959:2952]} - {1'b0, layer_2_2[2959:2952]};
      btm_2[1] = {1'b0,layer_3_2[2967:2960]} - {1'b0, layer_2_2[2967:2960]};
      btm_2[2] = {1'b0,layer_3_2[2975:2968]} - {1'b0, layer_2_2[2975:2968]};
    end
    'd371: begin
      top_0[0] = {1'b0,layer_1_0[2967:2960]} - {1'b0, layer_0_0[2967:2960]};
      top_0[1] = {1'b0,layer_1_0[2975:2968]} - {1'b0, layer_0_0[2975:2968]};
      top_0[2] = {1'b0,layer_1_0[2983:2976]} - {1'b0, layer_0_0[2983:2976]};
      top_1[0] = {1'b0,layer_1_1[2967:2960]} - {1'b0, layer_0_1[2967:2960]};
      top_1[1] = {1'b0,layer_1_1[2975:2968]} - {1'b0, layer_0_1[2975:2968]};
      top_1[2] = {1'b0,layer_1_1[2983:2976]} - {1'b0, layer_0_1[2983:2976]};
      top_2[0] = {1'b0,layer_1_2[2967:2960]} - {1'b0, layer_0_2[2967:2960]};
      top_2[1] = {1'b0,layer_1_2[2975:2968]} - {1'b0, layer_0_2[2975:2968]};
      top_2[2] = {1'b0,layer_1_2[2983:2976]} - {1'b0, layer_0_2[2983:2976]};
      mid_0[0] = {1'b0,layer_2_0[2967:2960]} - {1'b0, layer_1_0[2967:2960]};
      mid_0[1] = {1'b0,layer_2_0[2975:2968]} - {1'b0, layer_1_0[2975:2968]};
      mid_0[2] = {1'b0,layer_2_0[2983:2976]} - {1'b0, layer_1_0[2983:2976]};
      mid_1[0] = {1'b0,layer_2_1[2967:2960]} - {1'b0, layer_1_1[2967:2960]};
      mid_1[1] = {1'b0,layer_2_1[2975:2968]} - {1'b0, layer_1_1[2975:2968]};
      mid_1[2] = {1'b0,layer_2_1[2983:2976]} - {1'b0, layer_1_1[2983:2976]};
      mid_2[0] = {1'b0,layer_2_2[2967:2960]} - {1'b0, layer_1_2[2967:2960]};
      mid_2[1] = {1'b0,layer_2_2[2975:2968]} - {1'b0, layer_1_2[2975:2968]};
      mid_2[2] = {1'b0,layer_2_2[2983:2976]} - {1'b0, layer_1_2[2983:2976]};
      btm_0[0] = {1'b0,layer_3_0[2967:2960]} - {1'b0, layer_2_0[2967:2960]};
      btm_0[1] = {1'b0,layer_3_0[2975:2968]} - {1'b0, layer_2_0[2975:2968]};
      btm_0[2] = {1'b0,layer_3_0[2983:2976]} - {1'b0, layer_2_0[2983:2976]};
      btm_1[0] = {1'b0,layer_3_1[2967:2960]} - {1'b0, layer_2_1[2967:2960]};
      btm_1[1] = {1'b0,layer_3_1[2975:2968]} - {1'b0, layer_2_1[2975:2968]};
      btm_1[2] = {1'b0,layer_3_1[2983:2976]} - {1'b0, layer_2_1[2983:2976]};
      btm_2[0] = {1'b0,layer_3_2[2967:2960]} - {1'b0, layer_2_2[2967:2960]};
      btm_2[1] = {1'b0,layer_3_2[2975:2968]} - {1'b0, layer_2_2[2975:2968]};
      btm_2[2] = {1'b0,layer_3_2[2983:2976]} - {1'b0, layer_2_2[2983:2976]};
    end
    'd372: begin
      top_0[0] = {1'b0,layer_1_0[2975:2968]} - {1'b0, layer_0_0[2975:2968]};
      top_0[1] = {1'b0,layer_1_0[2983:2976]} - {1'b0, layer_0_0[2983:2976]};
      top_0[2] = {1'b0,layer_1_0[2991:2984]} - {1'b0, layer_0_0[2991:2984]};
      top_1[0] = {1'b0,layer_1_1[2975:2968]} - {1'b0, layer_0_1[2975:2968]};
      top_1[1] = {1'b0,layer_1_1[2983:2976]} - {1'b0, layer_0_1[2983:2976]};
      top_1[2] = {1'b0,layer_1_1[2991:2984]} - {1'b0, layer_0_1[2991:2984]};
      top_2[0] = {1'b0,layer_1_2[2975:2968]} - {1'b0, layer_0_2[2975:2968]};
      top_2[1] = {1'b0,layer_1_2[2983:2976]} - {1'b0, layer_0_2[2983:2976]};
      top_2[2] = {1'b0,layer_1_2[2991:2984]} - {1'b0, layer_0_2[2991:2984]};
      mid_0[0] = {1'b0,layer_2_0[2975:2968]} - {1'b0, layer_1_0[2975:2968]};
      mid_0[1] = {1'b0,layer_2_0[2983:2976]} - {1'b0, layer_1_0[2983:2976]};
      mid_0[2] = {1'b0,layer_2_0[2991:2984]} - {1'b0, layer_1_0[2991:2984]};
      mid_1[0] = {1'b0,layer_2_1[2975:2968]} - {1'b0, layer_1_1[2975:2968]};
      mid_1[1] = {1'b0,layer_2_1[2983:2976]} - {1'b0, layer_1_1[2983:2976]};
      mid_1[2] = {1'b0,layer_2_1[2991:2984]} - {1'b0, layer_1_1[2991:2984]};
      mid_2[0] = {1'b0,layer_2_2[2975:2968]} - {1'b0, layer_1_2[2975:2968]};
      mid_2[1] = {1'b0,layer_2_2[2983:2976]} - {1'b0, layer_1_2[2983:2976]};
      mid_2[2] = {1'b0,layer_2_2[2991:2984]} - {1'b0, layer_1_2[2991:2984]};
      btm_0[0] = {1'b0,layer_3_0[2975:2968]} - {1'b0, layer_2_0[2975:2968]};
      btm_0[1] = {1'b0,layer_3_0[2983:2976]} - {1'b0, layer_2_0[2983:2976]};
      btm_0[2] = {1'b0,layer_3_0[2991:2984]} - {1'b0, layer_2_0[2991:2984]};
      btm_1[0] = {1'b0,layer_3_1[2975:2968]} - {1'b0, layer_2_1[2975:2968]};
      btm_1[1] = {1'b0,layer_3_1[2983:2976]} - {1'b0, layer_2_1[2983:2976]};
      btm_1[2] = {1'b0,layer_3_1[2991:2984]} - {1'b0, layer_2_1[2991:2984]};
      btm_2[0] = {1'b0,layer_3_2[2975:2968]} - {1'b0, layer_2_2[2975:2968]};
      btm_2[1] = {1'b0,layer_3_2[2983:2976]} - {1'b0, layer_2_2[2983:2976]};
      btm_2[2] = {1'b0,layer_3_2[2991:2984]} - {1'b0, layer_2_2[2991:2984]};
    end
    'd373: begin
      top_0[0] = {1'b0,layer_1_0[2983:2976]} - {1'b0, layer_0_0[2983:2976]};
      top_0[1] = {1'b0,layer_1_0[2991:2984]} - {1'b0, layer_0_0[2991:2984]};
      top_0[2] = {1'b0,layer_1_0[2999:2992]} - {1'b0, layer_0_0[2999:2992]};
      top_1[0] = {1'b0,layer_1_1[2983:2976]} - {1'b0, layer_0_1[2983:2976]};
      top_1[1] = {1'b0,layer_1_1[2991:2984]} - {1'b0, layer_0_1[2991:2984]};
      top_1[2] = {1'b0,layer_1_1[2999:2992]} - {1'b0, layer_0_1[2999:2992]};
      top_2[0] = {1'b0,layer_1_2[2983:2976]} - {1'b0, layer_0_2[2983:2976]};
      top_2[1] = {1'b0,layer_1_2[2991:2984]} - {1'b0, layer_0_2[2991:2984]};
      top_2[2] = {1'b0,layer_1_2[2999:2992]} - {1'b0, layer_0_2[2999:2992]};
      mid_0[0] = {1'b0,layer_2_0[2983:2976]} - {1'b0, layer_1_0[2983:2976]};
      mid_0[1] = {1'b0,layer_2_0[2991:2984]} - {1'b0, layer_1_0[2991:2984]};
      mid_0[2] = {1'b0,layer_2_0[2999:2992]} - {1'b0, layer_1_0[2999:2992]};
      mid_1[0] = {1'b0,layer_2_1[2983:2976]} - {1'b0, layer_1_1[2983:2976]};
      mid_1[1] = {1'b0,layer_2_1[2991:2984]} - {1'b0, layer_1_1[2991:2984]};
      mid_1[2] = {1'b0,layer_2_1[2999:2992]} - {1'b0, layer_1_1[2999:2992]};
      mid_2[0] = {1'b0,layer_2_2[2983:2976]} - {1'b0, layer_1_2[2983:2976]};
      mid_2[1] = {1'b0,layer_2_2[2991:2984]} - {1'b0, layer_1_2[2991:2984]};
      mid_2[2] = {1'b0,layer_2_2[2999:2992]} - {1'b0, layer_1_2[2999:2992]};
      btm_0[0] = {1'b0,layer_3_0[2983:2976]} - {1'b0, layer_2_0[2983:2976]};
      btm_0[1] = {1'b0,layer_3_0[2991:2984]} - {1'b0, layer_2_0[2991:2984]};
      btm_0[2] = {1'b0,layer_3_0[2999:2992]} - {1'b0, layer_2_0[2999:2992]};
      btm_1[0] = {1'b0,layer_3_1[2983:2976]} - {1'b0, layer_2_1[2983:2976]};
      btm_1[1] = {1'b0,layer_3_1[2991:2984]} - {1'b0, layer_2_1[2991:2984]};
      btm_1[2] = {1'b0,layer_3_1[2999:2992]} - {1'b0, layer_2_1[2999:2992]};
      btm_2[0] = {1'b0,layer_3_2[2983:2976]} - {1'b0, layer_2_2[2983:2976]};
      btm_2[1] = {1'b0,layer_3_2[2991:2984]} - {1'b0, layer_2_2[2991:2984]};
      btm_2[2] = {1'b0,layer_3_2[2999:2992]} - {1'b0, layer_2_2[2999:2992]};
    end
    'd374: begin
      top_0[0] = {1'b0,layer_1_0[2991:2984]} - {1'b0, layer_0_0[2991:2984]};
      top_0[1] = {1'b0,layer_1_0[2999:2992]} - {1'b0, layer_0_0[2999:2992]};
      top_0[2] = {1'b0,layer_1_0[3007:3000]} - {1'b0, layer_0_0[3007:3000]};
      top_1[0] = {1'b0,layer_1_1[2991:2984]} - {1'b0, layer_0_1[2991:2984]};
      top_1[1] = {1'b0,layer_1_1[2999:2992]} - {1'b0, layer_0_1[2999:2992]};
      top_1[2] = {1'b0,layer_1_1[3007:3000]} - {1'b0, layer_0_1[3007:3000]};
      top_2[0] = {1'b0,layer_1_2[2991:2984]} - {1'b0, layer_0_2[2991:2984]};
      top_2[1] = {1'b0,layer_1_2[2999:2992]} - {1'b0, layer_0_2[2999:2992]};
      top_2[2] = {1'b0,layer_1_2[3007:3000]} - {1'b0, layer_0_2[3007:3000]};
      mid_0[0] = {1'b0,layer_2_0[2991:2984]} - {1'b0, layer_1_0[2991:2984]};
      mid_0[1] = {1'b0,layer_2_0[2999:2992]} - {1'b0, layer_1_0[2999:2992]};
      mid_0[2] = {1'b0,layer_2_0[3007:3000]} - {1'b0, layer_1_0[3007:3000]};
      mid_1[0] = {1'b0,layer_2_1[2991:2984]} - {1'b0, layer_1_1[2991:2984]};
      mid_1[1] = {1'b0,layer_2_1[2999:2992]} - {1'b0, layer_1_1[2999:2992]};
      mid_1[2] = {1'b0,layer_2_1[3007:3000]} - {1'b0, layer_1_1[3007:3000]};
      mid_2[0] = {1'b0,layer_2_2[2991:2984]} - {1'b0, layer_1_2[2991:2984]};
      mid_2[1] = {1'b0,layer_2_2[2999:2992]} - {1'b0, layer_1_2[2999:2992]};
      mid_2[2] = {1'b0,layer_2_2[3007:3000]} - {1'b0, layer_1_2[3007:3000]};
      btm_0[0] = {1'b0,layer_3_0[2991:2984]} - {1'b0, layer_2_0[2991:2984]};
      btm_0[1] = {1'b0,layer_3_0[2999:2992]} - {1'b0, layer_2_0[2999:2992]};
      btm_0[2] = {1'b0,layer_3_0[3007:3000]} - {1'b0, layer_2_0[3007:3000]};
      btm_1[0] = {1'b0,layer_3_1[2991:2984]} - {1'b0, layer_2_1[2991:2984]};
      btm_1[1] = {1'b0,layer_3_1[2999:2992]} - {1'b0, layer_2_1[2999:2992]};
      btm_1[2] = {1'b0,layer_3_1[3007:3000]} - {1'b0, layer_2_1[3007:3000]};
      btm_2[0] = {1'b0,layer_3_2[2991:2984]} - {1'b0, layer_2_2[2991:2984]};
      btm_2[1] = {1'b0,layer_3_2[2999:2992]} - {1'b0, layer_2_2[2999:2992]};
      btm_2[2] = {1'b0,layer_3_2[3007:3000]} - {1'b0, layer_2_2[3007:3000]};
    end
    'd375: begin
      top_0[0] = {1'b0,layer_1_0[2999:2992]} - {1'b0, layer_0_0[2999:2992]};
      top_0[1] = {1'b0,layer_1_0[3007:3000]} - {1'b0, layer_0_0[3007:3000]};
      top_0[2] = {1'b0,layer_1_0[3015:3008]} - {1'b0, layer_0_0[3015:3008]};
      top_1[0] = {1'b0,layer_1_1[2999:2992]} - {1'b0, layer_0_1[2999:2992]};
      top_1[1] = {1'b0,layer_1_1[3007:3000]} - {1'b0, layer_0_1[3007:3000]};
      top_1[2] = {1'b0,layer_1_1[3015:3008]} - {1'b0, layer_0_1[3015:3008]};
      top_2[0] = {1'b0,layer_1_2[2999:2992]} - {1'b0, layer_0_2[2999:2992]};
      top_2[1] = {1'b0,layer_1_2[3007:3000]} - {1'b0, layer_0_2[3007:3000]};
      top_2[2] = {1'b0,layer_1_2[3015:3008]} - {1'b0, layer_0_2[3015:3008]};
      mid_0[0] = {1'b0,layer_2_0[2999:2992]} - {1'b0, layer_1_0[2999:2992]};
      mid_0[1] = {1'b0,layer_2_0[3007:3000]} - {1'b0, layer_1_0[3007:3000]};
      mid_0[2] = {1'b0,layer_2_0[3015:3008]} - {1'b0, layer_1_0[3015:3008]};
      mid_1[0] = {1'b0,layer_2_1[2999:2992]} - {1'b0, layer_1_1[2999:2992]};
      mid_1[1] = {1'b0,layer_2_1[3007:3000]} - {1'b0, layer_1_1[3007:3000]};
      mid_1[2] = {1'b0,layer_2_1[3015:3008]} - {1'b0, layer_1_1[3015:3008]};
      mid_2[0] = {1'b0,layer_2_2[2999:2992]} - {1'b0, layer_1_2[2999:2992]};
      mid_2[1] = {1'b0,layer_2_2[3007:3000]} - {1'b0, layer_1_2[3007:3000]};
      mid_2[2] = {1'b0,layer_2_2[3015:3008]} - {1'b0, layer_1_2[3015:3008]};
      btm_0[0] = {1'b0,layer_3_0[2999:2992]} - {1'b0, layer_2_0[2999:2992]};
      btm_0[1] = {1'b0,layer_3_0[3007:3000]} - {1'b0, layer_2_0[3007:3000]};
      btm_0[2] = {1'b0,layer_3_0[3015:3008]} - {1'b0, layer_2_0[3015:3008]};
      btm_1[0] = {1'b0,layer_3_1[2999:2992]} - {1'b0, layer_2_1[2999:2992]};
      btm_1[1] = {1'b0,layer_3_1[3007:3000]} - {1'b0, layer_2_1[3007:3000]};
      btm_1[2] = {1'b0,layer_3_1[3015:3008]} - {1'b0, layer_2_1[3015:3008]};
      btm_2[0] = {1'b0,layer_3_2[2999:2992]} - {1'b0, layer_2_2[2999:2992]};
      btm_2[1] = {1'b0,layer_3_2[3007:3000]} - {1'b0, layer_2_2[3007:3000]};
      btm_2[2] = {1'b0,layer_3_2[3015:3008]} - {1'b0, layer_2_2[3015:3008]};
    end
    'd376: begin
      top_0[0] = {1'b0,layer_1_0[3007:3000]} - {1'b0, layer_0_0[3007:3000]};
      top_0[1] = {1'b0,layer_1_0[3015:3008]} - {1'b0, layer_0_0[3015:3008]};
      top_0[2] = {1'b0,layer_1_0[3023:3016]} - {1'b0, layer_0_0[3023:3016]};
      top_1[0] = {1'b0,layer_1_1[3007:3000]} - {1'b0, layer_0_1[3007:3000]};
      top_1[1] = {1'b0,layer_1_1[3015:3008]} - {1'b0, layer_0_1[3015:3008]};
      top_1[2] = {1'b0,layer_1_1[3023:3016]} - {1'b0, layer_0_1[3023:3016]};
      top_2[0] = {1'b0,layer_1_2[3007:3000]} - {1'b0, layer_0_2[3007:3000]};
      top_2[1] = {1'b0,layer_1_2[3015:3008]} - {1'b0, layer_0_2[3015:3008]};
      top_2[2] = {1'b0,layer_1_2[3023:3016]} - {1'b0, layer_0_2[3023:3016]};
      mid_0[0] = {1'b0,layer_2_0[3007:3000]} - {1'b0, layer_1_0[3007:3000]};
      mid_0[1] = {1'b0,layer_2_0[3015:3008]} - {1'b0, layer_1_0[3015:3008]};
      mid_0[2] = {1'b0,layer_2_0[3023:3016]} - {1'b0, layer_1_0[3023:3016]};
      mid_1[0] = {1'b0,layer_2_1[3007:3000]} - {1'b0, layer_1_1[3007:3000]};
      mid_1[1] = {1'b0,layer_2_1[3015:3008]} - {1'b0, layer_1_1[3015:3008]};
      mid_1[2] = {1'b0,layer_2_1[3023:3016]} - {1'b0, layer_1_1[3023:3016]};
      mid_2[0] = {1'b0,layer_2_2[3007:3000]} - {1'b0, layer_1_2[3007:3000]};
      mid_2[1] = {1'b0,layer_2_2[3015:3008]} - {1'b0, layer_1_2[3015:3008]};
      mid_2[2] = {1'b0,layer_2_2[3023:3016]} - {1'b0, layer_1_2[3023:3016]};
      btm_0[0] = {1'b0,layer_3_0[3007:3000]} - {1'b0, layer_2_0[3007:3000]};
      btm_0[1] = {1'b0,layer_3_0[3015:3008]} - {1'b0, layer_2_0[3015:3008]};
      btm_0[2] = {1'b0,layer_3_0[3023:3016]} - {1'b0, layer_2_0[3023:3016]};
      btm_1[0] = {1'b0,layer_3_1[3007:3000]} - {1'b0, layer_2_1[3007:3000]};
      btm_1[1] = {1'b0,layer_3_1[3015:3008]} - {1'b0, layer_2_1[3015:3008]};
      btm_1[2] = {1'b0,layer_3_1[3023:3016]} - {1'b0, layer_2_1[3023:3016]};
      btm_2[0] = {1'b0,layer_3_2[3007:3000]} - {1'b0, layer_2_2[3007:3000]};
      btm_2[1] = {1'b0,layer_3_2[3015:3008]} - {1'b0, layer_2_2[3015:3008]};
      btm_2[2] = {1'b0,layer_3_2[3023:3016]} - {1'b0, layer_2_2[3023:3016]};
    end
    'd377: begin
      top_0[0] = {1'b0,layer_1_0[3015:3008]} - {1'b0, layer_0_0[3015:3008]};
      top_0[1] = {1'b0,layer_1_0[3023:3016]} - {1'b0, layer_0_0[3023:3016]};
      top_0[2] = {1'b0,layer_1_0[3031:3024]} - {1'b0, layer_0_0[3031:3024]};
      top_1[0] = {1'b0,layer_1_1[3015:3008]} - {1'b0, layer_0_1[3015:3008]};
      top_1[1] = {1'b0,layer_1_1[3023:3016]} - {1'b0, layer_0_1[3023:3016]};
      top_1[2] = {1'b0,layer_1_1[3031:3024]} - {1'b0, layer_0_1[3031:3024]};
      top_2[0] = {1'b0,layer_1_2[3015:3008]} - {1'b0, layer_0_2[3015:3008]};
      top_2[1] = {1'b0,layer_1_2[3023:3016]} - {1'b0, layer_0_2[3023:3016]};
      top_2[2] = {1'b0,layer_1_2[3031:3024]} - {1'b0, layer_0_2[3031:3024]};
      mid_0[0] = {1'b0,layer_2_0[3015:3008]} - {1'b0, layer_1_0[3015:3008]};
      mid_0[1] = {1'b0,layer_2_0[3023:3016]} - {1'b0, layer_1_0[3023:3016]};
      mid_0[2] = {1'b0,layer_2_0[3031:3024]} - {1'b0, layer_1_0[3031:3024]};
      mid_1[0] = {1'b0,layer_2_1[3015:3008]} - {1'b0, layer_1_1[3015:3008]};
      mid_1[1] = {1'b0,layer_2_1[3023:3016]} - {1'b0, layer_1_1[3023:3016]};
      mid_1[2] = {1'b0,layer_2_1[3031:3024]} - {1'b0, layer_1_1[3031:3024]};
      mid_2[0] = {1'b0,layer_2_2[3015:3008]} - {1'b0, layer_1_2[3015:3008]};
      mid_2[1] = {1'b0,layer_2_2[3023:3016]} - {1'b0, layer_1_2[3023:3016]};
      mid_2[2] = {1'b0,layer_2_2[3031:3024]} - {1'b0, layer_1_2[3031:3024]};
      btm_0[0] = {1'b0,layer_3_0[3015:3008]} - {1'b0, layer_2_0[3015:3008]};
      btm_0[1] = {1'b0,layer_3_0[3023:3016]} - {1'b0, layer_2_0[3023:3016]};
      btm_0[2] = {1'b0,layer_3_0[3031:3024]} - {1'b0, layer_2_0[3031:3024]};
      btm_1[0] = {1'b0,layer_3_1[3015:3008]} - {1'b0, layer_2_1[3015:3008]};
      btm_1[1] = {1'b0,layer_3_1[3023:3016]} - {1'b0, layer_2_1[3023:3016]};
      btm_1[2] = {1'b0,layer_3_1[3031:3024]} - {1'b0, layer_2_1[3031:3024]};
      btm_2[0] = {1'b0,layer_3_2[3015:3008]} - {1'b0, layer_2_2[3015:3008]};
      btm_2[1] = {1'b0,layer_3_2[3023:3016]} - {1'b0, layer_2_2[3023:3016]};
      btm_2[2] = {1'b0,layer_3_2[3031:3024]} - {1'b0, layer_2_2[3031:3024]};
    end
    'd378: begin
      top_0[0] = {1'b0,layer_1_0[3023:3016]} - {1'b0, layer_0_0[3023:3016]};
      top_0[1] = {1'b0,layer_1_0[3031:3024]} - {1'b0, layer_0_0[3031:3024]};
      top_0[2] = {1'b0,layer_1_0[3039:3032]} - {1'b0, layer_0_0[3039:3032]};
      top_1[0] = {1'b0,layer_1_1[3023:3016]} - {1'b0, layer_0_1[3023:3016]};
      top_1[1] = {1'b0,layer_1_1[3031:3024]} - {1'b0, layer_0_1[3031:3024]};
      top_1[2] = {1'b0,layer_1_1[3039:3032]} - {1'b0, layer_0_1[3039:3032]};
      top_2[0] = {1'b0,layer_1_2[3023:3016]} - {1'b0, layer_0_2[3023:3016]};
      top_2[1] = {1'b0,layer_1_2[3031:3024]} - {1'b0, layer_0_2[3031:3024]};
      top_2[2] = {1'b0,layer_1_2[3039:3032]} - {1'b0, layer_0_2[3039:3032]};
      mid_0[0] = {1'b0,layer_2_0[3023:3016]} - {1'b0, layer_1_0[3023:3016]};
      mid_0[1] = {1'b0,layer_2_0[3031:3024]} - {1'b0, layer_1_0[3031:3024]};
      mid_0[2] = {1'b0,layer_2_0[3039:3032]} - {1'b0, layer_1_0[3039:3032]};
      mid_1[0] = {1'b0,layer_2_1[3023:3016]} - {1'b0, layer_1_1[3023:3016]};
      mid_1[1] = {1'b0,layer_2_1[3031:3024]} - {1'b0, layer_1_1[3031:3024]};
      mid_1[2] = {1'b0,layer_2_1[3039:3032]} - {1'b0, layer_1_1[3039:3032]};
      mid_2[0] = {1'b0,layer_2_2[3023:3016]} - {1'b0, layer_1_2[3023:3016]};
      mid_2[1] = {1'b0,layer_2_2[3031:3024]} - {1'b0, layer_1_2[3031:3024]};
      mid_2[2] = {1'b0,layer_2_2[3039:3032]} - {1'b0, layer_1_2[3039:3032]};
      btm_0[0] = {1'b0,layer_3_0[3023:3016]} - {1'b0, layer_2_0[3023:3016]};
      btm_0[1] = {1'b0,layer_3_0[3031:3024]} - {1'b0, layer_2_0[3031:3024]};
      btm_0[2] = {1'b0,layer_3_0[3039:3032]} - {1'b0, layer_2_0[3039:3032]};
      btm_1[0] = {1'b0,layer_3_1[3023:3016]} - {1'b0, layer_2_1[3023:3016]};
      btm_1[1] = {1'b0,layer_3_1[3031:3024]} - {1'b0, layer_2_1[3031:3024]};
      btm_1[2] = {1'b0,layer_3_1[3039:3032]} - {1'b0, layer_2_1[3039:3032]};
      btm_2[0] = {1'b0,layer_3_2[3023:3016]} - {1'b0, layer_2_2[3023:3016]};
      btm_2[1] = {1'b0,layer_3_2[3031:3024]} - {1'b0, layer_2_2[3031:3024]};
      btm_2[2] = {1'b0,layer_3_2[3039:3032]} - {1'b0, layer_2_2[3039:3032]};
    end
    'd379: begin
      top_0[0] = {1'b0,layer_1_0[3031:3024]} - {1'b0, layer_0_0[3031:3024]};
      top_0[1] = {1'b0,layer_1_0[3039:3032]} - {1'b0, layer_0_0[3039:3032]};
      top_0[2] = {1'b0,layer_1_0[3047:3040]} - {1'b0, layer_0_0[3047:3040]};
      top_1[0] = {1'b0,layer_1_1[3031:3024]} - {1'b0, layer_0_1[3031:3024]};
      top_1[1] = {1'b0,layer_1_1[3039:3032]} - {1'b0, layer_0_1[3039:3032]};
      top_1[2] = {1'b0,layer_1_1[3047:3040]} - {1'b0, layer_0_1[3047:3040]};
      top_2[0] = {1'b0,layer_1_2[3031:3024]} - {1'b0, layer_0_2[3031:3024]};
      top_2[1] = {1'b0,layer_1_2[3039:3032]} - {1'b0, layer_0_2[3039:3032]};
      top_2[2] = {1'b0,layer_1_2[3047:3040]} - {1'b0, layer_0_2[3047:3040]};
      mid_0[0] = {1'b0,layer_2_0[3031:3024]} - {1'b0, layer_1_0[3031:3024]};
      mid_0[1] = {1'b0,layer_2_0[3039:3032]} - {1'b0, layer_1_0[3039:3032]};
      mid_0[2] = {1'b0,layer_2_0[3047:3040]} - {1'b0, layer_1_0[3047:3040]};
      mid_1[0] = {1'b0,layer_2_1[3031:3024]} - {1'b0, layer_1_1[3031:3024]};
      mid_1[1] = {1'b0,layer_2_1[3039:3032]} - {1'b0, layer_1_1[3039:3032]};
      mid_1[2] = {1'b0,layer_2_1[3047:3040]} - {1'b0, layer_1_1[3047:3040]};
      mid_2[0] = {1'b0,layer_2_2[3031:3024]} - {1'b0, layer_1_2[3031:3024]};
      mid_2[1] = {1'b0,layer_2_2[3039:3032]} - {1'b0, layer_1_2[3039:3032]};
      mid_2[2] = {1'b0,layer_2_2[3047:3040]} - {1'b0, layer_1_2[3047:3040]};
      btm_0[0] = {1'b0,layer_3_0[3031:3024]} - {1'b0, layer_2_0[3031:3024]};
      btm_0[1] = {1'b0,layer_3_0[3039:3032]} - {1'b0, layer_2_0[3039:3032]};
      btm_0[2] = {1'b0,layer_3_0[3047:3040]} - {1'b0, layer_2_0[3047:3040]};
      btm_1[0] = {1'b0,layer_3_1[3031:3024]} - {1'b0, layer_2_1[3031:3024]};
      btm_1[1] = {1'b0,layer_3_1[3039:3032]} - {1'b0, layer_2_1[3039:3032]};
      btm_1[2] = {1'b0,layer_3_1[3047:3040]} - {1'b0, layer_2_1[3047:3040]};
      btm_2[0] = {1'b0,layer_3_2[3031:3024]} - {1'b0, layer_2_2[3031:3024]};
      btm_2[1] = {1'b0,layer_3_2[3039:3032]} - {1'b0, layer_2_2[3039:3032]};
      btm_2[2] = {1'b0,layer_3_2[3047:3040]} - {1'b0, layer_2_2[3047:3040]};
    end
    'd380: begin
      top_0[0] = {1'b0,layer_1_0[3039:3032]} - {1'b0, layer_0_0[3039:3032]};
      top_0[1] = {1'b0,layer_1_0[3047:3040]} - {1'b0, layer_0_0[3047:3040]};
      top_0[2] = {1'b0,layer_1_0[3055:3048]} - {1'b0, layer_0_0[3055:3048]};
      top_1[0] = {1'b0,layer_1_1[3039:3032]} - {1'b0, layer_0_1[3039:3032]};
      top_1[1] = {1'b0,layer_1_1[3047:3040]} - {1'b0, layer_0_1[3047:3040]};
      top_1[2] = {1'b0,layer_1_1[3055:3048]} - {1'b0, layer_0_1[3055:3048]};
      top_2[0] = {1'b0,layer_1_2[3039:3032]} - {1'b0, layer_0_2[3039:3032]};
      top_2[1] = {1'b0,layer_1_2[3047:3040]} - {1'b0, layer_0_2[3047:3040]};
      top_2[2] = {1'b0,layer_1_2[3055:3048]} - {1'b0, layer_0_2[3055:3048]};
      mid_0[0] = {1'b0,layer_2_0[3039:3032]} - {1'b0, layer_1_0[3039:3032]};
      mid_0[1] = {1'b0,layer_2_0[3047:3040]} - {1'b0, layer_1_0[3047:3040]};
      mid_0[2] = {1'b0,layer_2_0[3055:3048]} - {1'b0, layer_1_0[3055:3048]};
      mid_1[0] = {1'b0,layer_2_1[3039:3032]} - {1'b0, layer_1_1[3039:3032]};
      mid_1[1] = {1'b0,layer_2_1[3047:3040]} - {1'b0, layer_1_1[3047:3040]};
      mid_1[2] = {1'b0,layer_2_1[3055:3048]} - {1'b0, layer_1_1[3055:3048]};
      mid_2[0] = {1'b0,layer_2_2[3039:3032]} - {1'b0, layer_1_2[3039:3032]};
      mid_2[1] = {1'b0,layer_2_2[3047:3040]} - {1'b0, layer_1_2[3047:3040]};
      mid_2[2] = {1'b0,layer_2_2[3055:3048]} - {1'b0, layer_1_2[3055:3048]};
      btm_0[0] = {1'b0,layer_3_0[3039:3032]} - {1'b0, layer_2_0[3039:3032]};
      btm_0[1] = {1'b0,layer_3_0[3047:3040]} - {1'b0, layer_2_0[3047:3040]};
      btm_0[2] = {1'b0,layer_3_0[3055:3048]} - {1'b0, layer_2_0[3055:3048]};
      btm_1[0] = {1'b0,layer_3_1[3039:3032]} - {1'b0, layer_2_1[3039:3032]};
      btm_1[1] = {1'b0,layer_3_1[3047:3040]} - {1'b0, layer_2_1[3047:3040]};
      btm_1[2] = {1'b0,layer_3_1[3055:3048]} - {1'b0, layer_2_1[3055:3048]};
      btm_2[0] = {1'b0,layer_3_2[3039:3032]} - {1'b0, layer_2_2[3039:3032]};
      btm_2[1] = {1'b0,layer_3_2[3047:3040]} - {1'b0, layer_2_2[3047:3040]};
      btm_2[2] = {1'b0,layer_3_2[3055:3048]} - {1'b0, layer_2_2[3055:3048]};
    end
    'd381: begin
      top_0[0] = {1'b0,layer_1_0[3047:3040]} - {1'b0, layer_0_0[3047:3040]};
      top_0[1] = {1'b0,layer_1_0[3055:3048]} - {1'b0, layer_0_0[3055:3048]};
      top_0[2] = {1'b0,layer_1_0[3063:3056]} - {1'b0, layer_0_0[3063:3056]};
      top_1[0] = {1'b0,layer_1_1[3047:3040]} - {1'b0, layer_0_1[3047:3040]};
      top_1[1] = {1'b0,layer_1_1[3055:3048]} - {1'b0, layer_0_1[3055:3048]};
      top_1[2] = {1'b0,layer_1_1[3063:3056]} - {1'b0, layer_0_1[3063:3056]};
      top_2[0] = {1'b0,layer_1_2[3047:3040]} - {1'b0, layer_0_2[3047:3040]};
      top_2[1] = {1'b0,layer_1_2[3055:3048]} - {1'b0, layer_0_2[3055:3048]};
      top_2[2] = {1'b0,layer_1_2[3063:3056]} - {1'b0, layer_0_2[3063:3056]};
      mid_0[0] = {1'b0,layer_2_0[3047:3040]} - {1'b0, layer_1_0[3047:3040]};
      mid_0[1] = {1'b0,layer_2_0[3055:3048]} - {1'b0, layer_1_0[3055:3048]};
      mid_0[2] = {1'b0,layer_2_0[3063:3056]} - {1'b0, layer_1_0[3063:3056]};
      mid_1[0] = {1'b0,layer_2_1[3047:3040]} - {1'b0, layer_1_1[3047:3040]};
      mid_1[1] = {1'b0,layer_2_1[3055:3048]} - {1'b0, layer_1_1[3055:3048]};
      mid_1[2] = {1'b0,layer_2_1[3063:3056]} - {1'b0, layer_1_1[3063:3056]};
      mid_2[0] = {1'b0,layer_2_2[3047:3040]} - {1'b0, layer_1_2[3047:3040]};
      mid_2[1] = {1'b0,layer_2_2[3055:3048]} - {1'b0, layer_1_2[3055:3048]};
      mid_2[2] = {1'b0,layer_2_2[3063:3056]} - {1'b0, layer_1_2[3063:3056]};
      btm_0[0] = {1'b0,layer_3_0[3047:3040]} - {1'b0, layer_2_0[3047:3040]};
      btm_0[1] = {1'b0,layer_3_0[3055:3048]} - {1'b0, layer_2_0[3055:3048]};
      btm_0[2] = {1'b0,layer_3_0[3063:3056]} - {1'b0, layer_2_0[3063:3056]};
      btm_1[0] = {1'b0,layer_3_1[3047:3040]} - {1'b0, layer_2_1[3047:3040]};
      btm_1[1] = {1'b0,layer_3_1[3055:3048]} - {1'b0, layer_2_1[3055:3048]};
      btm_1[2] = {1'b0,layer_3_1[3063:3056]} - {1'b0, layer_2_1[3063:3056]};
      btm_2[0] = {1'b0,layer_3_2[3047:3040]} - {1'b0, layer_2_2[3047:3040]};
      btm_2[1] = {1'b0,layer_3_2[3055:3048]} - {1'b0, layer_2_2[3055:3048]};
      btm_2[2] = {1'b0,layer_3_2[3063:3056]} - {1'b0, layer_2_2[3063:3056]};
    end
    'd382: begin
      top_0[0] = {1'b0,layer_1_0[3055:3048]} - {1'b0, layer_0_0[3055:3048]};
      top_0[1] = {1'b0,layer_1_0[3063:3056]} - {1'b0, layer_0_0[3063:3056]};
      top_0[2] = {1'b0,layer_1_0[3071:3064]} - {1'b0, layer_0_0[3071:3064]};
      top_1[0] = {1'b0,layer_1_1[3055:3048]} - {1'b0, layer_0_1[3055:3048]};
      top_1[1] = {1'b0,layer_1_1[3063:3056]} - {1'b0, layer_0_1[3063:3056]};
      top_1[2] = {1'b0,layer_1_1[3071:3064]} - {1'b0, layer_0_1[3071:3064]};
      top_2[0] = {1'b0,layer_1_2[3055:3048]} - {1'b0, layer_0_2[3055:3048]};
      top_2[1] = {1'b0,layer_1_2[3063:3056]} - {1'b0, layer_0_2[3063:3056]};
      top_2[2] = {1'b0,layer_1_2[3071:3064]} - {1'b0, layer_0_2[3071:3064]};
      mid_0[0] = {1'b0,layer_2_0[3055:3048]} - {1'b0, layer_1_0[3055:3048]};
      mid_0[1] = {1'b0,layer_2_0[3063:3056]} - {1'b0, layer_1_0[3063:3056]};
      mid_0[2] = {1'b0,layer_2_0[3071:3064]} - {1'b0, layer_1_0[3071:3064]};
      mid_1[0] = {1'b0,layer_2_1[3055:3048]} - {1'b0, layer_1_1[3055:3048]};
      mid_1[1] = {1'b0,layer_2_1[3063:3056]} - {1'b0, layer_1_1[3063:3056]};
      mid_1[2] = {1'b0,layer_2_1[3071:3064]} - {1'b0, layer_1_1[3071:3064]};
      mid_2[0] = {1'b0,layer_2_2[3055:3048]} - {1'b0, layer_1_2[3055:3048]};
      mid_2[1] = {1'b0,layer_2_2[3063:3056]} - {1'b0, layer_1_2[3063:3056]};
      mid_2[2] = {1'b0,layer_2_2[3071:3064]} - {1'b0, layer_1_2[3071:3064]};
      btm_0[0] = {1'b0,layer_3_0[3055:3048]} - {1'b0, layer_2_0[3055:3048]};
      btm_0[1] = {1'b0,layer_3_0[3063:3056]} - {1'b0, layer_2_0[3063:3056]};
      btm_0[2] = {1'b0,layer_3_0[3071:3064]} - {1'b0, layer_2_0[3071:3064]};
      btm_1[0] = {1'b0,layer_3_1[3055:3048]} - {1'b0, layer_2_1[3055:3048]};
      btm_1[1] = {1'b0,layer_3_1[3063:3056]} - {1'b0, layer_2_1[3063:3056]};
      btm_1[2] = {1'b0,layer_3_1[3071:3064]} - {1'b0, layer_2_1[3071:3064]};
      btm_2[0] = {1'b0,layer_3_2[3055:3048]} - {1'b0, layer_2_2[3055:3048]};
      btm_2[1] = {1'b0,layer_3_2[3063:3056]} - {1'b0, layer_2_2[3063:3056]};
      btm_2[2] = {1'b0,layer_3_2[3071:3064]} - {1'b0, layer_2_2[3071:3064]};
    end
    'd383: begin
      top_0[0] = {1'b0,layer_1_0[3063:3056]} - {1'b0, layer_0_0[3063:3056]};
      top_0[1] = {1'b0,layer_1_0[3071:3064]} - {1'b0, layer_0_0[3071:3064]};
      top_0[2] = {1'b0,layer_1_0[3079:3072]} - {1'b0, layer_0_0[3079:3072]};
      top_1[0] = {1'b0,layer_1_1[3063:3056]} - {1'b0, layer_0_1[3063:3056]};
      top_1[1] = {1'b0,layer_1_1[3071:3064]} - {1'b0, layer_0_1[3071:3064]};
      top_1[2] = {1'b0,layer_1_1[3079:3072]} - {1'b0, layer_0_1[3079:3072]};
      top_2[0] = {1'b0,layer_1_2[3063:3056]} - {1'b0, layer_0_2[3063:3056]};
      top_2[1] = {1'b0,layer_1_2[3071:3064]} - {1'b0, layer_0_2[3071:3064]};
      top_2[2] = {1'b0,layer_1_2[3079:3072]} - {1'b0, layer_0_2[3079:3072]};
      mid_0[0] = {1'b0,layer_2_0[3063:3056]} - {1'b0, layer_1_0[3063:3056]};
      mid_0[1] = {1'b0,layer_2_0[3071:3064]} - {1'b0, layer_1_0[3071:3064]};
      mid_0[2] = {1'b0,layer_2_0[3079:3072]} - {1'b0, layer_1_0[3079:3072]};
      mid_1[0] = {1'b0,layer_2_1[3063:3056]} - {1'b0, layer_1_1[3063:3056]};
      mid_1[1] = {1'b0,layer_2_1[3071:3064]} - {1'b0, layer_1_1[3071:3064]};
      mid_1[2] = {1'b0,layer_2_1[3079:3072]} - {1'b0, layer_1_1[3079:3072]};
      mid_2[0] = {1'b0,layer_2_2[3063:3056]} - {1'b0, layer_1_2[3063:3056]};
      mid_2[1] = {1'b0,layer_2_2[3071:3064]} - {1'b0, layer_1_2[3071:3064]};
      mid_2[2] = {1'b0,layer_2_2[3079:3072]} - {1'b0, layer_1_2[3079:3072]};
      btm_0[0] = {1'b0,layer_3_0[3063:3056]} - {1'b0, layer_2_0[3063:3056]};
      btm_0[1] = {1'b0,layer_3_0[3071:3064]} - {1'b0, layer_2_0[3071:3064]};
      btm_0[2] = {1'b0,layer_3_0[3079:3072]} - {1'b0, layer_2_0[3079:3072]};
      btm_1[0] = {1'b0,layer_3_1[3063:3056]} - {1'b0, layer_2_1[3063:3056]};
      btm_1[1] = {1'b0,layer_3_1[3071:3064]} - {1'b0, layer_2_1[3071:3064]};
      btm_1[2] = {1'b0,layer_3_1[3079:3072]} - {1'b0, layer_2_1[3079:3072]};
      btm_2[0] = {1'b0,layer_3_2[3063:3056]} - {1'b0, layer_2_2[3063:3056]};
      btm_2[1] = {1'b0,layer_3_2[3071:3064]} - {1'b0, layer_2_2[3071:3064]};
      btm_2[2] = {1'b0,layer_3_2[3079:3072]} - {1'b0, layer_2_2[3079:3072]};
    end
    'd384: begin
      top_0[0] = {1'b0,layer_1_0[3071:3064]} - {1'b0, layer_0_0[3071:3064]};
      top_0[1] = {1'b0,layer_1_0[3079:3072]} - {1'b0, layer_0_0[3079:3072]};
      top_0[2] = {1'b0,layer_1_0[3087:3080]} - {1'b0, layer_0_0[3087:3080]};
      top_1[0] = {1'b0,layer_1_1[3071:3064]} - {1'b0, layer_0_1[3071:3064]};
      top_1[1] = {1'b0,layer_1_1[3079:3072]} - {1'b0, layer_0_1[3079:3072]};
      top_1[2] = {1'b0,layer_1_1[3087:3080]} - {1'b0, layer_0_1[3087:3080]};
      top_2[0] = {1'b0,layer_1_2[3071:3064]} - {1'b0, layer_0_2[3071:3064]};
      top_2[1] = {1'b0,layer_1_2[3079:3072]} - {1'b0, layer_0_2[3079:3072]};
      top_2[2] = {1'b0,layer_1_2[3087:3080]} - {1'b0, layer_0_2[3087:3080]};
      mid_0[0] = {1'b0,layer_2_0[3071:3064]} - {1'b0, layer_1_0[3071:3064]};
      mid_0[1] = {1'b0,layer_2_0[3079:3072]} - {1'b0, layer_1_0[3079:3072]};
      mid_0[2] = {1'b0,layer_2_0[3087:3080]} - {1'b0, layer_1_0[3087:3080]};
      mid_1[0] = {1'b0,layer_2_1[3071:3064]} - {1'b0, layer_1_1[3071:3064]};
      mid_1[1] = {1'b0,layer_2_1[3079:3072]} - {1'b0, layer_1_1[3079:3072]};
      mid_1[2] = {1'b0,layer_2_1[3087:3080]} - {1'b0, layer_1_1[3087:3080]};
      mid_2[0] = {1'b0,layer_2_2[3071:3064]} - {1'b0, layer_1_2[3071:3064]};
      mid_2[1] = {1'b0,layer_2_2[3079:3072]} - {1'b0, layer_1_2[3079:3072]};
      mid_2[2] = {1'b0,layer_2_2[3087:3080]} - {1'b0, layer_1_2[3087:3080]};
      btm_0[0] = {1'b0,layer_3_0[3071:3064]} - {1'b0, layer_2_0[3071:3064]};
      btm_0[1] = {1'b0,layer_3_0[3079:3072]} - {1'b0, layer_2_0[3079:3072]};
      btm_0[2] = {1'b0,layer_3_0[3087:3080]} - {1'b0, layer_2_0[3087:3080]};
      btm_1[0] = {1'b0,layer_3_1[3071:3064]} - {1'b0, layer_2_1[3071:3064]};
      btm_1[1] = {1'b0,layer_3_1[3079:3072]} - {1'b0, layer_2_1[3079:3072]};
      btm_1[2] = {1'b0,layer_3_1[3087:3080]} - {1'b0, layer_2_1[3087:3080]};
      btm_2[0] = {1'b0,layer_3_2[3071:3064]} - {1'b0, layer_2_2[3071:3064]};
      btm_2[1] = {1'b0,layer_3_2[3079:3072]} - {1'b0, layer_2_2[3079:3072]};
      btm_2[2] = {1'b0,layer_3_2[3087:3080]} - {1'b0, layer_2_2[3087:3080]};
    end
    'd385: begin
      top_0[0] = {1'b0,layer_1_0[3079:3072]} - {1'b0, layer_0_0[3079:3072]};
      top_0[1] = {1'b0,layer_1_0[3087:3080]} - {1'b0, layer_0_0[3087:3080]};
      top_0[2] = {1'b0,layer_1_0[3095:3088]} - {1'b0, layer_0_0[3095:3088]};
      top_1[0] = {1'b0,layer_1_1[3079:3072]} - {1'b0, layer_0_1[3079:3072]};
      top_1[1] = {1'b0,layer_1_1[3087:3080]} - {1'b0, layer_0_1[3087:3080]};
      top_1[2] = {1'b0,layer_1_1[3095:3088]} - {1'b0, layer_0_1[3095:3088]};
      top_2[0] = {1'b0,layer_1_2[3079:3072]} - {1'b0, layer_0_2[3079:3072]};
      top_2[1] = {1'b0,layer_1_2[3087:3080]} - {1'b0, layer_0_2[3087:3080]};
      top_2[2] = {1'b0,layer_1_2[3095:3088]} - {1'b0, layer_0_2[3095:3088]};
      mid_0[0] = {1'b0,layer_2_0[3079:3072]} - {1'b0, layer_1_0[3079:3072]};
      mid_0[1] = {1'b0,layer_2_0[3087:3080]} - {1'b0, layer_1_0[3087:3080]};
      mid_0[2] = {1'b0,layer_2_0[3095:3088]} - {1'b0, layer_1_0[3095:3088]};
      mid_1[0] = {1'b0,layer_2_1[3079:3072]} - {1'b0, layer_1_1[3079:3072]};
      mid_1[1] = {1'b0,layer_2_1[3087:3080]} - {1'b0, layer_1_1[3087:3080]};
      mid_1[2] = {1'b0,layer_2_1[3095:3088]} - {1'b0, layer_1_1[3095:3088]};
      mid_2[0] = {1'b0,layer_2_2[3079:3072]} - {1'b0, layer_1_2[3079:3072]};
      mid_2[1] = {1'b0,layer_2_2[3087:3080]} - {1'b0, layer_1_2[3087:3080]};
      mid_2[2] = {1'b0,layer_2_2[3095:3088]} - {1'b0, layer_1_2[3095:3088]};
      btm_0[0] = {1'b0,layer_3_0[3079:3072]} - {1'b0, layer_2_0[3079:3072]};
      btm_0[1] = {1'b0,layer_3_0[3087:3080]} - {1'b0, layer_2_0[3087:3080]};
      btm_0[2] = {1'b0,layer_3_0[3095:3088]} - {1'b0, layer_2_0[3095:3088]};
      btm_1[0] = {1'b0,layer_3_1[3079:3072]} - {1'b0, layer_2_1[3079:3072]};
      btm_1[1] = {1'b0,layer_3_1[3087:3080]} - {1'b0, layer_2_1[3087:3080]};
      btm_1[2] = {1'b0,layer_3_1[3095:3088]} - {1'b0, layer_2_1[3095:3088]};
      btm_2[0] = {1'b0,layer_3_2[3079:3072]} - {1'b0, layer_2_2[3079:3072]};
      btm_2[1] = {1'b0,layer_3_2[3087:3080]} - {1'b0, layer_2_2[3087:3080]};
      btm_2[2] = {1'b0,layer_3_2[3095:3088]} - {1'b0, layer_2_2[3095:3088]};
    end
    'd386: begin
      top_0[0] = {1'b0,layer_1_0[3087:3080]} - {1'b0, layer_0_0[3087:3080]};
      top_0[1] = {1'b0,layer_1_0[3095:3088]} - {1'b0, layer_0_0[3095:3088]};
      top_0[2] = {1'b0,layer_1_0[3103:3096]} - {1'b0, layer_0_0[3103:3096]};
      top_1[0] = {1'b0,layer_1_1[3087:3080]} - {1'b0, layer_0_1[3087:3080]};
      top_1[1] = {1'b0,layer_1_1[3095:3088]} - {1'b0, layer_0_1[3095:3088]};
      top_1[2] = {1'b0,layer_1_1[3103:3096]} - {1'b0, layer_0_1[3103:3096]};
      top_2[0] = {1'b0,layer_1_2[3087:3080]} - {1'b0, layer_0_2[3087:3080]};
      top_2[1] = {1'b0,layer_1_2[3095:3088]} - {1'b0, layer_0_2[3095:3088]};
      top_2[2] = {1'b0,layer_1_2[3103:3096]} - {1'b0, layer_0_2[3103:3096]};
      mid_0[0] = {1'b0,layer_2_0[3087:3080]} - {1'b0, layer_1_0[3087:3080]};
      mid_0[1] = {1'b0,layer_2_0[3095:3088]} - {1'b0, layer_1_0[3095:3088]};
      mid_0[2] = {1'b0,layer_2_0[3103:3096]} - {1'b0, layer_1_0[3103:3096]};
      mid_1[0] = {1'b0,layer_2_1[3087:3080]} - {1'b0, layer_1_1[3087:3080]};
      mid_1[1] = {1'b0,layer_2_1[3095:3088]} - {1'b0, layer_1_1[3095:3088]};
      mid_1[2] = {1'b0,layer_2_1[3103:3096]} - {1'b0, layer_1_1[3103:3096]};
      mid_2[0] = {1'b0,layer_2_2[3087:3080]} - {1'b0, layer_1_2[3087:3080]};
      mid_2[1] = {1'b0,layer_2_2[3095:3088]} - {1'b0, layer_1_2[3095:3088]};
      mid_2[2] = {1'b0,layer_2_2[3103:3096]} - {1'b0, layer_1_2[3103:3096]};
      btm_0[0] = {1'b0,layer_3_0[3087:3080]} - {1'b0, layer_2_0[3087:3080]};
      btm_0[1] = {1'b0,layer_3_0[3095:3088]} - {1'b0, layer_2_0[3095:3088]};
      btm_0[2] = {1'b0,layer_3_0[3103:3096]} - {1'b0, layer_2_0[3103:3096]};
      btm_1[0] = {1'b0,layer_3_1[3087:3080]} - {1'b0, layer_2_1[3087:3080]};
      btm_1[1] = {1'b0,layer_3_1[3095:3088]} - {1'b0, layer_2_1[3095:3088]};
      btm_1[2] = {1'b0,layer_3_1[3103:3096]} - {1'b0, layer_2_1[3103:3096]};
      btm_2[0] = {1'b0,layer_3_2[3087:3080]} - {1'b0, layer_2_2[3087:3080]};
      btm_2[1] = {1'b0,layer_3_2[3095:3088]} - {1'b0, layer_2_2[3095:3088]};
      btm_2[2] = {1'b0,layer_3_2[3103:3096]} - {1'b0, layer_2_2[3103:3096]};
    end
    'd387: begin
      top_0[0] = {1'b0,layer_1_0[3095:3088]} - {1'b0, layer_0_0[3095:3088]};
      top_0[1] = {1'b0,layer_1_0[3103:3096]} - {1'b0, layer_0_0[3103:3096]};
      top_0[2] = {1'b0,layer_1_0[3111:3104]} - {1'b0, layer_0_0[3111:3104]};
      top_1[0] = {1'b0,layer_1_1[3095:3088]} - {1'b0, layer_0_1[3095:3088]};
      top_1[1] = {1'b0,layer_1_1[3103:3096]} - {1'b0, layer_0_1[3103:3096]};
      top_1[2] = {1'b0,layer_1_1[3111:3104]} - {1'b0, layer_0_1[3111:3104]};
      top_2[0] = {1'b0,layer_1_2[3095:3088]} - {1'b0, layer_0_2[3095:3088]};
      top_2[1] = {1'b0,layer_1_2[3103:3096]} - {1'b0, layer_0_2[3103:3096]};
      top_2[2] = {1'b0,layer_1_2[3111:3104]} - {1'b0, layer_0_2[3111:3104]};
      mid_0[0] = {1'b0,layer_2_0[3095:3088]} - {1'b0, layer_1_0[3095:3088]};
      mid_0[1] = {1'b0,layer_2_0[3103:3096]} - {1'b0, layer_1_0[3103:3096]};
      mid_0[2] = {1'b0,layer_2_0[3111:3104]} - {1'b0, layer_1_0[3111:3104]};
      mid_1[0] = {1'b0,layer_2_1[3095:3088]} - {1'b0, layer_1_1[3095:3088]};
      mid_1[1] = {1'b0,layer_2_1[3103:3096]} - {1'b0, layer_1_1[3103:3096]};
      mid_1[2] = {1'b0,layer_2_1[3111:3104]} - {1'b0, layer_1_1[3111:3104]};
      mid_2[0] = {1'b0,layer_2_2[3095:3088]} - {1'b0, layer_1_2[3095:3088]};
      mid_2[1] = {1'b0,layer_2_2[3103:3096]} - {1'b0, layer_1_2[3103:3096]};
      mid_2[2] = {1'b0,layer_2_2[3111:3104]} - {1'b0, layer_1_2[3111:3104]};
      btm_0[0] = {1'b0,layer_3_0[3095:3088]} - {1'b0, layer_2_0[3095:3088]};
      btm_0[1] = {1'b0,layer_3_0[3103:3096]} - {1'b0, layer_2_0[3103:3096]};
      btm_0[2] = {1'b0,layer_3_0[3111:3104]} - {1'b0, layer_2_0[3111:3104]};
      btm_1[0] = {1'b0,layer_3_1[3095:3088]} - {1'b0, layer_2_1[3095:3088]};
      btm_1[1] = {1'b0,layer_3_1[3103:3096]} - {1'b0, layer_2_1[3103:3096]};
      btm_1[2] = {1'b0,layer_3_1[3111:3104]} - {1'b0, layer_2_1[3111:3104]};
      btm_2[0] = {1'b0,layer_3_2[3095:3088]} - {1'b0, layer_2_2[3095:3088]};
      btm_2[1] = {1'b0,layer_3_2[3103:3096]} - {1'b0, layer_2_2[3103:3096]};
      btm_2[2] = {1'b0,layer_3_2[3111:3104]} - {1'b0, layer_2_2[3111:3104]};
    end
    'd388: begin
      top_0[0] = {1'b0,layer_1_0[3103:3096]} - {1'b0, layer_0_0[3103:3096]};
      top_0[1] = {1'b0,layer_1_0[3111:3104]} - {1'b0, layer_0_0[3111:3104]};
      top_0[2] = {1'b0,layer_1_0[3119:3112]} - {1'b0, layer_0_0[3119:3112]};
      top_1[0] = {1'b0,layer_1_1[3103:3096]} - {1'b0, layer_0_1[3103:3096]};
      top_1[1] = {1'b0,layer_1_1[3111:3104]} - {1'b0, layer_0_1[3111:3104]};
      top_1[2] = {1'b0,layer_1_1[3119:3112]} - {1'b0, layer_0_1[3119:3112]};
      top_2[0] = {1'b0,layer_1_2[3103:3096]} - {1'b0, layer_0_2[3103:3096]};
      top_2[1] = {1'b0,layer_1_2[3111:3104]} - {1'b0, layer_0_2[3111:3104]};
      top_2[2] = {1'b0,layer_1_2[3119:3112]} - {1'b0, layer_0_2[3119:3112]};
      mid_0[0] = {1'b0,layer_2_0[3103:3096]} - {1'b0, layer_1_0[3103:3096]};
      mid_0[1] = {1'b0,layer_2_0[3111:3104]} - {1'b0, layer_1_0[3111:3104]};
      mid_0[2] = {1'b0,layer_2_0[3119:3112]} - {1'b0, layer_1_0[3119:3112]};
      mid_1[0] = {1'b0,layer_2_1[3103:3096]} - {1'b0, layer_1_1[3103:3096]};
      mid_1[1] = {1'b0,layer_2_1[3111:3104]} - {1'b0, layer_1_1[3111:3104]};
      mid_1[2] = {1'b0,layer_2_1[3119:3112]} - {1'b0, layer_1_1[3119:3112]};
      mid_2[0] = {1'b0,layer_2_2[3103:3096]} - {1'b0, layer_1_2[3103:3096]};
      mid_2[1] = {1'b0,layer_2_2[3111:3104]} - {1'b0, layer_1_2[3111:3104]};
      mid_2[2] = {1'b0,layer_2_2[3119:3112]} - {1'b0, layer_1_2[3119:3112]};
      btm_0[0] = {1'b0,layer_3_0[3103:3096]} - {1'b0, layer_2_0[3103:3096]};
      btm_0[1] = {1'b0,layer_3_0[3111:3104]} - {1'b0, layer_2_0[3111:3104]};
      btm_0[2] = {1'b0,layer_3_0[3119:3112]} - {1'b0, layer_2_0[3119:3112]};
      btm_1[0] = {1'b0,layer_3_1[3103:3096]} - {1'b0, layer_2_1[3103:3096]};
      btm_1[1] = {1'b0,layer_3_1[3111:3104]} - {1'b0, layer_2_1[3111:3104]};
      btm_1[2] = {1'b0,layer_3_1[3119:3112]} - {1'b0, layer_2_1[3119:3112]};
      btm_2[0] = {1'b0,layer_3_2[3103:3096]} - {1'b0, layer_2_2[3103:3096]};
      btm_2[1] = {1'b0,layer_3_2[3111:3104]} - {1'b0, layer_2_2[3111:3104]};
      btm_2[2] = {1'b0,layer_3_2[3119:3112]} - {1'b0, layer_2_2[3119:3112]};
    end
    'd389: begin
      top_0[0] = {1'b0,layer_1_0[3111:3104]} - {1'b0, layer_0_0[3111:3104]};
      top_0[1] = {1'b0,layer_1_0[3119:3112]} - {1'b0, layer_0_0[3119:3112]};
      top_0[2] = {1'b0,layer_1_0[3127:3120]} - {1'b0, layer_0_0[3127:3120]};
      top_1[0] = {1'b0,layer_1_1[3111:3104]} - {1'b0, layer_0_1[3111:3104]};
      top_1[1] = {1'b0,layer_1_1[3119:3112]} - {1'b0, layer_0_1[3119:3112]};
      top_1[2] = {1'b0,layer_1_1[3127:3120]} - {1'b0, layer_0_1[3127:3120]};
      top_2[0] = {1'b0,layer_1_2[3111:3104]} - {1'b0, layer_0_2[3111:3104]};
      top_2[1] = {1'b0,layer_1_2[3119:3112]} - {1'b0, layer_0_2[3119:3112]};
      top_2[2] = {1'b0,layer_1_2[3127:3120]} - {1'b0, layer_0_2[3127:3120]};
      mid_0[0] = {1'b0,layer_2_0[3111:3104]} - {1'b0, layer_1_0[3111:3104]};
      mid_0[1] = {1'b0,layer_2_0[3119:3112]} - {1'b0, layer_1_0[3119:3112]};
      mid_0[2] = {1'b0,layer_2_0[3127:3120]} - {1'b0, layer_1_0[3127:3120]};
      mid_1[0] = {1'b0,layer_2_1[3111:3104]} - {1'b0, layer_1_1[3111:3104]};
      mid_1[1] = {1'b0,layer_2_1[3119:3112]} - {1'b0, layer_1_1[3119:3112]};
      mid_1[2] = {1'b0,layer_2_1[3127:3120]} - {1'b0, layer_1_1[3127:3120]};
      mid_2[0] = {1'b0,layer_2_2[3111:3104]} - {1'b0, layer_1_2[3111:3104]};
      mid_2[1] = {1'b0,layer_2_2[3119:3112]} - {1'b0, layer_1_2[3119:3112]};
      mid_2[2] = {1'b0,layer_2_2[3127:3120]} - {1'b0, layer_1_2[3127:3120]};
      btm_0[0] = {1'b0,layer_3_0[3111:3104]} - {1'b0, layer_2_0[3111:3104]};
      btm_0[1] = {1'b0,layer_3_0[3119:3112]} - {1'b0, layer_2_0[3119:3112]};
      btm_0[2] = {1'b0,layer_3_0[3127:3120]} - {1'b0, layer_2_0[3127:3120]};
      btm_1[0] = {1'b0,layer_3_1[3111:3104]} - {1'b0, layer_2_1[3111:3104]};
      btm_1[1] = {1'b0,layer_3_1[3119:3112]} - {1'b0, layer_2_1[3119:3112]};
      btm_1[2] = {1'b0,layer_3_1[3127:3120]} - {1'b0, layer_2_1[3127:3120]};
      btm_2[0] = {1'b0,layer_3_2[3111:3104]} - {1'b0, layer_2_2[3111:3104]};
      btm_2[1] = {1'b0,layer_3_2[3119:3112]} - {1'b0, layer_2_2[3119:3112]};
      btm_2[2] = {1'b0,layer_3_2[3127:3120]} - {1'b0, layer_2_2[3127:3120]};
    end
    'd390: begin
      top_0[0] = {1'b0,layer_1_0[3119:3112]} - {1'b0, layer_0_0[3119:3112]};
      top_0[1] = {1'b0,layer_1_0[3127:3120]} - {1'b0, layer_0_0[3127:3120]};
      top_0[2] = {1'b0,layer_1_0[3135:3128]} - {1'b0, layer_0_0[3135:3128]};
      top_1[0] = {1'b0,layer_1_1[3119:3112]} - {1'b0, layer_0_1[3119:3112]};
      top_1[1] = {1'b0,layer_1_1[3127:3120]} - {1'b0, layer_0_1[3127:3120]};
      top_1[2] = {1'b0,layer_1_1[3135:3128]} - {1'b0, layer_0_1[3135:3128]};
      top_2[0] = {1'b0,layer_1_2[3119:3112]} - {1'b0, layer_0_2[3119:3112]};
      top_2[1] = {1'b0,layer_1_2[3127:3120]} - {1'b0, layer_0_2[3127:3120]};
      top_2[2] = {1'b0,layer_1_2[3135:3128]} - {1'b0, layer_0_2[3135:3128]};
      mid_0[0] = {1'b0,layer_2_0[3119:3112]} - {1'b0, layer_1_0[3119:3112]};
      mid_0[1] = {1'b0,layer_2_0[3127:3120]} - {1'b0, layer_1_0[3127:3120]};
      mid_0[2] = {1'b0,layer_2_0[3135:3128]} - {1'b0, layer_1_0[3135:3128]};
      mid_1[0] = {1'b0,layer_2_1[3119:3112]} - {1'b0, layer_1_1[3119:3112]};
      mid_1[1] = {1'b0,layer_2_1[3127:3120]} - {1'b0, layer_1_1[3127:3120]};
      mid_1[2] = {1'b0,layer_2_1[3135:3128]} - {1'b0, layer_1_1[3135:3128]};
      mid_2[0] = {1'b0,layer_2_2[3119:3112]} - {1'b0, layer_1_2[3119:3112]};
      mid_2[1] = {1'b0,layer_2_2[3127:3120]} - {1'b0, layer_1_2[3127:3120]};
      mid_2[2] = {1'b0,layer_2_2[3135:3128]} - {1'b0, layer_1_2[3135:3128]};
      btm_0[0] = {1'b0,layer_3_0[3119:3112]} - {1'b0, layer_2_0[3119:3112]};
      btm_0[1] = {1'b0,layer_3_0[3127:3120]} - {1'b0, layer_2_0[3127:3120]};
      btm_0[2] = {1'b0,layer_3_0[3135:3128]} - {1'b0, layer_2_0[3135:3128]};
      btm_1[0] = {1'b0,layer_3_1[3119:3112]} - {1'b0, layer_2_1[3119:3112]};
      btm_1[1] = {1'b0,layer_3_1[3127:3120]} - {1'b0, layer_2_1[3127:3120]};
      btm_1[2] = {1'b0,layer_3_1[3135:3128]} - {1'b0, layer_2_1[3135:3128]};
      btm_2[0] = {1'b0,layer_3_2[3119:3112]} - {1'b0, layer_2_2[3119:3112]};
      btm_2[1] = {1'b0,layer_3_2[3127:3120]} - {1'b0, layer_2_2[3127:3120]};
      btm_2[2] = {1'b0,layer_3_2[3135:3128]} - {1'b0, layer_2_2[3135:3128]};
    end
    'd391: begin
      top_0[0] = {1'b0,layer_1_0[3127:3120]} - {1'b0, layer_0_0[3127:3120]};
      top_0[1] = {1'b0,layer_1_0[3135:3128]} - {1'b0, layer_0_0[3135:3128]};
      top_0[2] = {1'b0,layer_1_0[3143:3136]} - {1'b0, layer_0_0[3143:3136]};
      top_1[0] = {1'b0,layer_1_1[3127:3120]} - {1'b0, layer_0_1[3127:3120]};
      top_1[1] = {1'b0,layer_1_1[3135:3128]} - {1'b0, layer_0_1[3135:3128]};
      top_1[2] = {1'b0,layer_1_1[3143:3136]} - {1'b0, layer_0_1[3143:3136]};
      top_2[0] = {1'b0,layer_1_2[3127:3120]} - {1'b0, layer_0_2[3127:3120]};
      top_2[1] = {1'b0,layer_1_2[3135:3128]} - {1'b0, layer_0_2[3135:3128]};
      top_2[2] = {1'b0,layer_1_2[3143:3136]} - {1'b0, layer_0_2[3143:3136]};
      mid_0[0] = {1'b0,layer_2_0[3127:3120]} - {1'b0, layer_1_0[3127:3120]};
      mid_0[1] = {1'b0,layer_2_0[3135:3128]} - {1'b0, layer_1_0[3135:3128]};
      mid_0[2] = {1'b0,layer_2_0[3143:3136]} - {1'b0, layer_1_0[3143:3136]};
      mid_1[0] = {1'b0,layer_2_1[3127:3120]} - {1'b0, layer_1_1[3127:3120]};
      mid_1[1] = {1'b0,layer_2_1[3135:3128]} - {1'b0, layer_1_1[3135:3128]};
      mid_1[2] = {1'b0,layer_2_1[3143:3136]} - {1'b0, layer_1_1[3143:3136]};
      mid_2[0] = {1'b0,layer_2_2[3127:3120]} - {1'b0, layer_1_2[3127:3120]};
      mid_2[1] = {1'b0,layer_2_2[3135:3128]} - {1'b0, layer_1_2[3135:3128]};
      mid_2[2] = {1'b0,layer_2_2[3143:3136]} - {1'b0, layer_1_2[3143:3136]};
      btm_0[0] = {1'b0,layer_3_0[3127:3120]} - {1'b0, layer_2_0[3127:3120]};
      btm_0[1] = {1'b0,layer_3_0[3135:3128]} - {1'b0, layer_2_0[3135:3128]};
      btm_0[2] = {1'b0,layer_3_0[3143:3136]} - {1'b0, layer_2_0[3143:3136]};
      btm_1[0] = {1'b0,layer_3_1[3127:3120]} - {1'b0, layer_2_1[3127:3120]};
      btm_1[1] = {1'b0,layer_3_1[3135:3128]} - {1'b0, layer_2_1[3135:3128]};
      btm_1[2] = {1'b0,layer_3_1[3143:3136]} - {1'b0, layer_2_1[3143:3136]};
      btm_2[0] = {1'b0,layer_3_2[3127:3120]} - {1'b0, layer_2_2[3127:3120]};
      btm_2[1] = {1'b0,layer_3_2[3135:3128]} - {1'b0, layer_2_2[3135:3128]};
      btm_2[2] = {1'b0,layer_3_2[3143:3136]} - {1'b0, layer_2_2[3143:3136]};
    end
    'd392: begin
      top_0[0] = {1'b0,layer_1_0[3135:3128]} - {1'b0, layer_0_0[3135:3128]};
      top_0[1] = {1'b0,layer_1_0[3143:3136]} - {1'b0, layer_0_0[3143:3136]};
      top_0[2] = {1'b0,layer_1_0[3151:3144]} - {1'b0, layer_0_0[3151:3144]};
      top_1[0] = {1'b0,layer_1_1[3135:3128]} - {1'b0, layer_0_1[3135:3128]};
      top_1[1] = {1'b0,layer_1_1[3143:3136]} - {1'b0, layer_0_1[3143:3136]};
      top_1[2] = {1'b0,layer_1_1[3151:3144]} - {1'b0, layer_0_1[3151:3144]};
      top_2[0] = {1'b0,layer_1_2[3135:3128]} - {1'b0, layer_0_2[3135:3128]};
      top_2[1] = {1'b0,layer_1_2[3143:3136]} - {1'b0, layer_0_2[3143:3136]};
      top_2[2] = {1'b0,layer_1_2[3151:3144]} - {1'b0, layer_0_2[3151:3144]};
      mid_0[0] = {1'b0,layer_2_0[3135:3128]} - {1'b0, layer_1_0[3135:3128]};
      mid_0[1] = {1'b0,layer_2_0[3143:3136]} - {1'b0, layer_1_0[3143:3136]};
      mid_0[2] = {1'b0,layer_2_0[3151:3144]} - {1'b0, layer_1_0[3151:3144]};
      mid_1[0] = {1'b0,layer_2_1[3135:3128]} - {1'b0, layer_1_1[3135:3128]};
      mid_1[1] = {1'b0,layer_2_1[3143:3136]} - {1'b0, layer_1_1[3143:3136]};
      mid_1[2] = {1'b0,layer_2_1[3151:3144]} - {1'b0, layer_1_1[3151:3144]};
      mid_2[0] = {1'b0,layer_2_2[3135:3128]} - {1'b0, layer_1_2[3135:3128]};
      mid_2[1] = {1'b0,layer_2_2[3143:3136]} - {1'b0, layer_1_2[3143:3136]};
      mid_2[2] = {1'b0,layer_2_2[3151:3144]} - {1'b0, layer_1_2[3151:3144]};
      btm_0[0] = {1'b0,layer_3_0[3135:3128]} - {1'b0, layer_2_0[3135:3128]};
      btm_0[1] = {1'b0,layer_3_0[3143:3136]} - {1'b0, layer_2_0[3143:3136]};
      btm_0[2] = {1'b0,layer_3_0[3151:3144]} - {1'b0, layer_2_0[3151:3144]};
      btm_1[0] = {1'b0,layer_3_1[3135:3128]} - {1'b0, layer_2_1[3135:3128]};
      btm_1[1] = {1'b0,layer_3_1[3143:3136]} - {1'b0, layer_2_1[3143:3136]};
      btm_1[2] = {1'b0,layer_3_1[3151:3144]} - {1'b0, layer_2_1[3151:3144]};
      btm_2[0] = {1'b0,layer_3_2[3135:3128]} - {1'b0, layer_2_2[3135:3128]};
      btm_2[1] = {1'b0,layer_3_2[3143:3136]} - {1'b0, layer_2_2[3143:3136]};
      btm_2[2] = {1'b0,layer_3_2[3151:3144]} - {1'b0, layer_2_2[3151:3144]};
    end
    'd393: begin
      top_0[0] = {1'b0,layer_1_0[3143:3136]} - {1'b0, layer_0_0[3143:3136]};
      top_0[1] = {1'b0,layer_1_0[3151:3144]} - {1'b0, layer_0_0[3151:3144]};
      top_0[2] = {1'b0,layer_1_0[3159:3152]} - {1'b0, layer_0_0[3159:3152]};
      top_1[0] = {1'b0,layer_1_1[3143:3136]} - {1'b0, layer_0_1[3143:3136]};
      top_1[1] = {1'b0,layer_1_1[3151:3144]} - {1'b0, layer_0_1[3151:3144]};
      top_1[2] = {1'b0,layer_1_1[3159:3152]} - {1'b0, layer_0_1[3159:3152]};
      top_2[0] = {1'b0,layer_1_2[3143:3136]} - {1'b0, layer_0_2[3143:3136]};
      top_2[1] = {1'b0,layer_1_2[3151:3144]} - {1'b0, layer_0_2[3151:3144]};
      top_2[2] = {1'b0,layer_1_2[3159:3152]} - {1'b0, layer_0_2[3159:3152]};
      mid_0[0] = {1'b0,layer_2_0[3143:3136]} - {1'b0, layer_1_0[3143:3136]};
      mid_0[1] = {1'b0,layer_2_0[3151:3144]} - {1'b0, layer_1_0[3151:3144]};
      mid_0[2] = {1'b0,layer_2_0[3159:3152]} - {1'b0, layer_1_0[3159:3152]};
      mid_1[0] = {1'b0,layer_2_1[3143:3136]} - {1'b0, layer_1_1[3143:3136]};
      mid_1[1] = {1'b0,layer_2_1[3151:3144]} - {1'b0, layer_1_1[3151:3144]};
      mid_1[2] = {1'b0,layer_2_1[3159:3152]} - {1'b0, layer_1_1[3159:3152]};
      mid_2[0] = {1'b0,layer_2_2[3143:3136]} - {1'b0, layer_1_2[3143:3136]};
      mid_2[1] = {1'b0,layer_2_2[3151:3144]} - {1'b0, layer_1_2[3151:3144]};
      mid_2[2] = {1'b0,layer_2_2[3159:3152]} - {1'b0, layer_1_2[3159:3152]};
      btm_0[0] = {1'b0,layer_3_0[3143:3136]} - {1'b0, layer_2_0[3143:3136]};
      btm_0[1] = {1'b0,layer_3_0[3151:3144]} - {1'b0, layer_2_0[3151:3144]};
      btm_0[2] = {1'b0,layer_3_0[3159:3152]} - {1'b0, layer_2_0[3159:3152]};
      btm_1[0] = {1'b0,layer_3_1[3143:3136]} - {1'b0, layer_2_1[3143:3136]};
      btm_1[1] = {1'b0,layer_3_1[3151:3144]} - {1'b0, layer_2_1[3151:3144]};
      btm_1[2] = {1'b0,layer_3_1[3159:3152]} - {1'b0, layer_2_1[3159:3152]};
      btm_2[0] = {1'b0,layer_3_2[3143:3136]} - {1'b0, layer_2_2[3143:3136]};
      btm_2[1] = {1'b0,layer_3_2[3151:3144]} - {1'b0, layer_2_2[3151:3144]};
      btm_2[2] = {1'b0,layer_3_2[3159:3152]} - {1'b0, layer_2_2[3159:3152]};
    end
    'd394: begin
      top_0[0] = {1'b0,layer_1_0[3151:3144]} - {1'b0, layer_0_0[3151:3144]};
      top_0[1] = {1'b0,layer_1_0[3159:3152]} - {1'b0, layer_0_0[3159:3152]};
      top_0[2] = {1'b0,layer_1_0[3167:3160]} - {1'b0, layer_0_0[3167:3160]};
      top_1[0] = {1'b0,layer_1_1[3151:3144]} - {1'b0, layer_0_1[3151:3144]};
      top_1[1] = {1'b0,layer_1_1[3159:3152]} - {1'b0, layer_0_1[3159:3152]};
      top_1[2] = {1'b0,layer_1_1[3167:3160]} - {1'b0, layer_0_1[3167:3160]};
      top_2[0] = {1'b0,layer_1_2[3151:3144]} - {1'b0, layer_0_2[3151:3144]};
      top_2[1] = {1'b0,layer_1_2[3159:3152]} - {1'b0, layer_0_2[3159:3152]};
      top_2[2] = {1'b0,layer_1_2[3167:3160]} - {1'b0, layer_0_2[3167:3160]};
      mid_0[0] = {1'b0,layer_2_0[3151:3144]} - {1'b0, layer_1_0[3151:3144]};
      mid_0[1] = {1'b0,layer_2_0[3159:3152]} - {1'b0, layer_1_0[3159:3152]};
      mid_0[2] = {1'b0,layer_2_0[3167:3160]} - {1'b0, layer_1_0[3167:3160]};
      mid_1[0] = {1'b0,layer_2_1[3151:3144]} - {1'b0, layer_1_1[3151:3144]};
      mid_1[1] = {1'b0,layer_2_1[3159:3152]} - {1'b0, layer_1_1[3159:3152]};
      mid_1[2] = {1'b0,layer_2_1[3167:3160]} - {1'b0, layer_1_1[3167:3160]};
      mid_2[0] = {1'b0,layer_2_2[3151:3144]} - {1'b0, layer_1_2[3151:3144]};
      mid_2[1] = {1'b0,layer_2_2[3159:3152]} - {1'b0, layer_1_2[3159:3152]};
      mid_2[2] = {1'b0,layer_2_2[3167:3160]} - {1'b0, layer_1_2[3167:3160]};
      btm_0[0] = {1'b0,layer_3_0[3151:3144]} - {1'b0, layer_2_0[3151:3144]};
      btm_0[1] = {1'b0,layer_3_0[3159:3152]} - {1'b0, layer_2_0[3159:3152]};
      btm_0[2] = {1'b0,layer_3_0[3167:3160]} - {1'b0, layer_2_0[3167:3160]};
      btm_1[0] = {1'b0,layer_3_1[3151:3144]} - {1'b0, layer_2_1[3151:3144]};
      btm_1[1] = {1'b0,layer_3_1[3159:3152]} - {1'b0, layer_2_1[3159:3152]};
      btm_1[2] = {1'b0,layer_3_1[3167:3160]} - {1'b0, layer_2_1[3167:3160]};
      btm_2[0] = {1'b0,layer_3_2[3151:3144]} - {1'b0, layer_2_2[3151:3144]};
      btm_2[1] = {1'b0,layer_3_2[3159:3152]} - {1'b0, layer_2_2[3159:3152]};
      btm_2[2] = {1'b0,layer_3_2[3167:3160]} - {1'b0, layer_2_2[3167:3160]};
    end
    'd395: begin
      top_0[0] = {1'b0,layer_1_0[3159:3152]} - {1'b0, layer_0_0[3159:3152]};
      top_0[1] = {1'b0,layer_1_0[3167:3160]} - {1'b0, layer_0_0[3167:3160]};
      top_0[2] = {1'b0,layer_1_0[3175:3168]} - {1'b0, layer_0_0[3175:3168]};
      top_1[0] = {1'b0,layer_1_1[3159:3152]} - {1'b0, layer_0_1[3159:3152]};
      top_1[1] = {1'b0,layer_1_1[3167:3160]} - {1'b0, layer_0_1[3167:3160]};
      top_1[2] = {1'b0,layer_1_1[3175:3168]} - {1'b0, layer_0_1[3175:3168]};
      top_2[0] = {1'b0,layer_1_2[3159:3152]} - {1'b0, layer_0_2[3159:3152]};
      top_2[1] = {1'b0,layer_1_2[3167:3160]} - {1'b0, layer_0_2[3167:3160]};
      top_2[2] = {1'b0,layer_1_2[3175:3168]} - {1'b0, layer_0_2[3175:3168]};
      mid_0[0] = {1'b0,layer_2_0[3159:3152]} - {1'b0, layer_1_0[3159:3152]};
      mid_0[1] = {1'b0,layer_2_0[3167:3160]} - {1'b0, layer_1_0[3167:3160]};
      mid_0[2] = {1'b0,layer_2_0[3175:3168]} - {1'b0, layer_1_0[3175:3168]};
      mid_1[0] = {1'b0,layer_2_1[3159:3152]} - {1'b0, layer_1_1[3159:3152]};
      mid_1[1] = {1'b0,layer_2_1[3167:3160]} - {1'b0, layer_1_1[3167:3160]};
      mid_1[2] = {1'b0,layer_2_1[3175:3168]} - {1'b0, layer_1_1[3175:3168]};
      mid_2[0] = {1'b0,layer_2_2[3159:3152]} - {1'b0, layer_1_2[3159:3152]};
      mid_2[1] = {1'b0,layer_2_2[3167:3160]} - {1'b0, layer_1_2[3167:3160]};
      mid_2[2] = {1'b0,layer_2_2[3175:3168]} - {1'b0, layer_1_2[3175:3168]};
      btm_0[0] = {1'b0,layer_3_0[3159:3152]} - {1'b0, layer_2_0[3159:3152]};
      btm_0[1] = {1'b0,layer_3_0[3167:3160]} - {1'b0, layer_2_0[3167:3160]};
      btm_0[2] = {1'b0,layer_3_0[3175:3168]} - {1'b0, layer_2_0[3175:3168]};
      btm_1[0] = {1'b0,layer_3_1[3159:3152]} - {1'b0, layer_2_1[3159:3152]};
      btm_1[1] = {1'b0,layer_3_1[3167:3160]} - {1'b0, layer_2_1[3167:3160]};
      btm_1[2] = {1'b0,layer_3_1[3175:3168]} - {1'b0, layer_2_1[3175:3168]};
      btm_2[0] = {1'b0,layer_3_2[3159:3152]} - {1'b0, layer_2_2[3159:3152]};
      btm_2[1] = {1'b0,layer_3_2[3167:3160]} - {1'b0, layer_2_2[3167:3160]};
      btm_2[2] = {1'b0,layer_3_2[3175:3168]} - {1'b0, layer_2_2[3175:3168]};
    end
    'd396: begin
      top_0[0] = {1'b0,layer_1_0[3167:3160]} - {1'b0, layer_0_0[3167:3160]};
      top_0[1] = {1'b0,layer_1_0[3175:3168]} - {1'b0, layer_0_0[3175:3168]};
      top_0[2] = {1'b0,layer_1_0[3183:3176]} - {1'b0, layer_0_0[3183:3176]};
      top_1[0] = {1'b0,layer_1_1[3167:3160]} - {1'b0, layer_0_1[3167:3160]};
      top_1[1] = {1'b0,layer_1_1[3175:3168]} - {1'b0, layer_0_1[3175:3168]};
      top_1[2] = {1'b0,layer_1_1[3183:3176]} - {1'b0, layer_0_1[3183:3176]};
      top_2[0] = {1'b0,layer_1_2[3167:3160]} - {1'b0, layer_0_2[3167:3160]};
      top_2[1] = {1'b0,layer_1_2[3175:3168]} - {1'b0, layer_0_2[3175:3168]};
      top_2[2] = {1'b0,layer_1_2[3183:3176]} - {1'b0, layer_0_2[3183:3176]};
      mid_0[0] = {1'b0,layer_2_0[3167:3160]} - {1'b0, layer_1_0[3167:3160]};
      mid_0[1] = {1'b0,layer_2_0[3175:3168]} - {1'b0, layer_1_0[3175:3168]};
      mid_0[2] = {1'b0,layer_2_0[3183:3176]} - {1'b0, layer_1_0[3183:3176]};
      mid_1[0] = {1'b0,layer_2_1[3167:3160]} - {1'b0, layer_1_1[3167:3160]};
      mid_1[1] = {1'b0,layer_2_1[3175:3168]} - {1'b0, layer_1_1[3175:3168]};
      mid_1[2] = {1'b0,layer_2_1[3183:3176]} - {1'b0, layer_1_1[3183:3176]};
      mid_2[0] = {1'b0,layer_2_2[3167:3160]} - {1'b0, layer_1_2[3167:3160]};
      mid_2[1] = {1'b0,layer_2_2[3175:3168]} - {1'b0, layer_1_2[3175:3168]};
      mid_2[2] = {1'b0,layer_2_2[3183:3176]} - {1'b0, layer_1_2[3183:3176]};
      btm_0[0] = {1'b0,layer_3_0[3167:3160]} - {1'b0, layer_2_0[3167:3160]};
      btm_0[1] = {1'b0,layer_3_0[3175:3168]} - {1'b0, layer_2_0[3175:3168]};
      btm_0[2] = {1'b0,layer_3_0[3183:3176]} - {1'b0, layer_2_0[3183:3176]};
      btm_1[0] = {1'b0,layer_3_1[3167:3160]} - {1'b0, layer_2_1[3167:3160]};
      btm_1[1] = {1'b0,layer_3_1[3175:3168]} - {1'b0, layer_2_1[3175:3168]};
      btm_1[2] = {1'b0,layer_3_1[3183:3176]} - {1'b0, layer_2_1[3183:3176]};
      btm_2[0] = {1'b0,layer_3_2[3167:3160]} - {1'b0, layer_2_2[3167:3160]};
      btm_2[1] = {1'b0,layer_3_2[3175:3168]} - {1'b0, layer_2_2[3175:3168]};
      btm_2[2] = {1'b0,layer_3_2[3183:3176]} - {1'b0, layer_2_2[3183:3176]};
    end
    'd397: begin
      top_0[0] = {1'b0,layer_1_0[3175:3168]} - {1'b0, layer_0_0[3175:3168]};
      top_0[1] = {1'b0,layer_1_0[3183:3176]} - {1'b0, layer_0_0[3183:3176]};
      top_0[2] = {1'b0,layer_1_0[3191:3184]} - {1'b0, layer_0_0[3191:3184]};
      top_1[0] = {1'b0,layer_1_1[3175:3168]} - {1'b0, layer_0_1[3175:3168]};
      top_1[1] = {1'b0,layer_1_1[3183:3176]} - {1'b0, layer_0_1[3183:3176]};
      top_1[2] = {1'b0,layer_1_1[3191:3184]} - {1'b0, layer_0_1[3191:3184]};
      top_2[0] = {1'b0,layer_1_2[3175:3168]} - {1'b0, layer_0_2[3175:3168]};
      top_2[1] = {1'b0,layer_1_2[3183:3176]} - {1'b0, layer_0_2[3183:3176]};
      top_2[2] = {1'b0,layer_1_2[3191:3184]} - {1'b0, layer_0_2[3191:3184]};
      mid_0[0] = {1'b0,layer_2_0[3175:3168]} - {1'b0, layer_1_0[3175:3168]};
      mid_0[1] = {1'b0,layer_2_0[3183:3176]} - {1'b0, layer_1_0[3183:3176]};
      mid_0[2] = {1'b0,layer_2_0[3191:3184]} - {1'b0, layer_1_0[3191:3184]};
      mid_1[0] = {1'b0,layer_2_1[3175:3168]} - {1'b0, layer_1_1[3175:3168]};
      mid_1[1] = {1'b0,layer_2_1[3183:3176]} - {1'b0, layer_1_1[3183:3176]};
      mid_1[2] = {1'b0,layer_2_1[3191:3184]} - {1'b0, layer_1_1[3191:3184]};
      mid_2[0] = {1'b0,layer_2_2[3175:3168]} - {1'b0, layer_1_2[3175:3168]};
      mid_2[1] = {1'b0,layer_2_2[3183:3176]} - {1'b0, layer_1_2[3183:3176]};
      mid_2[2] = {1'b0,layer_2_2[3191:3184]} - {1'b0, layer_1_2[3191:3184]};
      btm_0[0] = {1'b0,layer_3_0[3175:3168]} - {1'b0, layer_2_0[3175:3168]};
      btm_0[1] = {1'b0,layer_3_0[3183:3176]} - {1'b0, layer_2_0[3183:3176]};
      btm_0[2] = {1'b0,layer_3_0[3191:3184]} - {1'b0, layer_2_0[3191:3184]};
      btm_1[0] = {1'b0,layer_3_1[3175:3168]} - {1'b0, layer_2_1[3175:3168]};
      btm_1[1] = {1'b0,layer_3_1[3183:3176]} - {1'b0, layer_2_1[3183:3176]};
      btm_1[2] = {1'b0,layer_3_1[3191:3184]} - {1'b0, layer_2_1[3191:3184]};
      btm_2[0] = {1'b0,layer_3_2[3175:3168]} - {1'b0, layer_2_2[3175:3168]};
      btm_2[1] = {1'b0,layer_3_2[3183:3176]} - {1'b0, layer_2_2[3183:3176]};
      btm_2[2] = {1'b0,layer_3_2[3191:3184]} - {1'b0, layer_2_2[3191:3184]};
    end
    'd398: begin
      top_0[0] = {1'b0,layer_1_0[3183:3176]} - {1'b0, layer_0_0[3183:3176]};
      top_0[1] = {1'b0,layer_1_0[3191:3184]} - {1'b0, layer_0_0[3191:3184]};
      top_0[2] = {1'b0,layer_1_0[3199:3192]} - {1'b0, layer_0_0[3199:3192]};
      top_1[0] = {1'b0,layer_1_1[3183:3176]} - {1'b0, layer_0_1[3183:3176]};
      top_1[1] = {1'b0,layer_1_1[3191:3184]} - {1'b0, layer_0_1[3191:3184]};
      top_1[2] = {1'b0,layer_1_1[3199:3192]} - {1'b0, layer_0_1[3199:3192]};
      top_2[0] = {1'b0,layer_1_2[3183:3176]} - {1'b0, layer_0_2[3183:3176]};
      top_2[1] = {1'b0,layer_1_2[3191:3184]} - {1'b0, layer_0_2[3191:3184]};
      top_2[2] = {1'b0,layer_1_2[3199:3192]} - {1'b0, layer_0_2[3199:3192]};
      mid_0[0] = {1'b0,layer_2_0[3183:3176]} - {1'b0, layer_1_0[3183:3176]};
      mid_0[1] = {1'b0,layer_2_0[3191:3184]} - {1'b0, layer_1_0[3191:3184]};
      mid_0[2] = {1'b0,layer_2_0[3199:3192]} - {1'b0, layer_1_0[3199:3192]};
      mid_1[0] = {1'b0,layer_2_1[3183:3176]} - {1'b0, layer_1_1[3183:3176]};
      mid_1[1] = {1'b0,layer_2_1[3191:3184]} - {1'b0, layer_1_1[3191:3184]};
      mid_1[2] = {1'b0,layer_2_1[3199:3192]} - {1'b0, layer_1_1[3199:3192]};
      mid_2[0] = {1'b0,layer_2_2[3183:3176]} - {1'b0, layer_1_2[3183:3176]};
      mid_2[1] = {1'b0,layer_2_2[3191:3184]} - {1'b0, layer_1_2[3191:3184]};
      mid_2[2] = {1'b0,layer_2_2[3199:3192]} - {1'b0, layer_1_2[3199:3192]};
      btm_0[0] = {1'b0,layer_3_0[3183:3176]} - {1'b0, layer_2_0[3183:3176]};
      btm_0[1] = {1'b0,layer_3_0[3191:3184]} - {1'b0, layer_2_0[3191:3184]};
      btm_0[2] = {1'b0,layer_3_0[3199:3192]} - {1'b0, layer_2_0[3199:3192]};
      btm_1[0] = {1'b0,layer_3_1[3183:3176]} - {1'b0, layer_2_1[3183:3176]};
      btm_1[1] = {1'b0,layer_3_1[3191:3184]} - {1'b0, layer_2_1[3191:3184]};
      btm_1[2] = {1'b0,layer_3_1[3199:3192]} - {1'b0, layer_2_1[3199:3192]};
      btm_2[0] = {1'b0,layer_3_2[3183:3176]} - {1'b0, layer_2_2[3183:3176]};
      btm_2[1] = {1'b0,layer_3_2[3191:3184]} - {1'b0, layer_2_2[3191:3184]};
      btm_2[2] = {1'b0,layer_3_2[3199:3192]} - {1'b0, layer_2_2[3199:3192]};
    end
    'd399: begin
      top_0[0] = {1'b0,layer_1_0[3191:3184]} - {1'b0, layer_0_0[3191:3184]};
      top_0[1] = {1'b0,layer_1_0[3199:3192]} - {1'b0, layer_0_0[3199:3192]};
      top_0[2] = {1'b0,layer_1_0[3207:3200]} - {1'b0, layer_0_0[3207:3200]};
      top_1[0] = {1'b0,layer_1_1[3191:3184]} - {1'b0, layer_0_1[3191:3184]};
      top_1[1] = {1'b0,layer_1_1[3199:3192]} - {1'b0, layer_0_1[3199:3192]};
      top_1[2] = {1'b0,layer_1_1[3207:3200]} - {1'b0, layer_0_1[3207:3200]};
      top_2[0] = {1'b0,layer_1_2[3191:3184]} - {1'b0, layer_0_2[3191:3184]};
      top_2[1] = {1'b0,layer_1_2[3199:3192]} - {1'b0, layer_0_2[3199:3192]};
      top_2[2] = {1'b0,layer_1_2[3207:3200]} - {1'b0, layer_0_2[3207:3200]};
      mid_0[0] = {1'b0,layer_2_0[3191:3184]} - {1'b0, layer_1_0[3191:3184]};
      mid_0[1] = {1'b0,layer_2_0[3199:3192]} - {1'b0, layer_1_0[3199:3192]};
      mid_0[2] = {1'b0,layer_2_0[3207:3200]} - {1'b0, layer_1_0[3207:3200]};
      mid_1[0] = {1'b0,layer_2_1[3191:3184]} - {1'b0, layer_1_1[3191:3184]};
      mid_1[1] = {1'b0,layer_2_1[3199:3192]} - {1'b0, layer_1_1[3199:3192]};
      mid_1[2] = {1'b0,layer_2_1[3207:3200]} - {1'b0, layer_1_1[3207:3200]};
      mid_2[0] = {1'b0,layer_2_2[3191:3184]} - {1'b0, layer_1_2[3191:3184]};
      mid_2[1] = {1'b0,layer_2_2[3199:3192]} - {1'b0, layer_1_2[3199:3192]};
      mid_2[2] = {1'b0,layer_2_2[3207:3200]} - {1'b0, layer_1_2[3207:3200]};
      btm_0[0] = {1'b0,layer_3_0[3191:3184]} - {1'b0, layer_2_0[3191:3184]};
      btm_0[1] = {1'b0,layer_3_0[3199:3192]} - {1'b0, layer_2_0[3199:3192]};
      btm_0[2] = {1'b0,layer_3_0[3207:3200]} - {1'b0, layer_2_0[3207:3200]};
      btm_1[0] = {1'b0,layer_3_1[3191:3184]} - {1'b0, layer_2_1[3191:3184]};
      btm_1[1] = {1'b0,layer_3_1[3199:3192]} - {1'b0, layer_2_1[3199:3192]};
      btm_1[2] = {1'b0,layer_3_1[3207:3200]} - {1'b0, layer_2_1[3207:3200]};
      btm_2[0] = {1'b0,layer_3_2[3191:3184]} - {1'b0, layer_2_2[3191:3184]};
      btm_2[1] = {1'b0,layer_3_2[3199:3192]} - {1'b0, layer_2_2[3199:3192]};
      btm_2[2] = {1'b0,layer_3_2[3207:3200]} - {1'b0, layer_2_2[3207:3200]};
    end
    'd400: begin
      top_0[0] = {1'b0,layer_1_0[3199:3192]} - {1'b0, layer_0_0[3199:3192]};
      top_0[1] = {1'b0,layer_1_0[3207:3200]} - {1'b0, layer_0_0[3207:3200]};
      top_0[2] = {1'b0,layer_1_0[3215:3208]} - {1'b0, layer_0_0[3215:3208]};
      top_1[0] = {1'b0,layer_1_1[3199:3192]} - {1'b0, layer_0_1[3199:3192]};
      top_1[1] = {1'b0,layer_1_1[3207:3200]} - {1'b0, layer_0_1[3207:3200]};
      top_1[2] = {1'b0,layer_1_1[3215:3208]} - {1'b0, layer_0_1[3215:3208]};
      top_2[0] = {1'b0,layer_1_2[3199:3192]} - {1'b0, layer_0_2[3199:3192]};
      top_2[1] = {1'b0,layer_1_2[3207:3200]} - {1'b0, layer_0_2[3207:3200]};
      top_2[2] = {1'b0,layer_1_2[3215:3208]} - {1'b0, layer_0_2[3215:3208]};
      mid_0[0] = {1'b0,layer_2_0[3199:3192]} - {1'b0, layer_1_0[3199:3192]};
      mid_0[1] = {1'b0,layer_2_0[3207:3200]} - {1'b0, layer_1_0[3207:3200]};
      mid_0[2] = {1'b0,layer_2_0[3215:3208]} - {1'b0, layer_1_0[3215:3208]};
      mid_1[0] = {1'b0,layer_2_1[3199:3192]} - {1'b0, layer_1_1[3199:3192]};
      mid_1[1] = {1'b0,layer_2_1[3207:3200]} - {1'b0, layer_1_1[3207:3200]};
      mid_1[2] = {1'b0,layer_2_1[3215:3208]} - {1'b0, layer_1_1[3215:3208]};
      mid_2[0] = {1'b0,layer_2_2[3199:3192]} - {1'b0, layer_1_2[3199:3192]};
      mid_2[1] = {1'b0,layer_2_2[3207:3200]} - {1'b0, layer_1_2[3207:3200]};
      mid_2[2] = {1'b0,layer_2_2[3215:3208]} - {1'b0, layer_1_2[3215:3208]};
      btm_0[0] = {1'b0,layer_3_0[3199:3192]} - {1'b0, layer_2_0[3199:3192]};
      btm_0[1] = {1'b0,layer_3_0[3207:3200]} - {1'b0, layer_2_0[3207:3200]};
      btm_0[2] = {1'b0,layer_3_0[3215:3208]} - {1'b0, layer_2_0[3215:3208]};
      btm_1[0] = {1'b0,layer_3_1[3199:3192]} - {1'b0, layer_2_1[3199:3192]};
      btm_1[1] = {1'b0,layer_3_1[3207:3200]} - {1'b0, layer_2_1[3207:3200]};
      btm_1[2] = {1'b0,layer_3_1[3215:3208]} - {1'b0, layer_2_1[3215:3208]};
      btm_2[0] = {1'b0,layer_3_2[3199:3192]} - {1'b0, layer_2_2[3199:3192]};
      btm_2[1] = {1'b0,layer_3_2[3207:3200]} - {1'b0, layer_2_2[3207:3200]};
      btm_2[2] = {1'b0,layer_3_2[3215:3208]} - {1'b0, layer_2_2[3215:3208]};
    end
    'd401: begin
      top_0[0] = {1'b0,layer_1_0[3207:3200]} - {1'b0, layer_0_0[3207:3200]};
      top_0[1] = {1'b0,layer_1_0[3215:3208]} - {1'b0, layer_0_0[3215:3208]};
      top_0[2] = {1'b0,layer_1_0[3223:3216]} - {1'b0, layer_0_0[3223:3216]};
      top_1[0] = {1'b0,layer_1_1[3207:3200]} - {1'b0, layer_0_1[3207:3200]};
      top_1[1] = {1'b0,layer_1_1[3215:3208]} - {1'b0, layer_0_1[3215:3208]};
      top_1[2] = {1'b0,layer_1_1[3223:3216]} - {1'b0, layer_0_1[3223:3216]};
      top_2[0] = {1'b0,layer_1_2[3207:3200]} - {1'b0, layer_0_2[3207:3200]};
      top_2[1] = {1'b0,layer_1_2[3215:3208]} - {1'b0, layer_0_2[3215:3208]};
      top_2[2] = {1'b0,layer_1_2[3223:3216]} - {1'b0, layer_0_2[3223:3216]};
      mid_0[0] = {1'b0,layer_2_0[3207:3200]} - {1'b0, layer_1_0[3207:3200]};
      mid_0[1] = {1'b0,layer_2_0[3215:3208]} - {1'b0, layer_1_0[3215:3208]};
      mid_0[2] = {1'b0,layer_2_0[3223:3216]} - {1'b0, layer_1_0[3223:3216]};
      mid_1[0] = {1'b0,layer_2_1[3207:3200]} - {1'b0, layer_1_1[3207:3200]};
      mid_1[1] = {1'b0,layer_2_1[3215:3208]} - {1'b0, layer_1_1[3215:3208]};
      mid_1[2] = {1'b0,layer_2_1[3223:3216]} - {1'b0, layer_1_1[3223:3216]};
      mid_2[0] = {1'b0,layer_2_2[3207:3200]} - {1'b0, layer_1_2[3207:3200]};
      mid_2[1] = {1'b0,layer_2_2[3215:3208]} - {1'b0, layer_1_2[3215:3208]};
      mid_2[2] = {1'b0,layer_2_2[3223:3216]} - {1'b0, layer_1_2[3223:3216]};
      btm_0[0] = {1'b0,layer_3_0[3207:3200]} - {1'b0, layer_2_0[3207:3200]};
      btm_0[1] = {1'b0,layer_3_0[3215:3208]} - {1'b0, layer_2_0[3215:3208]};
      btm_0[2] = {1'b0,layer_3_0[3223:3216]} - {1'b0, layer_2_0[3223:3216]};
      btm_1[0] = {1'b0,layer_3_1[3207:3200]} - {1'b0, layer_2_1[3207:3200]};
      btm_1[1] = {1'b0,layer_3_1[3215:3208]} - {1'b0, layer_2_1[3215:3208]};
      btm_1[2] = {1'b0,layer_3_1[3223:3216]} - {1'b0, layer_2_1[3223:3216]};
      btm_2[0] = {1'b0,layer_3_2[3207:3200]} - {1'b0, layer_2_2[3207:3200]};
      btm_2[1] = {1'b0,layer_3_2[3215:3208]} - {1'b0, layer_2_2[3215:3208]};
      btm_2[2] = {1'b0,layer_3_2[3223:3216]} - {1'b0, layer_2_2[3223:3216]};
    end
    'd402: begin
      top_0[0] = {1'b0,layer_1_0[3215:3208]} - {1'b0, layer_0_0[3215:3208]};
      top_0[1] = {1'b0,layer_1_0[3223:3216]} - {1'b0, layer_0_0[3223:3216]};
      top_0[2] = {1'b0,layer_1_0[3231:3224]} - {1'b0, layer_0_0[3231:3224]};
      top_1[0] = {1'b0,layer_1_1[3215:3208]} - {1'b0, layer_0_1[3215:3208]};
      top_1[1] = {1'b0,layer_1_1[3223:3216]} - {1'b0, layer_0_1[3223:3216]};
      top_1[2] = {1'b0,layer_1_1[3231:3224]} - {1'b0, layer_0_1[3231:3224]};
      top_2[0] = {1'b0,layer_1_2[3215:3208]} - {1'b0, layer_0_2[3215:3208]};
      top_2[1] = {1'b0,layer_1_2[3223:3216]} - {1'b0, layer_0_2[3223:3216]};
      top_2[2] = {1'b0,layer_1_2[3231:3224]} - {1'b0, layer_0_2[3231:3224]};
      mid_0[0] = {1'b0,layer_2_0[3215:3208]} - {1'b0, layer_1_0[3215:3208]};
      mid_0[1] = {1'b0,layer_2_0[3223:3216]} - {1'b0, layer_1_0[3223:3216]};
      mid_0[2] = {1'b0,layer_2_0[3231:3224]} - {1'b0, layer_1_0[3231:3224]};
      mid_1[0] = {1'b0,layer_2_1[3215:3208]} - {1'b0, layer_1_1[3215:3208]};
      mid_1[1] = {1'b0,layer_2_1[3223:3216]} - {1'b0, layer_1_1[3223:3216]};
      mid_1[2] = {1'b0,layer_2_1[3231:3224]} - {1'b0, layer_1_1[3231:3224]};
      mid_2[0] = {1'b0,layer_2_2[3215:3208]} - {1'b0, layer_1_2[3215:3208]};
      mid_2[1] = {1'b0,layer_2_2[3223:3216]} - {1'b0, layer_1_2[3223:3216]};
      mid_2[2] = {1'b0,layer_2_2[3231:3224]} - {1'b0, layer_1_2[3231:3224]};
      btm_0[0] = {1'b0,layer_3_0[3215:3208]} - {1'b0, layer_2_0[3215:3208]};
      btm_0[1] = {1'b0,layer_3_0[3223:3216]} - {1'b0, layer_2_0[3223:3216]};
      btm_0[2] = {1'b0,layer_3_0[3231:3224]} - {1'b0, layer_2_0[3231:3224]};
      btm_1[0] = {1'b0,layer_3_1[3215:3208]} - {1'b0, layer_2_1[3215:3208]};
      btm_1[1] = {1'b0,layer_3_1[3223:3216]} - {1'b0, layer_2_1[3223:3216]};
      btm_1[2] = {1'b0,layer_3_1[3231:3224]} - {1'b0, layer_2_1[3231:3224]};
      btm_2[0] = {1'b0,layer_3_2[3215:3208]} - {1'b0, layer_2_2[3215:3208]};
      btm_2[1] = {1'b0,layer_3_2[3223:3216]} - {1'b0, layer_2_2[3223:3216]};
      btm_2[2] = {1'b0,layer_3_2[3231:3224]} - {1'b0, layer_2_2[3231:3224]};
    end
    'd403: begin
      top_0[0] = {1'b0,layer_1_0[3223:3216]} - {1'b0, layer_0_0[3223:3216]};
      top_0[1] = {1'b0,layer_1_0[3231:3224]} - {1'b0, layer_0_0[3231:3224]};
      top_0[2] = {1'b0,layer_1_0[3239:3232]} - {1'b0, layer_0_0[3239:3232]};
      top_1[0] = {1'b0,layer_1_1[3223:3216]} - {1'b0, layer_0_1[3223:3216]};
      top_1[1] = {1'b0,layer_1_1[3231:3224]} - {1'b0, layer_0_1[3231:3224]};
      top_1[2] = {1'b0,layer_1_1[3239:3232]} - {1'b0, layer_0_1[3239:3232]};
      top_2[0] = {1'b0,layer_1_2[3223:3216]} - {1'b0, layer_0_2[3223:3216]};
      top_2[1] = {1'b0,layer_1_2[3231:3224]} - {1'b0, layer_0_2[3231:3224]};
      top_2[2] = {1'b0,layer_1_2[3239:3232]} - {1'b0, layer_0_2[3239:3232]};
      mid_0[0] = {1'b0,layer_2_0[3223:3216]} - {1'b0, layer_1_0[3223:3216]};
      mid_0[1] = {1'b0,layer_2_0[3231:3224]} - {1'b0, layer_1_0[3231:3224]};
      mid_0[2] = {1'b0,layer_2_0[3239:3232]} - {1'b0, layer_1_0[3239:3232]};
      mid_1[0] = {1'b0,layer_2_1[3223:3216]} - {1'b0, layer_1_1[3223:3216]};
      mid_1[1] = {1'b0,layer_2_1[3231:3224]} - {1'b0, layer_1_1[3231:3224]};
      mid_1[2] = {1'b0,layer_2_1[3239:3232]} - {1'b0, layer_1_1[3239:3232]};
      mid_2[0] = {1'b0,layer_2_2[3223:3216]} - {1'b0, layer_1_2[3223:3216]};
      mid_2[1] = {1'b0,layer_2_2[3231:3224]} - {1'b0, layer_1_2[3231:3224]};
      mid_2[2] = {1'b0,layer_2_2[3239:3232]} - {1'b0, layer_1_2[3239:3232]};
      btm_0[0] = {1'b0,layer_3_0[3223:3216]} - {1'b0, layer_2_0[3223:3216]};
      btm_0[1] = {1'b0,layer_3_0[3231:3224]} - {1'b0, layer_2_0[3231:3224]};
      btm_0[2] = {1'b0,layer_3_0[3239:3232]} - {1'b0, layer_2_0[3239:3232]};
      btm_1[0] = {1'b0,layer_3_1[3223:3216]} - {1'b0, layer_2_1[3223:3216]};
      btm_1[1] = {1'b0,layer_3_1[3231:3224]} - {1'b0, layer_2_1[3231:3224]};
      btm_1[2] = {1'b0,layer_3_1[3239:3232]} - {1'b0, layer_2_1[3239:3232]};
      btm_2[0] = {1'b0,layer_3_2[3223:3216]} - {1'b0, layer_2_2[3223:3216]};
      btm_2[1] = {1'b0,layer_3_2[3231:3224]} - {1'b0, layer_2_2[3231:3224]};
      btm_2[2] = {1'b0,layer_3_2[3239:3232]} - {1'b0, layer_2_2[3239:3232]};
    end
    'd404: begin
      top_0[0] = {1'b0,layer_1_0[3231:3224]} - {1'b0, layer_0_0[3231:3224]};
      top_0[1] = {1'b0,layer_1_0[3239:3232]} - {1'b0, layer_0_0[3239:3232]};
      top_0[2] = {1'b0,layer_1_0[3247:3240]} - {1'b0, layer_0_0[3247:3240]};
      top_1[0] = {1'b0,layer_1_1[3231:3224]} - {1'b0, layer_0_1[3231:3224]};
      top_1[1] = {1'b0,layer_1_1[3239:3232]} - {1'b0, layer_0_1[3239:3232]};
      top_1[2] = {1'b0,layer_1_1[3247:3240]} - {1'b0, layer_0_1[3247:3240]};
      top_2[0] = {1'b0,layer_1_2[3231:3224]} - {1'b0, layer_0_2[3231:3224]};
      top_2[1] = {1'b0,layer_1_2[3239:3232]} - {1'b0, layer_0_2[3239:3232]};
      top_2[2] = {1'b0,layer_1_2[3247:3240]} - {1'b0, layer_0_2[3247:3240]};
      mid_0[0] = {1'b0,layer_2_0[3231:3224]} - {1'b0, layer_1_0[3231:3224]};
      mid_0[1] = {1'b0,layer_2_0[3239:3232]} - {1'b0, layer_1_0[3239:3232]};
      mid_0[2] = {1'b0,layer_2_0[3247:3240]} - {1'b0, layer_1_0[3247:3240]};
      mid_1[0] = {1'b0,layer_2_1[3231:3224]} - {1'b0, layer_1_1[3231:3224]};
      mid_1[1] = {1'b0,layer_2_1[3239:3232]} - {1'b0, layer_1_1[3239:3232]};
      mid_1[2] = {1'b0,layer_2_1[3247:3240]} - {1'b0, layer_1_1[3247:3240]};
      mid_2[0] = {1'b0,layer_2_2[3231:3224]} - {1'b0, layer_1_2[3231:3224]};
      mid_2[1] = {1'b0,layer_2_2[3239:3232]} - {1'b0, layer_1_2[3239:3232]};
      mid_2[2] = {1'b0,layer_2_2[3247:3240]} - {1'b0, layer_1_2[3247:3240]};
      btm_0[0] = {1'b0,layer_3_0[3231:3224]} - {1'b0, layer_2_0[3231:3224]};
      btm_0[1] = {1'b0,layer_3_0[3239:3232]} - {1'b0, layer_2_0[3239:3232]};
      btm_0[2] = {1'b0,layer_3_0[3247:3240]} - {1'b0, layer_2_0[3247:3240]};
      btm_1[0] = {1'b0,layer_3_1[3231:3224]} - {1'b0, layer_2_1[3231:3224]};
      btm_1[1] = {1'b0,layer_3_1[3239:3232]} - {1'b0, layer_2_1[3239:3232]};
      btm_1[2] = {1'b0,layer_3_1[3247:3240]} - {1'b0, layer_2_1[3247:3240]};
      btm_2[0] = {1'b0,layer_3_2[3231:3224]} - {1'b0, layer_2_2[3231:3224]};
      btm_2[1] = {1'b0,layer_3_2[3239:3232]} - {1'b0, layer_2_2[3239:3232]};
      btm_2[2] = {1'b0,layer_3_2[3247:3240]} - {1'b0, layer_2_2[3247:3240]};
    end
    'd405: begin
      top_0[0] = {1'b0,layer_1_0[3239:3232]} - {1'b0, layer_0_0[3239:3232]};
      top_0[1] = {1'b0,layer_1_0[3247:3240]} - {1'b0, layer_0_0[3247:3240]};
      top_0[2] = {1'b0,layer_1_0[3255:3248]} - {1'b0, layer_0_0[3255:3248]};
      top_1[0] = {1'b0,layer_1_1[3239:3232]} - {1'b0, layer_0_1[3239:3232]};
      top_1[1] = {1'b0,layer_1_1[3247:3240]} - {1'b0, layer_0_1[3247:3240]};
      top_1[2] = {1'b0,layer_1_1[3255:3248]} - {1'b0, layer_0_1[3255:3248]};
      top_2[0] = {1'b0,layer_1_2[3239:3232]} - {1'b0, layer_0_2[3239:3232]};
      top_2[1] = {1'b0,layer_1_2[3247:3240]} - {1'b0, layer_0_2[3247:3240]};
      top_2[2] = {1'b0,layer_1_2[3255:3248]} - {1'b0, layer_0_2[3255:3248]};
      mid_0[0] = {1'b0,layer_2_0[3239:3232]} - {1'b0, layer_1_0[3239:3232]};
      mid_0[1] = {1'b0,layer_2_0[3247:3240]} - {1'b0, layer_1_0[3247:3240]};
      mid_0[2] = {1'b0,layer_2_0[3255:3248]} - {1'b0, layer_1_0[3255:3248]};
      mid_1[0] = {1'b0,layer_2_1[3239:3232]} - {1'b0, layer_1_1[3239:3232]};
      mid_1[1] = {1'b0,layer_2_1[3247:3240]} - {1'b0, layer_1_1[3247:3240]};
      mid_1[2] = {1'b0,layer_2_1[3255:3248]} - {1'b0, layer_1_1[3255:3248]};
      mid_2[0] = {1'b0,layer_2_2[3239:3232]} - {1'b0, layer_1_2[3239:3232]};
      mid_2[1] = {1'b0,layer_2_2[3247:3240]} - {1'b0, layer_1_2[3247:3240]};
      mid_2[2] = {1'b0,layer_2_2[3255:3248]} - {1'b0, layer_1_2[3255:3248]};
      btm_0[0] = {1'b0,layer_3_0[3239:3232]} - {1'b0, layer_2_0[3239:3232]};
      btm_0[1] = {1'b0,layer_3_0[3247:3240]} - {1'b0, layer_2_0[3247:3240]};
      btm_0[2] = {1'b0,layer_3_0[3255:3248]} - {1'b0, layer_2_0[3255:3248]};
      btm_1[0] = {1'b0,layer_3_1[3239:3232]} - {1'b0, layer_2_1[3239:3232]};
      btm_1[1] = {1'b0,layer_3_1[3247:3240]} - {1'b0, layer_2_1[3247:3240]};
      btm_1[2] = {1'b0,layer_3_1[3255:3248]} - {1'b0, layer_2_1[3255:3248]};
      btm_2[0] = {1'b0,layer_3_2[3239:3232]} - {1'b0, layer_2_2[3239:3232]};
      btm_2[1] = {1'b0,layer_3_2[3247:3240]} - {1'b0, layer_2_2[3247:3240]};
      btm_2[2] = {1'b0,layer_3_2[3255:3248]} - {1'b0, layer_2_2[3255:3248]};
    end
    'd406: begin
      top_0[0] = {1'b0,layer_1_0[3247:3240]} - {1'b0, layer_0_0[3247:3240]};
      top_0[1] = {1'b0,layer_1_0[3255:3248]} - {1'b0, layer_0_0[3255:3248]};
      top_0[2] = {1'b0,layer_1_0[3263:3256]} - {1'b0, layer_0_0[3263:3256]};
      top_1[0] = {1'b0,layer_1_1[3247:3240]} - {1'b0, layer_0_1[3247:3240]};
      top_1[1] = {1'b0,layer_1_1[3255:3248]} - {1'b0, layer_0_1[3255:3248]};
      top_1[2] = {1'b0,layer_1_1[3263:3256]} - {1'b0, layer_0_1[3263:3256]};
      top_2[0] = {1'b0,layer_1_2[3247:3240]} - {1'b0, layer_0_2[3247:3240]};
      top_2[1] = {1'b0,layer_1_2[3255:3248]} - {1'b0, layer_0_2[3255:3248]};
      top_2[2] = {1'b0,layer_1_2[3263:3256]} - {1'b0, layer_0_2[3263:3256]};
      mid_0[0] = {1'b0,layer_2_0[3247:3240]} - {1'b0, layer_1_0[3247:3240]};
      mid_0[1] = {1'b0,layer_2_0[3255:3248]} - {1'b0, layer_1_0[3255:3248]};
      mid_0[2] = {1'b0,layer_2_0[3263:3256]} - {1'b0, layer_1_0[3263:3256]};
      mid_1[0] = {1'b0,layer_2_1[3247:3240]} - {1'b0, layer_1_1[3247:3240]};
      mid_1[1] = {1'b0,layer_2_1[3255:3248]} - {1'b0, layer_1_1[3255:3248]};
      mid_1[2] = {1'b0,layer_2_1[3263:3256]} - {1'b0, layer_1_1[3263:3256]};
      mid_2[0] = {1'b0,layer_2_2[3247:3240]} - {1'b0, layer_1_2[3247:3240]};
      mid_2[1] = {1'b0,layer_2_2[3255:3248]} - {1'b0, layer_1_2[3255:3248]};
      mid_2[2] = {1'b0,layer_2_2[3263:3256]} - {1'b0, layer_1_2[3263:3256]};
      btm_0[0] = {1'b0,layer_3_0[3247:3240]} - {1'b0, layer_2_0[3247:3240]};
      btm_0[1] = {1'b0,layer_3_0[3255:3248]} - {1'b0, layer_2_0[3255:3248]};
      btm_0[2] = {1'b0,layer_3_0[3263:3256]} - {1'b0, layer_2_0[3263:3256]};
      btm_1[0] = {1'b0,layer_3_1[3247:3240]} - {1'b0, layer_2_1[3247:3240]};
      btm_1[1] = {1'b0,layer_3_1[3255:3248]} - {1'b0, layer_2_1[3255:3248]};
      btm_1[2] = {1'b0,layer_3_1[3263:3256]} - {1'b0, layer_2_1[3263:3256]};
      btm_2[0] = {1'b0,layer_3_2[3247:3240]} - {1'b0, layer_2_2[3247:3240]};
      btm_2[1] = {1'b0,layer_3_2[3255:3248]} - {1'b0, layer_2_2[3255:3248]};
      btm_2[2] = {1'b0,layer_3_2[3263:3256]} - {1'b0, layer_2_2[3263:3256]};
    end
    'd407: begin
      top_0[0] = {1'b0,layer_1_0[3255:3248]} - {1'b0, layer_0_0[3255:3248]};
      top_0[1] = {1'b0,layer_1_0[3263:3256]} - {1'b0, layer_0_0[3263:3256]};
      top_0[2] = {1'b0,layer_1_0[3271:3264]} - {1'b0, layer_0_0[3271:3264]};
      top_1[0] = {1'b0,layer_1_1[3255:3248]} - {1'b0, layer_0_1[3255:3248]};
      top_1[1] = {1'b0,layer_1_1[3263:3256]} - {1'b0, layer_0_1[3263:3256]};
      top_1[2] = {1'b0,layer_1_1[3271:3264]} - {1'b0, layer_0_1[3271:3264]};
      top_2[0] = {1'b0,layer_1_2[3255:3248]} - {1'b0, layer_0_2[3255:3248]};
      top_2[1] = {1'b0,layer_1_2[3263:3256]} - {1'b0, layer_0_2[3263:3256]};
      top_2[2] = {1'b0,layer_1_2[3271:3264]} - {1'b0, layer_0_2[3271:3264]};
      mid_0[0] = {1'b0,layer_2_0[3255:3248]} - {1'b0, layer_1_0[3255:3248]};
      mid_0[1] = {1'b0,layer_2_0[3263:3256]} - {1'b0, layer_1_0[3263:3256]};
      mid_0[2] = {1'b0,layer_2_0[3271:3264]} - {1'b0, layer_1_0[3271:3264]};
      mid_1[0] = {1'b0,layer_2_1[3255:3248]} - {1'b0, layer_1_1[3255:3248]};
      mid_1[1] = {1'b0,layer_2_1[3263:3256]} - {1'b0, layer_1_1[3263:3256]};
      mid_1[2] = {1'b0,layer_2_1[3271:3264]} - {1'b0, layer_1_1[3271:3264]};
      mid_2[0] = {1'b0,layer_2_2[3255:3248]} - {1'b0, layer_1_2[3255:3248]};
      mid_2[1] = {1'b0,layer_2_2[3263:3256]} - {1'b0, layer_1_2[3263:3256]};
      mid_2[2] = {1'b0,layer_2_2[3271:3264]} - {1'b0, layer_1_2[3271:3264]};
      btm_0[0] = {1'b0,layer_3_0[3255:3248]} - {1'b0, layer_2_0[3255:3248]};
      btm_0[1] = {1'b0,layer_3_0[3263:3256]} - {1'b0, layer_2_0[3263:3256]};
      btm_0[2] = {1'b0,layer_3_0[3271:3264]} - {1'b0, layer_2_0[3271:3264]};
      btm_1[0] = {1'b0,layer_3_1[3255:3248]} - {1'b0, layer_2_1[3255:3248]};
      btm_1[1] = {1'b0,layer_3_1[3263:3256]} - {1'b0, layer_2_1[3263:3256]};
      btm_1[2] = {1'b0,layer_3_1[3271:3264]} - {1'b0, layer_2_1[3271:3264]};
      btm_2[0] = {1'b0,layer_3_2[3255:3248]} - {1'b0, layer_2_2[3255:3248]};
      btm_2[1] = {1'b0,layer_3_2[3263:3256]} - {1'b0, layer_2_2[3263:3256]};
      btm_2[2] = {1'b0,layer_3_2[3271:3264]} - {1'b0, layer_2_2[3271:3264]};
    end
    'd408: begin
      top_0[0] = {1'b0,layer_1_0[3263:3256]} - {1'b0, layer_0_0[3263:3256]};
      top_0[1] = {1'b0,layer_1_0[3271:3264]} - {1'b0, layer_0_0[3271:3264]};
      top_0[2] = {1'b0,layer_1_0[3279:3272]} - {1'b0, layer_0_0[3279:3272]};
      top_1[0] = {1'b0,layer_1_1[3263:3256]} - {1'b0, layer_0_1[3263:3256]};
      top_1[1] = {1'b0,layer_1_1[3271:3264]} - {1'b0, layer_0_1[3271:3264]};
      top_1[2] = {1'b0,layer_1_1[3279:3272]} - {1'b0, layer_0_1[3279:3272]};
      top_2[0] = {1'b0,layer_1_2[3263:3256]} - {1'b0, layer_0_2[3263:3256]};
      top_2[1] = {1'b0,layer_1_2[3271:3264]} - {1'b0, layer_0_2[3271:3264]};
      top_2[2] = {1'b0,layer_1_2[3279:3272]} - {1'b0, layer_0_2[3279:3272]};
      mid_0[0] = {1'b0,layer_2_0[3263:3256]} - {1'b0, layer_1_0[3263:3256]};
      mid_0[1] = {1'b0,layer_2_0[3271:3264]} - {1'b0, layer_1_0[3271:3264]};
      mid_0[2] = {1'b0,layer_2_0[3279:3272]} - {1'b0, layer_1_0[3279:3272]};
      mid_1[0] = {1'b0,layer_2_1[3263:3256]} - {1'b0, layer_1_1[3263:3256]};
      mid_1[1] = {1'b0,layer_2_1[3271:3264]} - {1'b0, layer_1_1[3271:3264]};
      mid_1[2] = {1'b0,layer_2_1[3279:3272]} - {1'b0, layer_1_1[3279:3272]};
      mid_2[0] = {1'b0,layer_2_2[3263:3256]} - {1'b0, layer_1_2[3263:3256]};
      mid_2[1] = {1'b0,layer_2_2[3271:3264]} - {1'b0, layer_1_2[3271:3264]};
      mid_2[2] = {1'b0,layer_2_2[3279:3272]} - {1'b0, layer_1_2[3279:3272]};
      btm_0[0] = {1'b0,layer_3_0[3263:3256]} - {1'b0, layer_2_0[3263:3256]};
      btm_0[1] = {1'b0,layer_3_0[3271:3264]} - {1'b0, layer_2_0[3271:3264]};
      btm_0[2] = {1'b0,layer_3_0[3279:3272]} - {1'b0, layer_2_0[3279:3272]};
      btm_1[0] = {1'b0,layer_3_1[3263:3256]} - {1'b0, layer_2_1[3263:3256]};
      btm_1[1] = {1'b0,layer_3_1[3271:3264]} - {1'b0, layer_2_1[3271:3264]};
      btm_1[2] = {1'b0,layer_3_1[3279:3272]} - {1'b0, layer_2_1[3279:3272]};
      btm_2[0] = {1'b0,layer_3_2[3263:3256]} - {1'b0, layer_2_2[3263:3256]};
      btm_2[1] = {1'b0,layer_3_2[3271:3264]} - {1'b0, layer_2_2[3271:3264]};
      btm_2[2] = {1'b0,layer_3_2[3279:3272]} - {1'b0, layer_2_2[3279:3272]};
    end
    'd409: begin
      top_0[0] = {1'b0,layer_1_0[3271:3264]} - {1'b0, layer_0_0[3271:3264]};
      top_0[1] = {1'b0,layer_1_0[3279:3272]} - {1'b0, layer_0_0[3279:3272]};
      top_0[2] = {1'b0,layer_1_0[3287:3280]} - {1'b0, layer_0_0[3287:3280]};
      top_1[0] = {1'b0,layer_1_1[3271:3264]} - {1'b0, layer_0_1[3271:3264]};
      top_1[1] = {1'b0,layer_1_1[3279:3272]} - {1'b0, layer_0_1[3279:3272]};
      top_1[2] = {1'b0,layer_1_1[3287:3280]} - {1'b0, layer_0_1[3287:3280]};
      top_2[0] = {1'b0,layer_1_2[3271:3264]} - {1'b0, layer_0_2[3271:3264]};
      top_2[1] = {1'b0,layer_1_2[3279:3272]} - {1'b0, layer_0_2[3279:3272]};
      top_2[2] = {1'b0,layer_1_2[3287:3280]} - {1'b0, layer_0_2[3287:3280]};
      mid_0[0] = {1'b0,layer_2_0[3271:3264]} - {1'b0, layer_1_0[3271:3264]};
      mid_0[1] = {1'b0,layer_2_0[3279:3272]} - {1'b0, layer_1_0[3279:3272]};
      mid_0[2] = {1'b0,layer_2_0[3287:3280]} - {1'b0, layer_1_0[3287:3280]};
      mid_1[0] = {1'b0,layer_2_1[3271:3264]} - {1'b0, layer_1_1[3271:3264]};
      mid_1[1] = {1'b0,layer_2_1[3279:3272]} - {1'b0, layer_1_1[3279:3272]};
      mid_1[2] = {1'b0,layer_2_1[3287:3280]} - {1'b0, layer_1_1[3287:3280]};
      mid_2[0] = {1'b0,layer_2_2[3271:3264]} - {1'b0, layer_1_2[3271:3264]};
      mid_2[1] = {1'b0,layer_2_2[3279:3272]} - {1'b0, layer_1_2[3279:3272]};
      mid_2[2] = {1'b0,layer_2_2[3287:3280]} - {1'b0, layer_1_2[3287:3280]};
      btm_0[0] = {1'b0,layer_3_0[3271:3264]} - {1'b0, layer_2_0[3271:3264]};
      btm_0[1] = {1'b0,layer_3_0[3279:3272]} - {1'b0, layer_2_0[3279:3272]};
      btm_0[2] = {1'b0,layer_3_0[3287:3280]} - {1'b0, layer_2_0[3287:3280]};
      btm_1[0] = {1'b0,layer_3_1[3271:3264]} - {1'b0, layer_2_1[3271:3264]};
      btm_1[1] = {1'b0,layer_3_1[3279:3272]} - {1'b0, layer_2_1[3279:3272]};
      btm_1[2] = {1'b0,layer_3_1[3287:3280]} - {1'b0, layer_2_1[3287:3280]};
      btm_2[0] = {1'b0,layer_3_2[3271:3264]} - {1'b0, layer_2_2[3271:3264]};
      btm_2[1] = {1'b0,layer_3_2[3279:3272]} - {1'b0, layer_2_2[3279:3272]};
      btm_2[2] = {1'b0,layer_3_2[3287:3280]} - {1'b0, layer_2_2[3287:3280]};
    end
    'd410: begin
      top_0[0] = {1'b0,layer_1_0[3279:3272]} - {1'b0, layer_0_0[3279:3272]};
      top_0[1] = {1'b0,layer_1_0[3287:3280]} - {1'b0, layer_0_0[3287:3280]};
      top_0[2] = {1'b0,layer_1_0[3295:3288]} - {1'b0, layer_0_0[3295:3288]};
      top_1[0] = {1'b0,layer_1_1[3279:3272]} - {1'b0, layer_0_1[3279:3272]};
      top_1[1] = {1'b0,layer_1_1[3287:3280]} - {1'b0, layer_0_1[3287:3280]};
      top_1[2] = {1'b0,layer_1_1[3295:3288]} - {1'b0, layer_0_1[3295:3288]};
      top_2[0] = {1'b0,layer_1_2[3279:3272]} - {1'b0, layer_0_2[3279:3272]};
      top_2[1] = {1'b0,layer_1_2[3287:3280]} - {1'b0, layer_0_2[3287:3280]};
      top_2[2] = {1'b0,layer_1_2[3295:3288]} - {1'b0, layer_0_2[3295:3288]};
      mid_0[0] = {1'b0,layer_2_0[3279:3272]} - {1'b0, layer_1_0[3279:3272]};
      mid_0[1] = {1'b0,layer_2_0[3287:3280]} - {1'b0, layer_1_0[3287:3280]};
      mid_0[2] = {1'b0,layer_2_0[3295:3288]} - {1'b0, layer_1_0[3295:3288]};
      mid_1[0] = {1'b0,layer_2_1[3279:3272]} - {1'b0, layer_1_1[3279:3272]};
      mid_1[1] = {1'b0,layer_2_1[3287:3280]} - {1'b0, layer_1_1[3287:3280]};
      mid_1[2] = {1'b0,layer_2_1[3295:3288]} - {1'b0, layer_1_1[3295:3288]};
      mid_2[0] = {1'b0,layer_2_2[3279:3272]} - {1'b0, layer_1_2[3279:3272]};
      mid_2[1] = {1'b0,layer_2_2[3287:3280]} - {1'b0, layer_1_2[3287:3280]};
      mid_2[2] = {1'b0,layer_2_2[3295:3288]} - {1'b0, layer_1_2[3295:3288]};
      btm_0[0] = {1'b0,layer_3_0[3279:3272]} - {1'b0, layer_2_0[3279:3272]};
      btm_0[1] = {1'b0,layer_3_0[3287:3280]} - {1'b0, layer_2_0[3287:3280]};
      btm_0[2] = {1'b0,layer_3_0[3295:3288]} - {1'b0, layer_2_0[3295:3288]};
      btm_1[0] = {1'b0,layer_3_1[3279:3272]} - {1'b0, layer_2_1[3279:3272]};
      btm_1[1] = {1'b0,layer_3_1[3287:3280]} - {1'b0, layer_2_1[3287:3280]};
      btm_1[2] = {1'b0,layer_3_1[3295:3288]} - {1'b0, layer_2_1[3295:3288]};
      btm_2[0] = {1'b0,layer_3_2[3279:3272]} - {1'b0, layer_2_2[3279:3272]};
      btm_2[1] = {1'b0,layer_3_2[3287:3280]} - {1'b0, layer_2_2[3287:3280]};
      btm_2[2] = {1'b0,layer_3_2[3295:3288]} - {1'b0, layer_2_2[3295:3288]};
    end
    'd411: begin
      top_0[0] = {1'b0,layer_1_0[3287:3280]} - {1'b0, layer_0_0[3287:3280]};
      top_0[1] = {1'b0,layer_1_0[3295:3288]} - {1'b0, layer_0_0[3295:3288]};
      top_0[2] = {1'b0,layer_1_0[3303:3296]} - {1'b0, layer_0_0[3303:3296]};
      top_1[0] = {1'b0,layer_1_1[3287:3280]} - {1'b0, layer_0_1[3287:3280]};
      top_1[1] = {1'b0,layer_1_1[3295:3288]} - {1'b0, layer_0_1[3295:3288]};
      top_1[2] = {1'b0,layer_1_1[3303:3296]} - {1'b0, layer_0_1[3303:3296]};
      top_2[0] = {1'b0,layer_1_2[3287:3280]} - {1'b0, layer_0_2[3287:3280]};
      top_2[1] = {1'b0,layer_1_2[3295:3288]} - {1'b0, layer_0_2[3295:3288]};
      top_2[2] = {1'b0,layer_1_2[3303:3296]} - {1'b0, layer_0_2[3303:3296]};
      mid_0[0] = {1'b0,layer_2_0[3287:3280]} - {1'b0, layer_1_0[3287:3280]};
      mid_0[1] = {1'b0,layer_2_0[3295:3288]} - {1'b0, layer_1_0[3295:3288]};
      mid_0[2] = {1'b0,layer_2_0[3303:3296]} - {1'b0, layer_1_0[3303:3296]};
      mid_1[0] = {1'b0,layer_2_1[3287:3280]} - {1'b0, layer_1_1[3287:3280]};
      mid_1[1] = {1'b0,layer_2_1[3295:3288]} - {1'b0, layer_1_1[3295:3288]};
      mid_1[2] = {1'b0,layer_2_1[3303:3296]} - {1'b0, layer_1_1[3303:3296]};
      mid_2[0] = {1'b0,layer_2_2[3287:3280]} - {1'b0, layer_1_2[3287:3280]};
      mid_2[1] = {1'b0,layer_2_2[3295:3288]} - {1'b0, layer_1_2[3295:3288]};
      mid_2[2] = {1'b0,layer_2_2[3303:3296]} - {1'b0, layer_1_2[3303:3296]};
      btm_0[0] = {1'b0,layer_3_0[3287:3280]} - {1'b0, layer_2_0[3287:3280]};
      btm_0[1] = {1'b0,layer_3_0[3295:3288]} - {1'b0, layer_2_0[3295:3288]};
      btm_0[2] = {1'b0,layer_3_0[3303:3296]} - {1'b0, layer_2_0[3303:3296]};
      btm_1[0] = {1'b0,layer_3_1[3287:3280]} - {1'b0, layer_2_1[3287:3280]};
      btm_1[1] = {1'b0,layer_3_1[3295:3288]} - {1'b0, layer_2_1[3295:3288]};
      btm_1[2] = {1'b0,layer_3_1[3303:3296]} - {1'b0, layer_2_1[3303:3296]};
      btm_2[0] = {1'b0,layer_3_2[3287:3280]} - {1'b0, layer_2_2[3287:3280]};
      btm_2[1] = {1'b0,layer_3_2[3295:3288]} - {1'b0, layer_2_2[3295:3288]};
      btm_2[2] = {1'b0,layer_3_2[3303:3296]} - {1'b0, layer_2_2[3303:3296]};
    end
    'd412: begin
      top_0[0] = {1'b0,layer_1_0[3295:3288]} - {1'b0, layer_0_0[3295:3288]};
      top_0[1] = {1'b0,layer_1_0[3303:3296]} - {1'b0, layer_0_0[3303:3296]};
      top_0[2] = {1'b0,layer_1_0[3311:3304]} - {1'b0, layer_0_0[3311:3304]};
      top_1[0] = {1'b0,layer_1_1[3295:3288]} - {1'b0, layer_0_1[3295:3288]};
      top_1[1] = {1'b0,layer_1_1[3303:3296]} - {1'b0, layer_0_1[3303:3296]};
      top_1[2] = {1'b0,layer_1_1[3311:3304]} - {1'b0, layer_0_1[3311:3304]};
      top_2[0] = {1'b0,layer_1_2[3295:3288]} - {1'b0, layer_0_2[3295:3288]};
      top_2[1] = {1'b0,layer_1_2[3303:3296]} - {1'b0, layer_0_2[3303:3296]};
      top_2[2] = {1'b0,layer_1_2[3311:3304]} - {1'b0, layer_0_2[3311:3304]};
      mid_0[0] = {1'b0,layer_2_0[3295:3288]} - {1'b0, layer_1_0[3295:3288]};
      mid_0[1] = {1'b0,layer_2_0[3303:3296]} - {1'b0, layer_1_0[3303:3296]};
      mid_0[2] = {1'b0,layer_2_0[3311:3304]} - {1'b0, layer_1_0[3311:3304]};
      mid_1[0] = {1'b0,layer_2_1[3295:3288]} - {1'b0, layer_1_1[3295:3288]};
      mid_1[1] = {1'b0,layer_2_1[3303:3296]} - {1'b0, layer_1_1[3303:3296]};
      mid_1[2] = {1'b0,layer_2_1[3311:3304]} - {1'b0, layer_1_1[3311:3304]};
      mid_2[0] = {1'b0,layer_2_2[3295:3288]} - {1'b0, layer_1_2[3295:3288]};
      mid_2[1] = {1'b0,layer_2_2[3303:3296]} - {1'b0, layer_1_2[3303:3296]};
      mid_2[2] = {1'b0,layer_2_2[3311:3304]} - {1'b0, layer_1_2[3311:3304]};
      btm_0[0] = {1'b0,layer_3_0[3295:3288]} - {1'b0, layer_2_0[3295:3288]};
      btm_0[1] = {1'b0,layer_3_0[3303:3296]} - {1'b0, layer_2_0[3303:3296]};
      btm_0[2] = {1'b0,layer_3_0[3311:3304]} - {1'b0, layer_2_0[3311:3304]};
      btm_1[0] = {1'b0,layer_3_1[3295:3288]} - {1'b0, layer_2_1[3295:3288]};
      btm_1[1] = {1'b0,layer_3_1[3303:3296]} - {1'b0, layer_2_1[3303:3296]};
      btm_1[2] = {1'b0,layer_3_1[3311:3304]} - {1'b0, layer_2_1[3311:3304]};
      btm_2[0] = {1'b0,layer_3_2[3295:3288]} - {1'b0, layer_2_2[3295:3288]};
      btm_2[1] = {1'b0,layer_3_2[3303:3296]} - {1'b0, layer_2_2[3303:3296]};
      btm_2[2] = {1'b0,layer_3_2[3311:3304]} - {1'b0, layer_2_2[3311:3304]};
    end
    'd413: begin
      top_0[0] = {1'b0,layer_1_0[3303:3296]} - {1'b0, layer_0_0[3303:3296]};
      top_0[1] = {1'b0,layer_1_0[3311:3304]} - {1'b0, layer_0_0[3311:3304]};
      top_0[2] = {1'b0,layer_1_0[3319:3312]} - {1'b0, layer_0_0[3319:3312]};
      top_1[0] = {1'b0,layer_1_1[3303:3296]} - {1'b0, layer_0_1[3303:3296]};
      top_1[1] = {1'b0,layer_1_1[3311:3304]} - {1'b0, layer_0_1[3311:3304]};
      top_1[2] = {1'b0,layer_1_1[3319:3312]} - {1'b0, layer_0_1[3319:3312]};
      top_2[0] = {1'b0,layer_1_2[3303:3296]} - {1'b0, layer_0_2[3303:3296]};
      top_2[1] = {1'b0,layer_1_2[3311:3304]} - {1'b0, layer_0_2[3311:3304]};
      top_2[2] = {1'b0,layer_1_2[3319:3312]} - {1'b0, layer_0_2[3319:3312]};
      mid_0[0] = {1'b0,layer_2_0[3303:3296]} - {1'b0, layer_1_0[3303:3296]};
      mid_0[1] = {1'b0,layer_2_0[3311:3304]} - {1'b0, layer_1_0[3311:3304]};
      mid_0[2] = {1'b0,layer_2_0[3319:3312]} - {1'b0, layer_1_0[3319:3312]};
      mid_1[0] = {1'b0,layer_2_1[3303:3296]} - {1'b0, layer_1_1[3303:3296]};
      mid_1[1] = {1'b0,layer_2_1[3311:3304]} - {1'b0, layer_1_1[3311:3304]};
      mid_1[2] = {1'b0,layer_2_1[3319:3312]} - {1'b0, layer_1_1[3319:3312]};
      mid_2[0] = {1'b0,layer_2_2[3303:3296]} - {1'b0, layer_1_2[3303:3296]};
      mid_2[1] = {1'b0,layer_2_2[3311:3304]} - {1'b0, layer_1_2[3311:3304]};
      mid_2[2] = {1'b0,layer_2_2[3319:3312]} - {1'b0, layer_1_2[3319:3312]};
      btm_0[0] = {1'b0,layer_3_0[3303:3296]} - {1'b0, layer_2_0[3303:3296]};
      btm_0[1] = {1'b0,layer_3_0[3311:3304]} - {1'b0, layer_2_0[3311:3304]};
      btm_0[2] = {1'b0,layer_3_0[3319:3312]} - {1'b0, layer_2_0[3319:3312]};
      btm_1[0] = {1'b0,layer_3_1[3303:3296]} - {1'b0, layer_2_1[3303:3296]};
      btm_1[1] = {1'b0,layer_3_1[3311:3304]} - {1'b0, layer_2_1[3311:3304]};
      btm_1[2] = {1'b0,layer_3_1[3319:3312]} - {1'b0, layer_2_1[3319:3312]};
      btm_2[0] = {1'b0,layer_3_2[3303:3296]} - {1'b0, layer_2_2[3303:3296]};
      btm_2[1] = {1'b0,layer_3_2[3311:3304]} - {1'b0, layer_2_2[3311:3304]};
      btm_2[2] = {1'b0,layer_3_2[3319:3312]} - {1'b0, layer_2_2[3319:3312]};
    end
    'd414: begin
      top_0[0] = {1'b0,layer_1_0[3311:3304]} - {1'b0, layer_0_0[3311:3304]};
      top_0[1] = {1'b0,layer_1_0[3319:3312]} - {1'b0, layer_0_0[3319:3312]};
      top_0[2] = {1'b0,layer_1_0[3327:3320]} - {1'b0, layer_0_0[3327:3320]};
      top_1[0] = {1'b0,layer_1_1[3311:3304]} - {1'b0, layer_0_1[3311:3304]};
      top_1[1] = {1'b0,layer_1_1[3319:3312]} - {1'b0, layer_0_1[3319:3312]};
      top_1[2] = {1'b0,layer_1_1[3327:3320]} - {1'b0, layer_0_1[3327:3320]};
      top_2[0] = {1'b0,layer_1_2[3311:3304]} - {1'b0, layer_0_2[3311:3304]};
      top_2[1] = {1'b0,layer_1_2[3319:3312]} - {1'b0, layer_0_2[3319:3312]};
      top_2[2] = {1'b0,layer_1_2[3327:3320]} - {1'b0, layer_0_2[3327:3320]};
      mid_0[0] = {1'b0,layer_2_0[3311:3304]} - {1'b0, layer_1_0[3311:3304]};
      mid_0[1] = {1'b0,layer_2_0[3319:3312]} - {1'b0, layer_1_0[3319:3312]};
      mid_0[2] = {1'b0,layer_2_0[3327:3320]} - {1'b0, layer_1_0[3327:3320]};
      mid_1[0] = {1'b0,layer_2_1[3311:3304]} - {1'b0, layer_1_1[3311:3304]};
      mid_1[1] = {1'b0,layer_2_1[3319:3312]} - {1'b0, layer_1_1[3319:3312]};
      mid_1[2] = {1'b0,layer_2_1[3327:3320]} - {1'b0, layer_1_1[3327:3320]};
      mid_2[0] = {1'b0,layer_2_2[3311:3304]} - {1'b0, layer_1_2[3311:3304]};
      mid_2[1] = {1'b0,layer_2_2[3319:3312]} - {1'b0, layer_1_2[3319:3312]};
      mid_2[2] = {1'b0,layer_2_2[3327:3320]} - {1'b0, layer_1_2[3327:3320]};
      btm_0[0] = {1'b0,layer_3_0[3311:3304]} - {1'b0, layer_2_0[3311:3304]};
      btm_0[1] = {1'b0,layer_3_0[3319:3312]} - {1'b0, layer_2_0[3319:3312]};
      btm_0[2] = {1'b0,layer_3_0[3327:3320]} - {1'b0, layer_2_0[3327:3320]};
      btm_1[0] = {1'b0,layer_3_1[3311:3304]} - {1'b0, layer_2_1[3311:3304]};
      btm_1[1] = {1'b0,layer_3_1[3319:3312]} - {1'b0, layer_2_1[3319:3312]};
      btm_1[2] = {1'b0,layer_3_1[3327:3320]} - {1'b0, layer_2_1[3327:3320]};
      btm_2[0] = {1'b0,layer_3_2[3311:3304]} - {1'b0, layer_2_2[3311:3304]};
      btm_2[1] = {1'b0,layer_3_2[3319:3312]} - {1'b0, layer_2_2[3319:3312]};
      btm_2[2] = {1'b0,layer_3_2[3327:3320]} - {1'b0, layer_2_2[3327:3320]};
    end
    'd415: begin
      top_0[0] = {1'b0,layer_1_0[3319:3312]} - {1'b0, layer_0_0[3319:3312]};
      top_0[1] = {1'b0,layer_1_0[3327:3320]} - {1'b0, layer_0_0[3327:3320]};
      top_0[2] = {1'b0,layer_1_0[3335:3328]} - {1'b0, layer_0_0[3335:3328]};
      top_1[0] = {1'b0,layer_1_1[3319:3312]} - {1'b0, layer_0_1[3319:3312]};
      top_1[1] = {1'b0,layer_1_1[3327:3320]} - {1'b0, layer_0_1[3327:3320]};
      top_1[2] = {1'b0,layer_1_1[3335:3328]} - {1'b0, layer_0_1[3335:3328]};
      top_2[0] = {1'b0,layer_1_2[3319:3312]} - {1'b0, layer_0_2[3319:3312]};
      top_2[1] = {1'b0,layer_1_2[3327:3320]} - {1'b0, layer_0_2[3327:3320]};
      top_2[2] = {1'b0,layer_1_2[3335:3328]} - {1'b0, layer_0_2[3335:3328]};
      mid_0[0] = {1'b0,layer_2_0[3319:3312]} - {1'b0, layer_1_0[3319:3312]};
      mid_0[1] = {1'b0,layer_2_0[3327:3320]} - {1'b0, layer_1_0[3327:3320]};
      mid_0[2] = {1'b0,layer_2_0[3335:3328]} - {1'b0, layer_1_0[3335:3328]};
      mid_1[0] = {1'b0,layer_2_1[3319:3312]} - {1'b0, layer_1_1[3319:3312]};
      mid_1[1] = {1'b0,layer_2_1[3327:3320]} - {1'b0, layer_1_1[3327:3320]};
      mid_1[2] = {1'b0,layer_2_1[3335:3328]} - {1'b0, layer_1_1[3335:3328]};
      mid_2[0] = {1'b0,layer_2_2[3319:3312]} - {1'b0, layer_1_2[3319:3312]};
      mid_2[1] = {1'b0,layer_2_2[3327:3320]} - {1'b0, layer_1_2[3327:3320]};
      mid_2[2] = {1'b0,layer_2_2[3335:3328]} - {1'b0, layer_1_2[3335:3328]};
      btm_0[0] = {1'b0,layer_3_0[3319:3312]} - {1'b0, layer_2_0[3319:3312]};
      btm_0[1] = {1'b0,layer_3_0[3327:3320]} - {1'b0, layer_2_0[3327:3320]};
      btm_0[2] = {1'b0,layer_3_0[3335:3328]} - {1'b0, layer_2_0[3335:3328]};
      btm_1[0] = {1'b0,layer_3_1[3319:3312]} - {1'b0, layer_2_1[3319:3312]};
      btm_1[1] = {1'b0,layer_3_1[3327:3320]} - {1'b0, layer_2_1[3327:3320]};
      btm_1[2] = {1'b0,layer_3_1[3335:3328]} - {1'b0, layer_2_1[3335:3328]};
      btm_2[0] = {1'b0,layer_3_2[3319:3312]} - {1'b0, layer_2_2[3319:3312]};
      btm_2[1] = {1'b0,layer_3_2[3327:3320]} - {1'b0, layer_2_2[3327:3320]};
      btm_2[2] = {1'b0,layer_3_2[3335:3328]} - {1'b0, layer_2_2[3335:3328]};
    end
    'd416: begin
      top_0[0] = {1'b0,layer_1_0[3327:3320]} - {1'b0, layer_0_0[3327:3320]};
      top_0[1] = {1'b0,layer_1_0[3335:3328]} - {1'b0, layer_0_0[3335:3328]};
      top_0[2] = {1'b0,layer_1_0[3343:3336]} - {1'b0, layer_0_0[3343:3336]};
      top_1[0] = {1'b0,layer_1_1[3327:3320]} - {1'b0, layer_0_1[3327:3320]};
      top_1[1] = {1'b0,layer_1_1[3335:3328]} - {1'b0, layer_0_1[3335:3328]};
      top_1[2] = {1'b0,layer_1_1[3343:3336]} - {1'b0, layer_0_1[3343:3336]};
      top_2[0] = {1'b0,layer_1_2[3327:3320]} - {1'b0, layer_0_2[3327:3320]};
      top_2[1] = {1'b0,layer_1_2[3335:3328]} - {1'b0, layer_0_2[3335:3328]};
      top_2[2] = {1'b0,layer_1_2[3343:3336]} - {1'b0, layer_0_2[3343:3336]};
      mid_0[0] = {1'b0,layer_2_0[3327:3320]} - {1'b0, layer_1_0[3327:3320]};
      mid_0[1] = {1'b0,layer_2_0[3335:3328]} - {1'b0, layer_1_0[3335:3328]};
      mid_0[2] = {1'b0,layer_2_0[3343:3336]} - {1'b0, layer_1_0[3343:3336]};
      mid_1[0] = {1'b0,layer_2_1[3327:3320]} - {1'b0, layer_1_1[3327:3320]};
      mid_1[1] = {1'b0,layer_2_1[3335:3328]} - {1'b0, layer_1_1[3335:3328]};
      mid_1[2] = {1'b0,layer_2_1[3343:3336]} - {1'b0, layer_1_1[3343:3336]};
      mid_2[0] = {1'b0,layer_2_2[3327:3320]} - {1'b0, layer_1_2[3327:3320]};
      mid_2[1] = {1'b0,layer_2_2[3335:3328]} - {1'b0, layer_1_2[3335:3328]};
      mid_2[2] = {1'b0,layer_2_2[3343:3336]} - {1'b0, layer_1_2[3343:3336]};
      btm_0[0] = {1'b0,layer_3_0[3327:3320]} - {1'b0, layer_2_0[3327:3320]};
      btm_0[1] = {1'b0,layer_3_0[3335:3328]} - {1'b0, layer_2_0[3335:3328]};
      btm_0[2] = {1'b0,layer_3_0[3343:3336]} - {1'b0, layer_2_0[3343:3336]};
      btm_1[0] = {1'b0,layer_3_1[3327:3320]} - {1'b0, layer_2_1[3327:3320]};
      btm_1[1] = {1'b0,layer_3_1[3335:3328]} - {1'b0, layer_2_1[3335:3328]};
      btm_1[2] = {1'b0,layer_3_1[3343:3336]} - {1'b0, layer_2_1[3343:3336]};
      btm_2[0] = {1'b0,layer_3_2[3327:3320]} - {1'b0, layer_2_2[3327:3320]};
      btm_2[1] = {1'b0,layer_3_2[3335:3328]} - {1'b0, layer_2_2[3335:3328]};
      btm_2[2] = {1'b0,layer_3_2[3343:3336]} - {1'b0, layer_2_2[3343:3336]};
    end
    'd417: begin
      top_0[0] = {1'b0,layer_1_0[3335:3328]} - {1'b0, layer_0_0[3335:3328]};
      top_0[1] = {1'b0,layer_1_0[3343:3336]} - {1'b0, layer_0_0[3343:3336]};
      top_0[2] = {1'b0,layer_1_0[3351:3344]} - {1'b0, layer_0_0[3351:3344]};
      top_1[0] = {1'b0,layer_1_1[3335:3328]} - {1'b0, layer_0_1[3335:3328]};
      top_1[1] = {1'b0,layer_1_1[3343:3336]} - {1'b0, layer_0_1[3343:3336]};
      top_1[2] = {1'b0,layer_1_1[3351:3344]} - {1'b0, layer_0_1[3351:3344]};
      top_2[0] = {1'b0,layer_1_2[3335:3328]} - {1'b0, layer_0_2[3335:3328]};
      top_2[1] = {1'b0,layer_1_2[3343:3336]} - {1'b0, layer_0_2[3343:3336]};
      top_2[2] = {1'b0,layer_1_2[3351:3344]} - {1'b0, layer_0_2[3351:3344]};
      mid_0[0] = {1'b0,layer_2_0[3335:3328]} - {1'b0, layer_1_0[3335:3328]};
      mid_0[1] = {1'b0,layer_2_0[3343:3336]} - {1'b0, layer_1_0[3343:3336]};
      mid_0[2] = {1'b0,layer_2_0[3351:3344]} - {1'b0, layer_1_0[3351:3344]};
      mid_1[0] = {1'b0,layer_2_1[3335:3328]} - {1'b0, layer_1_1[3335:3328]};
      mid_1[1] = {1'b0,layer_2_1[3343:3336]} - {1'b0, layer_1_1[3343:3336]};
      mid_1[2] = {1'b0,layer_2_1[3351:3344]} - {1'b0, layer_1_1[3351:3344]};
      mid_2[0] = {1'b0,layer_2_2[3335:3328]} - {1'b0, layer_1_2[3335:3328]};
      mid_2[1] = {1'b0,layer_2_2[3343:3336]} - {1'b0, layer_1_2[3343:3336]};
      mid_2[2] = {1'b0,layer_2_2[3351:3344]} - {1'b0, layer_1_2[3351:3344]};
      btm_0[0] = {1'b0,layer_3_0[3335:3328]} - {1'b0, layer_2_0[3335:3328]};
      btm_0[1] = {1'b0,layer_3_0[3343:3336]} - {1'b0, layer_2_0[3343:3336]};
      btm_0[2] = {1'b0,layer_3_0[3351:3344]} - {1'b0, layer_2_0[3351:3344]};
      btm_1[0] = {1'b0,layer_3_1[3335:3328]} - {1'b0, layer_2_1[3335:3328]};
      btm_1[1] = {1'b0,layer_3_1[3343:3336]} - {1'b0, layer_2_1[3343:3336]};
      btm_1[2] = {1'b0,layer_3_1[3351:3344]} - {1'b0, layer_2_1[3351:3344]};
      btm_2[0] = {1'b0,layer_3_2[3335:3328]} - {1'b0, layer_2_2[3335:3328]};
      btm_2[1] = {1'b0,layer_3_2[3343:3336]} - {1'b0, layer_2_2[3343:3336]};
      btm_2[2] = {1'b0,layer_3_2[3351:3344]} - {1'b0, layer_2_2[3351:3344]};
    end
    'd418: begin
      top_0[0] = {1'b0,layer_1_0[3343:3336]} - {1'b0, layer_0_0[3343:3336]};
      top_0[1] = {1'b0,layer_1_0[3351:3344]} - {1'b0, layer_0_0[3351:3344]};
      top_0[2] = {1'b0,layer_1_0[3359:3352]} - {1'b0, layer_0_0[3359:3352]};
      top_1[0] = {1'b0,layer_1_1[3343:3336]} - {1'b0, layer_0_1[3343:3336]};
      top_1[1] = {1'b0,layer_1_1[3351:3344]} - {1'b0, layer_0_1[3351:3344]};
      top_1[2] = {1'b0,layer_1_1[3359:3352]} - {1'b0, layer_0_1[3359:3352]};
      top_2[0] = {1'b0,layer_1_2[3343:3336]} - {1'b0, layer_0_2[3343:3336]};
      top_2[1] = {1'b0,layer_1_2[3351:3344]} - {1'b0, layer_0_2[3351:3344]};
      top_2[2] = {1'b0,layer_1_2[3359:3352]} - {1'b0, layer_0_2[3359:3352]};
      mid_0[0] = {1'b0,layer_2_0[3343:3336]} - {1'b0, layer_1_0[3343:3336]};
      mid_0[1] = {1'b0,layer_2_0[3351:3344]} - {1'b0, layer_1_0[3351:3344]};
      mid_0[2] = {1'b0,layer_2_0[3359:3352]} - {1'b0, layer_1_0[3359:3352]};
      mid_1[0] = {1'b0,layer_2_1[3343:3336]} - {1'b0, layer_1_1[3343:3336]};
      mid_1[1] = {1'b0,layer_2_1[3351:3344]} - {1'b0, layer_1_1[3351:3344]};
      mid_1[2] = {1'b0,layer_2_1[3359:3352]} - {1'b0, layer_1_1[3359:3352]};
      mid_2[0] = {1'b0,layer_2_2[3343:3336]} - {1'b0, layer_1_2[3343:3336]};
      mid_2[1] = {1'b0,layer_2_2[3351:3344]} - {1'b0, layer_1_2[3351:3344]};
      mid_2[2] = {1'b0,layer_2_2[3359:3352]} - {1'b0, layer_1_2[3359:3352]};
      btm_0[0] = {1'b0,layer_3_0[3343:3336]} - {1'b0, layer_2_0[3343:3336]};
      btm_0[1] = {1'b0,layer_3_0[3351:3344]} - {1'b0, layer_2_0[3351:3344]};
      btm_0[2] = {1'b0,layer_3_0[3359:3352]} - {1'b0, layer_2_0[3359:3352]};
      btm_1[0] = {1'b0,layer_3_1[3343:3336]} - {1'b0, layer_2_1[3343:3336]};
      btm_1[1] = {1'b0,layer_3_1[3351:3344]} - {1'b0, layer_2_1[3351:3344]};
      btm_1[2] = {1'b0,layer_3_1[3359:3352]} - {1'b0, layer_2_1[3359:3352]};
      btm_2[0] = {1'b0,layer_3_2[3343:3336]} - {1'b0, layer_2_2[3343:3336]};
      btm_2[1] = {1'b0,layer_3_2[3351:3344]} - {1'b0, layer_2_2[3351:3344]};
      btm_2[2] = {1'b0,layer_3_2[3359:3352]} - {1'b0, layer_2_2[3359:3352]};
    end
    'd419: begin
      top_0[0] = {1'b0,layer_1_0[3351:3344]} - {1'b0, layer_0_0[3351:3344]};
      top_0[1] = {1'b0,layer_1_0[3359:3352]} - {1'b0, layer_0_0[3359:3352]};
      top_0[2] = {1'b0,layer_1_0[3367:3360]} - {1'b0, layer_0_0[3367:3360]};
      top_1[0] = {1'b0,layer_1_1[3351:3344]} - {1'b0, layer_0_1[3351:3344]};
      top_1[1] = {1'b0,layer_1_1[3359:3352]} - {1'b0, layer_0_1[3359:3352]};
      top_1[2] = {1'b0,layer_1_1[3367:3360]} - {1'b0, layer_0_1[3367:3360]};
      top_2[0] = {1'b0,layer_1_2[3351:3344]} - {1'b0, layer_0_2[3351:3344]};
      top_2[1] = {1'b0,layer_1_2[3359:3352]} - {1'b0, layer_0_2[3359:3352]};
      top_2[2] = {1'b0,layer_1_2[3367:3360]} - {1'b0, layer_0_2[3367:3360]};
      mid_0[0] = {1'b0,layer_2_0[3351:3344]} - {1'b0, layer_1_0[3351:3344]};
      mid_0[1] = {1'b0,layer_2_0[3359:3352]} - {1'b0, layer_1_0[3359:3352]};
      mid_0[2] = {1'b0,layer_2_0[3367:3360]} - {1'b0, layer_1_0[3367:3360]};
      mid_1[0] = {1'b0,layer_2_1[3351:3344]} - {1'b0, layer_1_1[3351:3344]};
      mid_1[1] = {1'b0,layer_2_1[3359:3352]} - {1'b0, layer_1_1[3359:3352]};
      mid_1[2] = {1'b0,layer_2_1[3367:3360]} - {1'b0, layer_1_1[3367:3360]};
      mid_2[0] = {1'b0,layer_2_2[3351:3344]} - {1'b0, layer_1_2[3351:3344]};
      mid_2[1] = {1'b0,layer_2_2[3359:3352]} - {1'b0, layer_1_2[3359:3352]};
      mid_2[2] = {1'b0,layer_2_2[3367:3360]} - {1'b0, layer_1_2[3367:3360]};
      btm_0[0] = {1'b0,layer_3_0[3351:3344]} - {1'b0, layer_2_0[3351:3344]};
      btm_0[1] = {1'b0,layer_3_0[3359:3352]} - {1'b0, layer_2_0[3359:3352]};
      btm_0[2] = {1'b0,layer_3_0[3367:3360]} - {1'b0, layer_2_0[3367:3360]};
      btm_1[0] = {1'b0,layer_3_1[3351:3344]} - {1'b0, layer_2_1[3351:3344]};
      btm_1[1] = {1'b0,layer_3_1[3359:3352]} - {1'b0, layer_2_1[3359:3352]};
      btm_1[2] = {1'b0,layer_3_1[3367:3360]} - {1'b0, layer_2_1[3367:3360]};
      btm_2[0] = {1'b0,layer_3_2[3351:3344]} - {1'b0, layer_2_2[3351:3344]};
      btm_2[1] = {1'b0,layer_3_2[3359:3352]} - {1'b0, layer_2_2[3359:3352]};
      btm_2[2] = {1'b0,layer_3_2[3367:3360]} - {1'b0, layer_2_2[3367:3360]};
    end
    'd420: begin
      top_0[0] = {1'b0,layer_1_0[3359:3352]} - {1'b0, layer_0_0[3359:3352]};
      top_0[1] = {1'b0,layer_1_0[3367:3360]} - {1'b0, layer_0_0[3367:3360]};
      top_0[2] = {1'b0,layer_1_0[3375:3368]} - {1'b0, layer_0_0[3375:3368]};
      top_1[0] = {1'b0,layer_1_1[3359:3352]} - {1'b0, layer_0_1[3359:3352]};
      top_1[1] = {1'b0,layer_1_1[3367:3360]} - {1'b0, layer_0_1[3367:3360]};
      top_1[2] = {1'b0,layer_1_1[3375:3368]} - {1'b0, layer_0_1[3375:3368]};
      top_2[0] = {1'b0,layer_1_2[3359:3352]} - {1'b0, layer_0_2[3359:3352]};
      top_2[1] = {1'b0,layer_1_2[3367:3360]} - {1'b0, layer_0_2[3367:3360]};
      top_2[2] = {1'b0,layer_1_2[3375:3368]} - {1'b0, layer_0_2[3375:3368]};
      mid_0[0] = {1'b0,layer_2_0[3359:3352]} - {1'b0, layer_1_0[3359:3352]};
      mid_0[1] = {1'b0,layer_2_0[3367:3360]} - {1'b0, layer_1_0[3367:3360]};
      mid_0[2] = {1'b0,layer_2_0[3375:3368]} - {1'b0, layer_1_0[3375:3368]};
      mid_1[0] = {1'b0,layer_2_1[3359:3352]} - {1'b0, layer_1_1[3359:3352]};
      mid_1[1] = {1'b0,layer_2_1[3367:3360]} - {1'b0, layer_1_1[3367:3360]};
      mid_1[2] = {1'b0,layer_2_1[3375:3368]} - {1'b0, layer_1_1[3375:3368]};
      mid_2[0] = {1'b0,layer_2_2[3359:3352]} - {1'b0, layer_1_2[3359:3352]};
      mid_2[1] = {1'b0,layer_2_2[3367:3360]} - {1'b0, layer_1_2[3367:3360]};
      mid_2[2] = {1'b0,layer_2_2[3375:3368]} - {1'b0, layer_1_2[3375:3368]};
      btm_0[0] = {1'b0,layer_3_0[3359:3352]} - {1'b0, layer_2_0[3359:3352]};
      btm_0[1] = {1'b0,layer_3_0[3367:3360]} - {1'b0, layer_2_0[3367:3360]};
      btm_0[2] = {1'b0,layer_3_0[3375:3368]} - {1'b0, layer_2_0[3375:3368]};
      btm_1[0] = {1'b0,layer_3_1[3359:3352]} - {1'b0, layer_2_1[3359:3352]};
      btm_1[1] = {1'b0,layer_3_1[3367:3360]} - {1'b0, layer_2_1[3367:3360]};
      btm_1[2] = {1'b0,layer_3_1[3375:3368]} - {1'b0, layer_2_1[3375:3368]};
      btm_2[0] = {1'b0,layer_3_2[3359:3352]} - {1'b0, layer_2_2[3359:3352]};
      btm_2[1] = {1'b0,layer_3_2[3367:3360]} - {1'b0, layer_2_2[3367:3360]};
      btm_2[2] = {1'b0,layer_3_2[3375:3368]} - {1'b0, layer_2_2[3375:3368]};
    end
    'd421: begin
      top_0[0] = {1'b0,layer_1_0[3367:3360]} - {1'b0, layer_0_0[3367:3360]};
      top_0[1] = {1'b0,layer_1_0[3375:3368]} - {1'b0, layer_0_0[3375:3368]};
      top_0[2] = {1'b0,layer_1_0[3383:3376]} - {1'b0, layer_0_0[3383:3376]};
      top_1[0] = {1'b0,layer_1_1[3367:3360]} - {1'b0, layer_0_1[3367:3360]};
      top_1[1] = {1'b0,layer_1_1[3375:3368]} - {1'b0, layer_0_1[3375:3368]};
      top_1[2] = {1'b0,layer_1_1[3383:3376]} - {1'b0, layer_0_1[3383:3376]};
      top_2[0] = {1'b0,layer_1_2[3367:3360]} - {1'b0, layer_0_2[3367:3360]};
      top_2[1] = {1'b0,layer_1_2[3375:3368]} - {1'b0, layer_0_2[3375:3368]};
      top_2[2] = {1'b0,layer_1_2[3383:3376]} - {1'b0, layer_0_2[3383:3376]};
      mid_0[0] = {1'b0,layer_2_0[3367:3360]} - {1'b0, layer_1_0[3367:3360]};
      mid_0[1] = {1'b0,layer_2_0[3375:3368]} - {1'b0, layer_1_0[3375:3368]};
      mid_0[2] = {1'b0,layer_2_0[3383:3376]} - {1'b0, layer_1_0[3383:3376]};
      mid_1[0] = {1'b0,layer_2_1[3367:3360]} - {1'b0, layer_1_1[3367:3360]};
      mid_1[1] = {1'b0,layer_2_1[3375:3368]} - {1'b0, layer_1_1[3375:3368]};
      mid_1[2] = {1'b0,layer_2_1[3383:3376]} - {1'b0, layer_1_1[3383:3376]};
      mid_2[0] = {1'b0,layer_2_2[3367:3360]} - {1'b0, layer_1_2[3367:3360]};
      mid_2[1] = {1'b0,layer_2_2[3375:3368]} - {1'b0, layer_1_2[3375:3368]};
      mid_2[2] = {1'b0,layer_2_2[3383:3376]} - {1'b0, layer_1_2[3383:3376]};
      btm_0[0] = {1'b0,layer_3_0[3367:3360]} - {1'b0, layer_2_0[3367:3360]};
      btm_0[1] = {1'b0,layer_3_0[3375:3368]} - {1'b0, layer_2_0[3375:3368]};
      btm_0[2] = {1'b0,layer_3_0[3383:3376]} - {1'b0, layer_2_0[3383:3376]};
      btm_1[0] = {1'b0,layer_3_1[3367:3360]} - {1'b0, layer_2_1[3367:3360]};
      btm_1[1] = {1'b0,layer_3_1[3375:3368]} - {1'b0, layer_2_1[3375:3368]};
      btm_1[2] = {1'b0,layer_3_1[3383:3376]} - {1'b0, layer_2_1[3383:3376]};
      btm_2[0] = {1'b0,layer_3_2[3367:3360]} - {1'b0, layer_2_2[3367:3360]};
      btm_2[1] = {1'b0,layer_3_2[3375:3368]} - {1'b0, layer_2_2[3375:3368]};
      btm_2[2] = {1'b0,layer_3_2[3383:3376]} - {1'b0, layer_2_2[3383:3376]};
    end
    'd422: begin
      top_0[0] = {1'b0,layer_1_0[3375:3368]} - {1'b0, layer_0_0[3375:3368]};
      top_0[1] = {1'b0,layer_1_0[3383:3376]} - {1'b0, layer_0_0[3383:3376]};
      top_0[2] = {1'b0,layer_1_0[3391:3384]} - {1'b0, layer_0_0[3391:3384]};
      top_1[0] = {1'b0,layer_1_1[3375:3368]} - {1'b0, layer_0_1[3375:3368]};
      top_1[1] = {1'b0,layer_1_1[3383:3376]} - {1'b0, layer_0_1[3383:3376]};
      top_1[2] = {1'b0,layer_1_1[3391:3384]} - {1'b0, layer_0_1[3391:3384]};
      top_2[0] = {1'b0,layer_1_2[3375:3368]} - {1'b0, layer_0_2[3375:3368]};
      top_2[1] = {1'b0,layer_1_2[3383:3376]} - {1'b0, layer_0_2[3383:3376]};
      top_2[2] = {1'b0,layer_1_2[3391:3384]} - {1'b0, layer_0_2[3391:3384]};
      mid_0[0] = {1'b0,layer_2_0[3375:3368]} - {1'b0, layer_1_0[3375:3368]};
      mid_0[1] = {1'b0,layer_2_0[3383:3376]} - {1'b0, layer_1_0[3383:3376]};
      mid_0[2] = {1'b0,layer_2_0[3391:3384]} - {1'b0, layer_1_0[3391:3384]};
      mid_1[0] = {1'b0,layer_2_1[3375:3368]} - {1'b0, layer_1_1[3375:3368]};
      mid_1[1] = {1'b0,layer_2_1[3383:3376]} - {1'b0, layer_1_1[3383:3376]};
      mid_1[2] = {1'b0,layer_2_1[3391:3384]} - {1'b0, layer_1_1[3391:3384]};
      mid_2[0] = {1'b0,layer_2_2[3375:3368]} - {1'b0, layer_1_2[3375:3368]};
      mid_2[1] = {1'b0,layer_2_2[3383:3376]} - {1'b0, layer_1_2[3383:3376]};
      mid_2[2] = {1'b0,layer_2_2[3391:3384]} - {1'b0, layer_1_2[3391:3384]};
      btm_0[0] = {1'b0,layer_3_0[3375:3368]} - {1'b0, layer_2_0[3375:3368]};
      btm_0[1] = {1'b0,layer_3_0[3383:3376]} - {1'b0, layer_2_0[3383:3376]};
      btm_0[2] = {1'b0,layer_3_0[3391:3384]} - {1'b0, layer_2_0[3391:3384]};
      btm_1[0] = {1'b0,layer_3_1[3375:3368]} - {1'b0, layer_2_1[3375:3368]};
      btm_1[1] = {1'b0,layer_3_1[3383:3376]} - {1'b0, layer_2_1[3383:3376]};
      btm_1[2] = {1'b0,layer_3_1[3391:3384]} - {1'b0, layer_2_1[3391:3384]};
      btm_2[0] = {1'b0,layer_3_2[3375:3368]} - {1'b0, layer_2_2[3375:3368]};
      btm_2[1] = {1'b0,layer_3_2[3383:3376]} - {1'b0, layer_2_2[3383:3376]};
      btm_2[2] = {1'b0,layer_3_2[3391:3384]} - {1'b0, layer_2_2[3391:3384]};
    end
    'd423: begin
      top_0[0] = {1'b0,layer_1_0[3383:3376]} - {1'b0, layer_0_0[3383:3376]};
      top_0[1] = {1'b0,layer_1_0[3391:3384]} - {1'b0, layer_0_0[3391:3384]};
      top_0[2] = {1'b0,layer_1_0[3399:3392]} - {1'b0, layer_0_0[3399:3392]};
      top_1[0] = {1'b0,layer_1_1[3383:3376]} - {1'b0, layer_0_1[3383:3376]};
      top_1[1] = {1'b0,layer_1_1[3391:3384]} - {1'b0, layer_0_1[3391:3384]};
      top_1[2] = {1'b0,layer_1_1[3399:3392]} - {1'b0, layer_0_1[3399:3392]};
      top_2[0] = {1'b0,layer_1_2[3383:3376]} - {1'b0, layer_0_2[3383:3376]};
      top_2[1] = {1'b0,layer_1_2[3391:3384]} - {1'b0, layer_0_2[3391:3384]};
      top_2[2] = {1'b0,layer_1_2[3399:3392]} - {1'b0, layer_0_2[3399:3392]};
      mid_0[0] = {1'b0,layer_2_0[3383:3376]} - {1'b0, layer_1_0[3383:3376]};
      mid_0[1] = {1'b0,layer_2_0[3391:3384]} - {1'b0, layer_1_0[3391:3384]};
      mid_0[2] = {1'b0,layer_2_0[3399:3392]} - {1'b0, layer_1_0[3399:3392]};
      mid_1[0] = {1'b0,layer_2_1[3383:3376]} - {1'b0, layer_1_1[3383:3376]};
      mid_1[1] = {1'b0,layer_2_1[3391:3384]} - {1'b0, layer_1_1[3391:3384]};
      mid_1[2] = {1'b0,layer_2_1[3399:3392]} - {1'b0, layer_1_1[3399:3392]};
      mid_2[0] = {1'b0,layer_2_2[3383:3376]} - {1'b0, layer_1_2[3383:3376]};
      mid_2[1] = {1'b0,layer_2_2[3391:3384]} - {1'b0, layer_1_2[3391:3384]};
      mid_2[2] = {1'b0,layer_2_2[3399:3392]} - {1'b0, layer_1_2[3399:3392]};
      btm_0[0] = {1'b0,layer_3_0[3383:3376]} - {1'b0, layer_2_0[3383:3376]};
      btm_0[1] = {1'b0,layer_3_0[3391:3384]} - {1'b0, layer_2_0[3391:3384]};
      btm_0[2] = {1'b0,layer_3_0[3399:3392]} - {1'b0, layer_2_0[3399:3392]};
      btm_1[0] = {1'b0,layer_3_1[3383:3376]} - {1'b0, layer_2_1[3383:3376]};
      btm_1[1] = {1'b0,layer_3_1[3391:3384]} - {1'b0, layer_2_1[3391:3384]};
      btm_1[2] = {1'b0,layer_3_1[3399:3392]} - {1'b0, layer_2_1[3399:3392]};
      btm_2[0] = {1'b0,layer_3_2[3383:3376]} - {1'b0, layer_2_2[3383:3376]};
      btm_2[1] = {1'b0,layer_3_2[3391:3384]} - {1'b0, layer_2_2[3391:3384]};
      btm_2[2] = {1'b0,layer_3_2[3399:3392]} - {1'b0, layer_2_2[3399:3392]};
    end
    'd424: begin
      top_0[0] = {1'b0,layer_1_0[3391:3384]} - {1'b0, layer_0_0[3391:3384]};
      top_0[1] = {1'b0,layer_1_0[3399:3392]} - {1'b0, layer_0_0[3399:3392]};
      top_0[2] = {1'b0,layer_1_0[3407:3400]} - {1'b0, layer_0_0[3407:3400]};
      top_1[0] = {1'b0,layer_1_1[3391:3384]} - {1'b0, layer_0_1[3391:3384]};
      top_1[1] = {1'b0,layer_1_1[3399:3392]} - {1'b0, layer_0_1[3399:3392]};
      top_1[2] = {1'b0,layer_1_1[3407:3400]} - {1'b0, layer_0_1[3407:3400]};
      top_2[0] = {1'b0,layer_1_2[3391:3384]} - {1'b0, layer_0_2[3391:3384]};
      top_2[1] = {1'b0,layer_1_2[3399:3392]} - {1'b0, layer_0_2[3399:3392]};
      top_2[2] = {1'b0,layer_1_2[3407:3400]} - {1'b0, layer_0_2[3407:3400]};
      mid_0[0] = {1'b0,layer_2_0[3391:3384]} - {1'b0, layer_1_0[3391:3384]};
      mid_0[1] = {1'b0,layer_2_0[3399:3392]} - {1'b0, layer_1_0[3399:3392]};
      mid_0[2] = {1'b0,layer_2_0[3407:3400]} - {1'b0, layer_1_0[3407:3400]};
      mid_1[0] = {1'b0,layer_2_1[3391:3384]} - {1'b0, layer_1_1[3391:3384]};
      mid_1[1] = {1'b0,layer_2_1[3399:3392]} - {1'b0, layer_1_1[3399:3392]};
      mid_1[2] = {1'b0,layer_2_1[3407:3400]} - {1'b0, layer_1_1[3407:3400]};
      mid_2[0] = {1'b0,layer_2_2[3391:3384]} - {1'b0, layer_1_2[3391:3384]};
      mid_2[1] = {1'b0,layer_2_2[3399:3392]} - {1'b0, layer_1_2[3399:3392]};
      mid_2[2] = {1'b0,layer_2_2[3407:3400]} - {1'b0, layer_1_2[3407:3400]};
      btm_0[0] = {1'b0,layer_3_0[3391:3384]} - {1'b0, layer_2_0[3391:3384]};
      btm_0[1] = {1'b0,layer_3_0[3399:3392]} - {1'b0, layer_2_0[3399:3392]};
      btm_0[2] = {1'b0,layer_3_0[3407:3400]} - {1'b0, layer_2_0[3407:3400]};
      btm_1[0] = {1'b0,layer_3_1[3391:3384]} - {1'b0, layer_2_1[3391:3384]};
      btm_1[1] = {1'b0,layer_3_1[3399:3392]} - {1'b0, layer_2_1[3399:3392]};
      btm_1[2] = {1'b0,layer_3_1[3407:3400]} - {1'b0, layer_2_1[3407:3400]};
      btm_2[0] = {1'b0,layer_3_2[3391:3384]} - {1'b0, layer_2_2[3391:3384]};
      btm_2[1] = {1'b0,layer_3_2[3399:3392]} - {1'b0, layer_2_2[3399:3392]};
      btm_2[2] = {1'b0,layer_3_2[3407:3400]} - {1'b0, layer_2_2[3407:3400]};
    end
    'd425: begin
      top_0[0] = {1'b0,layer_1_0[3399:3392]} - {1'b0, layer_0_0[3399:3392]};
      top_0[1] = {1'b0,layer_1_0[3407:3400]} - {1'b0, layer_0_0[3407:3400]};
      top_0[2] = {1'b0,layer_1_0[3415:3408]} - {1'b0, layer_0_0[3415:3408]};
      top_1[0] = {1'b0,layer_1_1[3399:3392]} - {1'b0, layer_0_1[3399:3392]};
      top_1[1] = {1'b0,layer_1_1[3407:3400]} - {1'b0, layer_0_1[3407:3400]};
      top_1[2] = {1'b0,layer_1_1[3415:3408]} - {1'b0, layer_0_1[3415:3408]};
      top_2[0] = {1'b0,layer_1_2[3399:3392]} - {1'b0, layer_0_2[3399:3392]};
      top_2[1] = {1'b0,layer_1_2[3407:3400]} - {1'b0, layer_0_2[3407:3400]};
      top_2[2] = {1'b0,layer_1_2[3415:3408]} - {1'b0, layer_0_2[3415:3408]};
      mid_0[0] = {1'b0,layer_2_0[3399:3392]} - {1'b0, layer_1_0[3399:3392]};
      mid_0[1] = {1'b0,layer_2_0[3407:3400]} - {1'b0, layer_1_0[3407:3400]};
      mid_0[2] = {1'b0,layer_2_0[3415:3408]} - {1'b0, layer_1_0[3415:3408]};
      mid_1[0] = {1'b0,layer_2_1[3399:3392]} - {1'b0, layer_1_1[3399:3392]};
      mid_1[1] = {1'b0,layer_2_1[3407:3400]} - {1'b0, layer_1_1[3407:3400]};
      mid_1[2] = {1'b0,layer_2_1[3415:3408]} - {1'b0, layer_1_1[3415:3408]};
      mid_2[0] = {1'b0,layer_2_2[3399:3392]} - {1'b0, layer_1_2[3399:3392]};
      mid_2[1] = {1'b0,layer_2_2[3407:3400]} - {1'b0, layer_1_2[3407:3400]};
      mid_2[2] = {1'b0,layer_2_2[3415:3408]} - {1'b0, layer_1_2[3415:3408]};
      btm_0[0] = {1'b0,layer_3_0[3399:3392]} - {1'b0, layer_2_0[3399:3392]};
      btm_0[1] = {1'b0,layer_3_0[3407:3400]} - {1'b0, layer_2_0[3407:3400]};
      btm_0[2] = {1'b0,layer_3_0[3415:3408]} - {1'b0, layer_2_0[3415:3408]};
      btm_1[0] = {1'b0,layer_3_1[3399:3392]} - {1'b0, layer_2_1[3399:3392]};
      btm_1[1] = {1'b0,layer_3_1[3407:3400]} - {1'b0, layer_2_1[3407:3400]};
      btm_1[2] = {1'b0,layer_3_1[3415:3408]} - {1'b0, layer_2_1[3415:3408]};
      btm_2[0] = {1'b0,layer_3_2[3399:3392]} - {1'b0, layer_2_2[3399:3392]};
      btm_2[1] = {1'b0,layer_3_2[3407:3400]} - {1'b0, layer_2_2[3407:3400]};
      btm_2[2] = {1'b0,layer_3_2[3415:3408]} - {1'b0, layer_2_2[3415:3408]};
    end
    'd426: begin
      top_0[0] = {1'b0,layer_1_0[3407:3400]} - {1'b0, layer_0_0[3407:3400]};
      top_0[1] = {1'b0,layer_1_0[3415:3408]} - {1'b0, layer_0_0[3415:3408]};
      top_0[2] = {1'b0,layer_1_0[3423:3416]} - {1'b0, layer_0_0[3423:3416]};
      top_1[0] = {1'b0,layer_1_1[3407:3400]} - {1'b0, layer_0_1[3407:3400]};
      top_1[1] = {1'b0,layer_1_1[3415:3408]} - {1'b0, layer_0_1[3415:3408]};
      top_1[2] = {1'b0,layer_1_1[3423:3416]} - {1'b0, layer_0_1[3423:3416]};
      top_2[0] = {1'b0,layer_1_2[3407:3400]} - {1'b0, layer_0_2[3407:3400]};
      top_2[1] = {1'b0,layer_1_2[3415:3408]} - {1'b0, layer_0_2[3415:3408]};
      top_2[2] = {1'b0,layer_1_2[3423:3416]} - {1'b0, layer_0_2[3423:3416]};
      mid_0[0] = {1'b0,layer_2_0[3407:3400]} - {1'b0, layer_1_0[3407:3400]};
      mid_0[1] = {1'b0,layer_2_0[3415:3408]} - {1'b0, layer_1_0[3415:3408]};
      mid_0[2] = {1'b0,layer_2_0[3423:3416]} - {1'b0, layer_1_0[3423:3416]};
      mid_1[0] = {1'b0,layer_2_1[3407:3400]} - {1'b0, layer_1_1[3407:3400]};
      mid_1[1] = {1'b0,layer_2_1[3415:3408]} - {1'b0, layer_1_1[3415:3408]};
      mid_1[2] = {1'b0,layer_2_1[3423:3416]} - {1'b0, layer_1_1[3423:3416]};
      mid_2[0] = {1'b0,layer_2_2[3407:3400]} - {1'b0, layer_1_2[3407:3400]};
      mid_2[1] = {1'b0,layer_2_2[3415:3408]} - {1'b0, layer_1_2[3415:3408]};
      mid_2[2] = {1'b0,layer_2_2[3423:3416]} - {1'b0, layer_1_2[3423:3416]};
      btm_0[0] = {1'b0,layer_3_0[3407:3400]} - {1'b0, layer_2_0[3407:3400]};
      btm_0[1] = {1'b0,layer_3_0[3415:3408]} - {1'b0, layer_2_0[3415:3408]};
      btm_0[2] = {1'b0,layer_3_0[3423:3416]} - {1'b0, layer_2_0[3423:3416]};
      btm_1[0] = {1'b0,layer_3_1[3407:3400]} - {1'b0, layer_2_1[3407:3400]};
      btm_1[1] = {1'b0,layer_3_1[3415:3408]} - {1'b0, layer_2_1[3415:3408]};
      btm_1[2] = {1'b0,layer_3_1[3423:3416]} - {1'b0, layer_2_1[3423:3416]};
      btm_2[0] = {1'b0,layer_3_2[3407:3400]} - {1'b0, layer_2_2[3407:3400]};
      btm_2[1] = {1'b0,layer_3_2[3415:3408]} - {1'b0, layer_2_2[3415:3408]};
      btm_2[2] = {1'b0,layer_3_2[3423:3416]} - {1'b0, layer_2_2[3423:3416]};
    end
    'd427: begin
      top_0[0] = {1'b0,layer_1_0[3415:3408]} - {1'b0, layer_0_0[3415:3408]};
      top_0[1] = {1'b0,layer_1_0[3423:3416]} - {1'b0, layer_0_0[3423:3416]};
      top_0[2] = {1'b0,layer_1_0[3431:3424]} - {1'b0, layer_0_0[3431:3424]};
      top_1[0] = {1'b0,layer_1_1[3415:3408]} - {1'b0, layer_0_1[3415:3408]};
      top_1[1] = {1'b0,layer_1_1[3423:3416]} - {1'b0, layer_0_1[3423:3416]};
      top_1[2] = {1'b0,layer_1_1[3431:3424]} - {1'b0, layer_0_1[3431:3424]};
      top_2[0] = {1'b0,layer_1_2[3415:3408]} - {1'b0, layer_0_2[3415:3408]};
      top_2[1] = {1'b0,layer_1_2[3423:3416]} - {1'b0, layer_0_2[3423:3416]};
      top_2[2] = {1'b0,layer_1_2[3431:3424]} - {1'b0, layer_0_2[3431:3424]};
      mid_0[0] = {1'b0,layer_2_0[3415:3408]} - {1'b0, layer_1_0[3415:3408]};
      mid_0[1] = {1'b0,layer_2_0[3423:3416]} - {1'b0, layer_1_0[3423:3416]};
      mid_0[2] = {1'b0,layer_2_0[3431:3424]} - {1'b0, layer_1_0[3431:3424]};
      mid_1[0] = {1'b0,layer_2_1[3415:3408]} - {1'b0, layer_1_1[3415:3408]};
      mid_1[1] = {1'b0,layer_2_1[3423:3416]} - {1'b0, layer_1_1[3423:3416]};
      mid_1[2] = {1'b0,layer_2_1[3431:3424]} - {1'b0, layer_1_1[3431:3424]};
      mid_2[0] = {1'b0,layer_2_2[3415:3408]} - {1'b0, layer_1_2[3415:3408]};
      mid_2[1] = {1'b0,layer_2_2[3423:3416]} - {1'b0, layer_1_2[3423:3416]};
      mid_2[2] = {1'b0,layer_2_2[3431:3424]} - {1'b0, layer_1_2[3431:3424]};
      btm_0[0] = {1'b0,layer_3_0[3415:3408]} - {1'b0, layer_2_0[3415:3408]};
      btm_0[1] = {1'b0,layer_3_0[3423:3416]} - {1'b0, layer_2_0[3423:3416]};
      btm_0[2] = {1'b0,layer_3_0[3431:3424]} - {1'b0, layer_2_0[3431:3424]};
      btm_1[0] = {1'b0,layer_3_1[3415:3408]} - {1'b0, layer_2_1[3415:3408]};
      btm_1[1] = {1'b0,layer_3_1[3423:3416]} - {1'b0, layer_2_1[3423:3416]};
      btm_1[2] = {1'b0,layer_3_1[3431:3424]} - {1'b0, layer_2_1[3431:3424]};
      btm_2[0] = {1'b0,layer_3_2[3415:3408]} - {1'b0, layer_2_2[3415:3408]};
      btm_2[1] = {1'b0,layer_3_2[3423:3416]} - {1'b0, layer_2_2[3423:3416]};
      btm_2[2] = {1'b0,layer_3_2[3431:3424]} - {1'b0, layer_2_2[3431:3424]};
    end
    'd428: begin
      top_0[0] = {1'b0,layer_1_0[3423:3416]} - {1'b0, layer_0_0[3423:3416]};
      top_0[1] = {1'b0,layer_1_0[3431:3424]} - {1'b0, layer_0_0[3431:3424]};
      top_0[2] = {1'b0,layer_1_0[3439:3432]} - {1'b0, layer_0_0[3439:3432]};
      top_1[0] = {1'b0,layer_1_1[3423:3416]} - {1'b0, layer_0_1[3423:3416]};
      top_1[1] = {1'b0,layer_1_1[3431:3424]} - {1'b0, layer_0_1[3431:3424]};
      top_1[2] = {1'b0,layer_1_1[3439:3432]} - {1'b0, layer_0_1[3439:3432]};
      top_2[0] = {1'b0,layer_1_2[3423:3416]} - {1'b0, layer_0_2[3423:3416]};
      top_2[1] = {1'b0,layer_1_2[3431:3424]} - {1'b0, layer_0_2[3431:3424]};
      top_2[2] = {1'b0,layer_1_2[3439:3432]} - {1'b0, layer_0_2[3439:3432]};
      mid_0[0] = {1'b0,layer_2_0[3423:3416]} - {1'b0, layer_1_0[3423:3416]};
      mid_0[1] = {1'b0,layer_2_0[3431:3424]} - {1'b0, layer_1_0[3431:3424]};
      mid_0[2] = {1'b0,layer_2_0[3439:3432]} - {1'b0, layer_1_0[3439:3432]};
      mid_1[0] = {1'b0,layer_2_1[3423:3416]} - {1'b0, layer_1_1[3423:3416]};
      mid_1[1] = {1'b0,layer_2_1[3431:3424]} - {1'b0, layer_1_1[3431:3424]};
      mid_1[2] = {1'b0,layer_2_1[3439:3432]} - {1'b0, layer_1_1[3439:3432]};
      mid_2[0] = {1'b0,layer_2_2[3423:3416]} - {1'b0, layer_1_2[3423:3416]};
      mid_2[1] = {1'b0,layer_2_2[3431:3424]} - {1'b0, layer_1_2[3431:3424]};
      mid_2[2] = {1'b0,layer_2_2[3439:3432]} - {1'b0, layer_1_2[3439:3432]};
      btm_0[0] = {1'b0,layer_3_0[3423:3416]} - {1'b0, layer_2_0[3423:3416]};
      btm_0[1] = {1'b0,layer_3_0[3431:3424]} - {1'b0, layer_2_0[3431:3424]};
      btm_0[2] = {1'b0,layer_3_0[3439:3432]} - {1'b0, layer_2_0[3439:3432]};
      btm_1[0] = {1'b0,layer_3_1[3423:3416]} - {1'b0, layer_2_1[3423:3416]};
      btm_1[1] = {1'b0,layer_3_1[3431:3424]} - {1'b0, layer_2_1[3431:3424]};
      btm_1[2] = {1'b0,layer_3_1[3439:3432]} - {1'b0, layer_2_1[3439:3432]};
      btm_2[0] = {1'b0,layer_3_2[3423:3416]} - {1'b0, layer_2_2[3423:3416]};
      btm_2[1] = {1'b0,layer_3_2[3431:3424]} - {1'b0, layer_2_2[3431:3424]};
      btm_2[2] = {1'b0,layer_3_2[3439:3432]} - {1'b0, layer_2_2[3439:3432]};
    end
    'd429: begin
      top_0[0] = {1'b0,layer_1_0[3431:3424]} - {1'b0, layer_0_0[3431:3424]};
      top_0[1] = {1'b0,layer_1_0[3439:3432]} - {1'b0, layer_0_0[3439:3432]};
      top_0[2] = {1'b0,layer_1_0[3447:3440]} - {1'b0, layer_0_0[3447:3440]};
      top_1[0] = {1'b0,layer_1_1[3431:3424]} - {1'b0, layer_0_1[3431:3424]};
      top_1[1] = {1'b0,layer_1_1[3439:3432]} - {1'b0, layer_0_1[3439:3432]};
      top_1[2] = {1'b0,layer_1_1[3447:3440]} - {1'b0, layer_0_1[3447:3440]};
      top_2[0] = {1'b0,layer_1_2[3431:3424]} - {1'b0, layer_0_2[3431:3424]};
      top_2[1] = {1'b0,layer_1_2[3439:3432]} - {1'b0, layer_0_2[3439:3432]};
      top_2[2] = {1'b0,layer_1_2[3447:3440]} - {1'b0, layer_0_2[3447:3440]};
      mid_0[0] = {1'b0,layer_2_0[3431:3424]} - {1'b0, layer_1_0[3431:3424]};
      mid_0[1] = {1'b0,layer_2_0[3439:3432]} - {1'b0, layer_1_0[3439:3432]};
      mid_0[2] = {1'b0,layer_2_0[3447:3440]} - {1'b0, layer_1_0[3447:3440]};
      mid_1[0] = {1'b0,layer_2_1[3431:3424]} - {1'b0, layer_1_1[3431:3424]};
      mid_1[1] = {1'b0,layer_2_1[3439:3432]} - {1'b0, layer_1_1[3439:3432]};
      mid_1[2] = {1'b0,layer_2_1[3447:3440]} - {1'b0, layer_1_1[3447:3440]};
      mid_2[0] = {1'b0,layer_2_2[3431:3424]} - {1'b0, layer_1_2[3431:3424]};
      mid_2[1] = {1'b0,layer_2_2[3439:3432]} - {1'b0, layer_1_2[3439:3432]};
      mid_2[2] = {1'b0,layer_2_2[3447:3440]} - {1'b0, layer_1_2[3447:3440]};
      btm_0[0] = {1'b0,layer_3_0[3431:3424]} - {1'b0, layer_2_0[3431:3424]};
      btm_0[1] = {1'b0,layer_3_0[3439:3432]} - {1'b0, layer_2_0[3439:3432]};
      btm_0[2] = {1'b0,layer_3_0[3447:3440]} - {1'b0, layer_2_0[3447:3440]};
      btm_1[0] = {1'b0,layer_3_1[3431:3424]} - {1'b0, layer_2_1[3431:3424]};
      btm_1[1] = {1'b0,layer_3_1[3439:3432]} - {1'b0, layer_2_1[3439:3432]};
      btm_1[2] = {1'b0,layer_3_1[3447:3440]} - {1'b0, layer_2_1[3447:3440]};
      btm_2[0] = {1'b0,layer_3_2[3431:3424]} - {1'b0, layer_2_2[3431:3424]};
      btm_2[1] = {1'b0,layer_3_2[3439:3432]} - {1'b0, layer_2_2[3439:3432]};
      btm_2[2] = {1'b0,layer_3_2[3447:3440]} - {1'b0, layer_2_2[3447:3440]};
    end
    'd430: begin
      top_0[0] = {1'b0,layer_1_0[3439:3432]} - {1'b0, layer_0_0[3439:3432]};
      top_0[1] = {1'b0,layer_1_0[3447:3440]} - {1'b0, layer_0_0[3447:3440]};
      top_0[2] = {1'b0,layer_1_0[3455:3448]} - {1'b0, layer_0_0[3455:3448]};
      top_1[0] = {1'b0,layer_1_1[3439:3432]} - {1'b0, layer_0_1[3439:3432]};
      top_1[1] = {1'b0,layer_1_1[3447:3440]} - {1'b0, layer_0_1[3447:3440]};
      top_1[2] = {1'b0,layer_1_1[3455:3448]} - {1'b0, layer_0_1[3455:3448]};
      top_2[0] = {1'b0,layer_1_2[3439:3432]} - {1'b0, layer_0_2[3439:3432]};
      top_2[1] = {1'b0,layer_1_2[3447:3440]} - {1'b0, layer_0_2[3447:3440]};
      top_2[2] = {1'b0,layer_1_2[3455:3448]} - {1'b0, layer_0_2[3455:3448]};
      mid_0[0] = {1'b0,layer_2_0[3439:3432]} - {1'b0, layer_1_0[3439:3432]};
      mid_0[1] = {1'b0,layer_2_0[3447:3440]} - {1'b0, layer_1_0[3447:3440]};
      mid_0[2] = {1'b0,layer_2_0[3455:3448]} - {1'b0, layer_1_0[3455:3448]};
      mid_1[0] = {1'b0,layer_2_1[3439:3432]} - {1'b0, layer_1_1[3439:3432]};
      mid_1[1] = {1'b0,layer_2_1[3447:3440]} - {1'b0, layer_1_1[3447:3440]};
      mid_1[2] = {1'b0,layer_2_1[3455:3448]} - {1'b0, layer_1_1[3455:3448]};
      mid_2[0] = {1'b0,layer_2_2[3439:3432]} - {1'b0, layer_1_2[3439:3432]};
      mid_2[1] = {1'b0,layer_2_2[3447:3440]} - {1'b0, layer_1_2[3447:3440]};
      mid_2[2] = {1'b0,layer_2_2[3455:3448]} - {1'b0, layer_1_2[3455:3448]};
      btm_0[0] = {1'b0,layer_3_0[3439:3432]} - {1'b0, layer_2_0[3439:3432]};
      btm_0[1] = {1'b0,layer_3_0[3447:3440]} - {1'b0, layer_2_0[3447:3440]};
      btm_0[2] = {1'b0,layer_3_0[3455:3448]} - {1'b0, layer_2_0[3455:3448]};
      btm_1[0] = {1'b0,layer_3_1[3439:3432]} - {1'b0, layer_2_1[3439:3432]};
      btm_1[1] = {1'b0,layer_3_1[3447:3440]} - {1'b0, layer_2_1[3447:3440]};
      btm_1[2] = {1'b0,layer_3_1[3455:3448]} - {1'b0, layer_2_1[3455:3448]};
      btm_2[0] = {1'b0,layer_3_2[3439:3432]} - {1'b0, layer_2_2[3439:3432]};
      btm_2[1] = {1'b0,layer_3_2[3447:3440]} - {1'b0, layer_2_2[3447:3440]};
      btm_2[2] = {1'b0,layer_3_2[3455:3448]} - {1'b0, layer_2_2[3455:3448]};
    end
    'd431: begin
      top_0[0] = {1'b0,layer_1_0[3447:3440]} - {1'b0, layer_0_0[3447:3440]};
      top_0[1] = {1'b0,layer_1_0[3455:3448]} - {1'b0, layer_0_0[3455:3448]};
      top_0[2] = {1'b0,layer_1_0[3463:3456]} - {1'b0, layer_0_0[3463:3456]};
      top_1[0] = {1'b0,layer_1_1[3447:3440]} - {1'b0, layer_0_1[3447:3440]};
      top_1[1] = {1'b0,layer_1_1[3455:3448]} - {1'b0, layer_0_1[3455:3448]};
      top_1[2] = {1'b0,layer_1_1[3463:3456]} - {1'b0, layer_0_1[3463:3456]};
      top_2[0] = {1'b0,layer_1_2[3447:3440]} - {1'b0, layer_0_2[3447:3440]};
      top_2[1] = {1'b0,layer_1_2[3455:3448]} - {1'b0, layer_0_2[3455:3448]};
      top_2[2] = {1'b0,layer_1_2[3463:3456]} - {1'b0, layer_0_2[3463:3456]};
      mid_0[0] = {1'b0,layer_2_0[3447:3440]} - {1'b0, layer_1_0[3447:3440]};
      mid_0[1] = {1'b0,layer_2_0[3455:3448]} - {1'b0, layer_1_0[3455:3448]};
      mid_0[2] = {1'b0,layer_2_0[3463:3456]} - {1'b0, layer_1_0[3463:3456]};
      mid_1[0] = {1'b0,layer_2_1[3447:3440]} - {1'b0, layer_1_1[3447:3440]};
      mid_1[1] = {1'b0,layer_2_1[3455:3448]} - {1'b0, layer_1_1[3455:3448]};
      mid_1[2] = {1'b0,layer_2_1[3463:3456]} - {1'b0, layer_1_1[3463:3456]};
      mid_2[0] = {1'b0,layer_2_2[3447:3440]} - {1'b0, layer_1_2[3447:3440]};
      mid_2[1] = {1'b0,layer_2_2[3455:3448]} - {1'b0, layer_1_2[3455:3448]};
      mid_2[2] = {1'b0,layer_2_2[3463:3456]} - {1'b0, layer_1_2[3463:3456]};
      btm_0[0] = {1'b0,layer_3_0[3447:3440]} - {1'b0, layer_2_0[3447:3440]};
      btm_0[1] = {1'b0,layer_3_0[3455:3448]} - {1'b0, layer_2_0[3455:3448]};
      btm_0[2] = {1'b0,layer_3_0[3463:3456]} - {1'b0, layer_2_0[3463:3456]};
      btm_1[0] = {1'b0,layer_3_1[3447:3440]} - {1'b0, layer_2_1[3447:3440]};
      btm_1[1] = {1'b0,layer_3_1[3455:3448]} - {1'b0, layer_2_1[3455:3448]};
      btm_1[2] = {1'b0,layer_3_1[3463:3456]} - {1'b0, layer_2_1[3463:3456]};
      btm_2[0] = {1'b0,layer_3_2[3447:3440]} - {1'b0, layer_2_2[3447:3440]};
      btm_2[1] = {1'b0,layer_3_2[3455:3448]} - {1'b0, layer_2_2[3455:3448]};
      btm_2[2] = {1'b0,layer_3_2[3463:3456]} - {1'b0, layer_2_2[3463:3456]};
    end
    'd432: begin
      top_0[0] = {1'b0,layer_1_0[3455:3448]} - {1'b0, layer_0_0[3455:3448]};
      top_0[1] = {1'b0,layer_1_0[3463:3456]} - {1'b0, layer_0_0[3463:3456]};
      top_0[2] = {1'b0,layer_1_0[3471:3464]} - {1'b0, layer_0_0[3471:3464]};
      top_1[0] = {1'b0,layer_1_1[3455:3448]} - {1'b0, layer_0_1[3455:3448]};
      top_1[1] = {1'b0,layer_1_1[3463:3456]} - {1'b0, layer_0_1[3463:3456]};
      top_1[2] = {1'b0,layer_1_1[3471:3464]} - {1'b0, layer_0_1[3471:3464]};
      top_2[0] = {1'b0,layer_1_2[3455:3448]} - {1'b0, layer_0_2[3455:3448]};
      top_2[1] = {1'b0,layer_1_2[3463:3456]} - {1'b0, layer_0_2[3463:3456]};
      top_2[2] = {1'b0,layer_1_2[3471:3464]} - {1'b0, layer_0_2[3471:3464]};
      mid_0[0] = {1'b0,layer_2_0[3455:3448]} - {1'b0, layer_1_0[3455:3448]};
      mid_0[1] = {1'b0,layer_2_0[3463:3456]} - {1'b0, layer_1_0[3463:3456]};
      mid_0[2] = {1'b0,layer_2_0[3471:3464]} - {1'b0, layer_1_0[3471:3464]};
      mid_1[0] = {1'b0,layer_2_1[3455:3448]} - {1'b0, layer_1_1[3455:3448]};
      mid_1[1] = {1'b0,layer_2_1[3463:3456]} - {1'b0, layer_1_1[3463:3456]};
      mid_1[2] = {1'b0,layer_2_1[3471:3464]} - {1'b0, layer_1_1[3471:3464]};
      mid_2[0] = {1'b0,layer_2_2[3455:3448]} - {1'b0, layer_1_2[3455:3448]};
      mid_2[1] = {1'b0,layer_2_2[3463:3456]} - {1'b0, layer_1_2[3463:3456]};
      mid_2[2] = {1'b0,layer_2_2[3471:3464]} - {1'b0, layer_1_2[3471:3464]};
      btm_0[0] = {1'b0,layer_3_0[3455:3448]} - {1'b0, layer_2_0[3455:3448]};
      btm_0[1] = {1'b0,layer_3_0[3463:3456]} - {1'b0, layer_2_0[3463:3456]};
      btm_0[2] = {1'b0,layer_3_0[3471:3464]} - {1'b0, layer_2_0[3471:3464]};
      btm_1[0] = {1'b0,layer_3_1[3455:3448]} - {1'b0, layer_2_1[3455:3448]};
      btm_1[1] = {1'b0,layer_3_1[3463:3456]} - {1'b0, layer_2_1[3463:3456]};
      btm_1[2] = {1'b0,layer_3_1[3471:3464]} - {1'b0, layer_2_1[3471:3464]};
      btm_2[0] = {1'b0,layer_3_2[3455:3448]} - {1'b0, layer_2_2[3455:3448]};
      btm_2[1] = {1'b0,layer_3_2[3463:3456]} - {1'b0, layer_2_2[3463:3456]};
      btm_2[2] = {1'b0,layer_3_2[3471:3464]} - {1'b0, layer_2_2[3471:3464]};
    end
    'd433: begin
      top_0[0] = {1'b0,layer_1_0[3463:3456]} - {1'b0, layer_0_0[3463:3456]};
      top_0[1] = {1'b0,layer_1_0[3471:3464]} - {1'b0, layer_0_0[3471:3464]};
      top_0[2] = {1'b0,layer_1_0[3479:3472]} - {1'b0, layer_0_0[3479:3472]};
      top_1[0] = {1'b0,layer_1_1[3463:3456]} - {1'b0, layer_0_1[3463:3456]};
      top_1[1] = {1'b0,layer_1_1[3471:3464]} - {1'b0, layer_0_1[3471:3464]};
      top_1[2] = {1'b0,layer_1_1[3479:3472]} - {1'b0, layer_0_1[3479:3472]};
      top_2[0] = {1'b0,layer_1_2[3463:3456]} - {1'b0, layer_0_2[3463:3456]};
      top_2[1] = {1'b0,layer_1_2[3471:3464]} - {1'b0, layer_0_2[3471:3464]};
      top_2[2] = {1'b0,layer_1_2[3479:3472]} - {1'b0, layer_0_2[3479:3472]};
      mid_0[0] = {1'b0,layer_2_0[3463:3456]} - {1'b0, layer_1_0[3463:3456]};
      mid_0[1] = {1'b0,layer_2_0[3471:3464]} - {1'b0, layer_1_0[3471:3464]};
      mid_0[2] = {1'b0,layer_2_0[3479:3472]} - {1'b0, layer_1_0[3479:3472]};
      mid_1[0] = {1'b0,layer_2_1[3463:3456]} - {1'b0, layer_1_1[3463:3456]};
      mid_1[1] = {1'b0,layer_2_1[3471:3464]} - {1'b0, layer_1_1[3471:3464]};
      mid_1[2] = {1'b0,layer_2_1[3479:3472]} - {1'b0, layer_1_1[3479:3472]};
      mid_2[0] = {1'b0,layer_2_2[3463:3456]} - {1'b0, layer_1_2[3463:3456]};
      mid_2[1] = {1'b0,layer_2_2[3471:3464]} - {1'b0, layer_1_2[3471:3464]};
      mid_2[2] = {1'b0,layer_2_2[3479:3472]} - {1'b0, layer_1_2[3479:3472]};
      btm_0[0] = {1'b0,layer_3_0[3463:3456]} - {1'b0, layer_2_0[3463:3456]};
      btm_0[1] = {1'b0,layer_3_0[3471:3464]} - {1'b0, layer_2_0[3471:3464]};
      btm_0[2] = {1'b0,layer_3_0[3479:3472]} - {1'b0, layer_2_0[3479:3472]};
      btm_1[0] = {1'b0,layer_3_1[3463:3456]} - {1'b0, layer_2_1[3463:3456]};
      btm_1[1] = {1'b0,layer_3_1[3471:3464]} - {1'b0, layer_2_1[3471:3464]};
      btm_1[2] = {1'b0,layer_3_1[3479:3472]} - {1'b0, layer_2_1[3479:3472]};
      btm_2[0] = {1'b0,layer_3_2[3463:3456]} - {1'b0, layer_2_2[3463:3456]};
      btm_2[1] = {1'b0,layer_3_2[3471:3464]} - {1'b0, layer_2_2[3471:3464]};
      btm_2[2] = {1'b0,layer_3_2[3479:3472]} - {1'b0, layer_2_2[3479:3472]};
    end
    'd434: begin
      top_0[0] = {1'b0,layer_1_0[3471:3464]} - {1'b0, layer_0_0[3471:3464]};
      top_0[1] = {1'b0,layer_1_0[3479:3472]} - {1'b0, layer_0_0[3479:3472]};
      top_0[2] = {1'b0,layer_1_0[3487:3480]} - {1'b0, layer_0_0[3487:3480]};
      top_1[0] = {1'b0,layer_1_1[3471:3464]} - {1'b0, layer_0_1[3471:3464]};
      top_1[1] = {1'b0,layer_1_1[3479:3472]} - {1'b0, layer_0_1[3479:3472]};
      top_1[2] = {1'b0,layer_1_1[3487:3480]} - {1'b0, layer_0_1[3487:3480]};
      top_2[0] = {1'b0,layer_1_2[3471:3464]} - {1'b0, layer_0_2[3471:3464]};
      top_2[1] = {1'b0,layer_1_2[3479:3472]} - {1'b0, layer_0_2[3479:3472]};
      top_2[2] = {1'b0,layer_1_2[3487:3480]} - {1'b0, layer_0_2[3487:3480]};
      mid_0[0] = {1'b0,layer_2_0[3471:3464]} - {1'b0, layer_1_0[3471:3464]};
      mid_0[1] = {1'b0,layer_2_0[3479:3472]} - {1'b0, layer_1_0[3479:3472]};
      mid_0[2] = {1'b0,layer_2_0[3487:3480]} - {1'b0, layer_1_0[3487:3480]};
      mid_1[0] = {1'b0,layer_2_1[3471:3464]} - {1'b0, layer_1_1[3471:3464]};
      mid_1[1] = {1'b0,layer_2_1[3479:3472]} - {1'b0, layer_1_1[3479:3472]};
      mid_1[2] = {1'b0,layer_2_1[3487:3480]} - {1'b0, layer_1_1[3487:3480]};
      mid_2[0] = {1'b0,layer_2_2[3471:3464]} - {1'b0, layer_1_2[3471:3464]};
      mid_2[1] = {1'b0,layer_2_2[3479:3472]} - {1'b0, layer_1_2[3479:3472]};
      mid_2[2] = {1'b0,layer_2_2[3487:3480]} - {1'b0, layer_1_2[3487:3480]};
      btm_0[0] = {1'b0,layer_3_0[3471:3464]} - {1'b0, layer_2_0[3471:3464]};
      btm_0[1] = {1'b0,layer_3_0[3479:3472]} - {1'b0, layer_2_0[3479:3472]};
      btm_0[2] = {1'b0,layer_3_0[3487:3480]} - {1'b0, layer_2_0[3487:3480]};
      btm_1[0] = {1'b0,layer_3_1[3471:3464]} - {1'b0, layer_2_1[3471:3464]};
      btm_1[1] = {1'b0,layer_3_1[3479:3472]} - {1'b0, layer_2_1[3479:3472]};
      btm_1[2] = {1'b0,layer_3_1[3487:3480]} - {1'b0, layer_2_1[3487:3480]};
      btm_2[0] = {1'b0,layer_3_2[3471:3464]} - {1'b0, layer_2_2[3471:3464]};
      btm_2[1] = {1'b0,layer_3_2[3479:3472]} - {1'b0, layer_2_2[3479:3472]};
      btm_2[2] = {1'b0,layer_3_2[3487:3480]} - {1'b0, layer_2_2[3487:3480]};
    end
    'd435: begin
      top_0[0] = {1'b0,layer_1_0[3479:3472]} - {1'b0, layer_0_0[3479:3472]};
      top_0[1] = {1'b0,layer_1_0[3487:3480]} - {1'b0, layer_0_0[3487:3480]};
      top_0[2] = {1'b0,layer_1_0[3495:3488]} - {1'b0, layer_0_0[3495:3488]};
      top_1[0] = {1'b0,layer_1_1[3479:3472]} - {1'b0, layer_0_1[3479:3472]};
      top_1[1] = {1'b0,layer_1_1[3487:3480]} - {1'b0, layer_0_1[3487:3480]};
      top_1[2] = {1'b0,layer_1_1[3495:3488]} - {1'b0, layer_0_1[3495:3488]};
      top_2[0] = {1'b0,layer_1_2[3479:3472]} - {1'b0, layer_0_2[3479:3472]};
      top_2[1] = {1'b0,layer_1_2[3487:3480]} - {1'b0, layer_0_2[3487:3480]};
      top_2[2] = {1'b0,layer_1_2[3495:3488]} - {1'b0, layer_0_2[3495:3488]};
      mid_0[0] = {1'b0,layer_2_0[3479:3472]} - {1'b0, layer_1_0[3479:3472]};
      mid_0[1] = {1'b0,layer_2_0[3487:3480]} - {1'b0, layer_1_0[3487:3480]};
      mid_0[2] = {1'b0,layer_2_0[3495:3488]} - {1'b0, layer_1_0[3495:3488]};
      mid_1[0] = {1'b0,layer_2_1[3479:3472]} - {1'b0, layer_1_1[3479:3472]};
      mid_1[1] = {1'b0,layer_2_1[3487:3480]} - {1'b0, layer_1_1[3487:3480]};
      mid_1[2] = {1'b0,layer_2_1[3495:3488]} - {1'b0, layer_1_1[3495:3488]};
      mid_2[0] = {1'b0,layer_2_2[3479:3472]} - {1'b0, layer_1_2[3479:3472]};
      mid_2[1] = {1'b0,layer_2_2[3487:3480]} - {1'b0, layer_1_2[3487:3480]};
      mid_2[2] = {1'b0,layer_2_2[3495:3488]} - {1'b0, layer_1_2[3495:3488]};
      btm_0[0] = {1'b0,layer_3_0[3479:3472]} - {1'b0, layer_2_0[3479:3472]};
      btm_0[1] = {1'b0,layer_3_0[3487:3480]} - {1'b0, layer_2_0[3487:3480]};
      btm_0[2] = {1'b0,layer_3_0[3495:3488]} - {1'b0, layer_2_0[3495:3488]};
      btm_1[0] = {1'b0,layer_3_1[3479:3472]} - {1'b0, layer_2_1[3479:3472]};
      btm_1[1] = {1'b0,layer_3_1[3487:3480]} - {1'b0, layer_2_1[3487:3480]};
      btm_1[2] = {1'b0,layer_3_1[3495:3488]} - {1'b0, layer_2_1[3495:3488]};
      btm_2[0] = {1'b0,layer_3_2[3479:3472]} - {1'b0, layer_2_2[3479:3472]};
      btm_2[1] = {1'b0,layer_3_2[3487:3480]} - {1'b0, layer_2_2[3487:3480]};
      btm_2[2] = {1'b0,layer_3_2[3495:3488]} - {1'b0, layer_2_2[3495:3488]};
    end
    'd436: begin
      top_0[0] = {1'b0,layer_1_0[3487:3480]} - {1'b0, layer_0_0[3487:3480]};
      top_0[1] = {1'b0,layer_1_0[3495:3488]} - {1'b0, layer_0_0[3495:3488]};
      top_0[2] = {1'b0,layer_1_0[3503:3496]} - {1'b0, layer_0_0[3503:3496]};
      top_1[0] = {1'b0,layer_1_1[3487:3480]} - {1'b0, layer_0_1[3487:3480]};
      top_1[1] = {1'b0,layer_1_1[3495:3488]} - {1'b0, layer_0_1[3495:3488]};
      top_1[2] = {1'b0,layer_1_1[3503:3496]} - {1'b0, layer_0_1[3503:3496]};
      top_2[0] = {1'b0,layer_1_2[3487:3480]} - {1'b0, layer_0_2[3487:3480]};
      top_2[1] = {1'b0,layer_1_2[3495:3488]} - {1'b0, layer_0_2[3495:3488]};
      top_2[2] = {1'b0,layer_1_2[3503:3496]} - {1'b0, layer_0_2[3503:3496]};
      mid_0[0] = {1'b0,layer_2_0[3487:3480]} - {1'b0, layer_1_0[3487:3480]};
      mid_0[1] = {1'b0,layer_2_0[3495:3488]} - {1'b0, layer_1_0[3495:3488]};
      mid_0[2] = {1'b0,layer_2_0[3503:3496]} - {1'b0, layer_1_0[3503:3496]};
      mid_1[0] = {1'b0,layer_2_1[3487:3480]} - {1'b0, layer_1_1[3487:3480]};
      mid_1[1] = {1'b0,layer_2_1[3495:3488]} - {1'b0, layer_1_1[3495:3488]};
      mid_1[2] = {1'b0,layer_2_1[3503:3496]} - {1'b0, layer_1_1[3503:3496]};
      mid_2[0] = {1'b0,layer_2_2[3487:3480]} - {1'b0, layer_1_2[3487:3480]};
      mid_2[1] = {1'b0,layer_2_2[3495:3488]} - {1'b0, layer_1_2[3495:3488]};
      mid_2[2] = {1'b0,layer_2_2[3503:3496]} - {1'b0, layer_1_2[3503:3496]};
      btm_0[0] = {1'b0,layer_3_0[3487:3480]} - {1'b0, layer_2_0[3487:3480]};
      btm_0[1] = {1'b0,layer_3_0[3495:3488]} - {1'b0, layer_2_0[3495:3488]};
      btm_0[2] = {1'b0,layer_3_0[3503:3496]} - {1'b0, layer_2_0[3503:3496]};
      btm_1[0] = {1'b0,layer_3_1[3487:3480]} - {1'b0, layer_2_1[3487:3480]};
      btm_1[1] = {1'b0,layer_3_1[3495:3488]} - {1'b0, layer_2_1[3495:3488]};
      btm_1[2] = {1'b0,layer_3_1[3503:3496]} - {1'b0, layer_2_1[3503:3496]};
      btm_2[0] = {1'b0,layer_3_2[3487:3480]} - {1'b0, layer_2_2[3487:3480]};
      btm_2[1] = {1'b0,layer_3_2[3495:3488]} - {1'b0, layer_2_2[3495:3488]};
      btm_2[2] = {1'b0,layer_3_2[3503:3496]} - {1'b0, layer_2_2[3503:3496]};
    end
    'd437: begin
      top_0[0] = {1'b0,layer_1_0[3495:3488]} - {1'b0, layer_0_0[3495:3488]};
      top_0[1] = {1'b0,layer_1_0[3503:3496]} - {1'b0, layer_0_0[3503:3496]};
      top_0[2] = {1'b0,layer_1_0[3511:3504]} - {1'b0, layer_0_0[3511:3504]};
      top_1[0] = {1'b0,layer_1_1[3495:3488]} - {1'b0, layer_0_1[3495:3488]};
      top_1[1] = {1'b0,layer_1_1[3503:3496]} - {1'b0, layer_0_1[3503:3496]};
      top_1[2] = {1'b0,layer_1_1[3511:3504]} - {1'b0, layer_0_1[3511:3504]};
      top_2[0] = {1'b0,layer_1_2[3495:3488]} - {1'b0, layer_0_2[3495:3488]};
      top_2[1] = {1'b0,layer_1_2[3503:3496]} - {1'b0, layer_0_2[3503:3496]};
      top_2[2] = {1'b0,layer_1_2[3511:3504]} - {1'b0, layer_0_2[3511:3504]};
      mid_0[0] = {1'b0,layer_2_0[3495:3488]} - {1'b0, layer_1_0[3495:3488]};
      mid_0[1] = {1'b0,layer_2_0[3503:3496]} - {1'b0, layer_1_0[3503:3496]};
      mid_0[2] = {1'b0,layer_2_0[3511:3504]} - {1'b0, layer_1_0[3511:3504]};
      mid_1[0] = {1'b0,layer_2_1[3495:3488]} - {1'b0, layer_1_1[3495:3488]};
      mid_1[1] = {1'b0,layer_2_1[3503:3496]} - {1'b0, layer_1_1[3503:3496]};
      mid_1[2] = {1'b0,layer_2_1[3511:3504]} - {1'b0, layer_1_1[3511:3504]};
      mid_2[0] = {1'b0,layer_2_2[3495:3488]} - {1'b0, layer_1_2[3495:3488]};
      mid_2[1] = {1'b0,layer_2_2[3503:3496]} - {1'b0, layer_1_2[3503:3496]};
      mid_2[2] = {1'b0,layer_2_2[3511:3504]} - {1'b0, layer_1_2[3511:3504]};
      btm_0[0] = {1'b0,layer_3_0[3495:3488]} - {1'b0, layer_2_0[3495:3488]};
      btm_0[1] = {1'b0,layer_3_0[3503:3496]} - {1'b0, layer_2_0[3503:3496]};
      btm_0[2] = {1'b0,layer_3_0[3511:3504]} - {1'b0, layer_2_0[3511:3504]};
      btm_1[0] = {1'b0,layer_3_1[3495:3488]} - {1'b0, layer_2_1[3495:3488]};
      btm_1[1] = {1'b0,layer_3_1[3503:3496]} - {1'b0, layer_2_1[3503:3496]};
      btm_1[2] = {1'b0,layer_3_1[3511:3504]} - {1'b0, layer_2_1[3511:3504]};
      btm_2[0] = {1'b0,layer_3_2[3495:3488]} - {1'b0, layer_2_2[3495:3488]};
      btm_2[1] = {1'b0,layer_3_2[3503:3496]} - {1'b0, layer_2_2[3503:3496]};
      btm_2[2] = {1'b0,layer_3_2[3511:3504]} - {1'b0, layer_2_2[3511:3504]};
    end
    'd438: begin
      top_0[0] = {1'b0,layer_1_0[3503:3496]} - {1'b0, layer_0_0[3503:3496]};
      top_0[1] = {1'b0,layer_1_0[3511:3504]} - {1'b0, layer_0_0[3511:3504]};
      top_0[2] = {1'b0,layer_1_0[3519:3512]} - {1'b0, layer_0_0[3519:3512]};
      top_1[0] = {1'b0,layer_1_1[3503:3496]} - {1'b0, layer_0_1[3503:3496]};
      top_1[1] = {1'b0,layer_1_1[3511:3504]} - {1'b0, layer_0_1[3511:3504]};
      top_1[2] = {1'b0,layer_1_1[3519:3512]} - {1'b0, layer_0_1[3519:3512]};
      top_2[0] = {1'b0,layer_1_2[3503:3496]} - {1'b0, layer_0_2[3503:3496]};
      top_2[1] = {1'b0,layer_1_2[3511:3504]} - {1'b0, layer_0_2[3511:3504]};
      top_2[2] = {1'b0,layer_1_2[3519:3512]} - {1'b0, layer_0_2[3519:3512]};
      mid_0[0] = {1'b0,layer_2_0[3503:3496]} - {1'b0, layer_1_0[3503:3496]};
      mid_0[1] = {1'b0,layer_2_0[3511:3504]} - {1'b0, layer_1_0[3511:3504]};
      mid_0[2] = {1'b0,layer_2_0[3519:3512]} - {1'b0, layer_1_0[3519:3512]};
      mid_1[0] = {1'b0,layer_2_1[3503:3496]} - {1'b0, layer_1_1[3503:3496]};
      mid_1[1] = {1'b0,layer_2_1[3511:3504]} - {1'b0, layer_1_1[3511:3504]};
      mid_1[2] = {1'b0,layer_2_1[3519:3512]} - {1'b0, layer_1_1[3519:3512]};
      mid_2[0] = {1'b0,layer_2_2[3503:3496]} - {1'b0, layer_1_2[3503:3496]};
      mid_2[1] = {1'b0,layer_2_2[3511:3504]} - {1'b0, layer_1_2[3511:3504]};
      mid_2[2] = {1'b0,layer_2_2[3519:3512]} - {1'b0, layer_1_2[3519:3512]};
      btm_0[0] = {1'b0,layer_3_0[3503:3496]} - {1'b0, layer_2_0[3503:3496]};
      btm_0[1] = {1'b0,layer_3_0[3511:3504]} - {1'b0, layer_2_0[3511:3504]};
      btm_0[2] = {1'b0,layer_3_0[3519:3512]} - {1'b0, layer_2_0[3519:3512]};
      btm_1[0] = {1'b0,layer_3_1[3503:3496]} - {1'b0, layer_2_1[3503:3496]};
      btm_1[1] = {1'b0,layer_3_1[3511:3504]} - {1'b0, layer_2_1[3511:3504]};
      btm_1[2] = {1'b0,layer_3_1[3519:3512]} - {1'b0, layer_2_1[3519:3512]};
      btm_2[0] = {1'b0,layer_3_2[3503:3496]} - {1'b0, layer_2_2[3503:3496]};
      btm_2[1] = {1'b0,layer_3_2[3511:3504]} - {1'b0, layer_2_2[3511:3504]};
      btm_2[2] = {1'b0,layer_3_2[3519:3512]} - {1'b0, layer_2_2[3519:3512]};
    end
    'd439: begin
      top_0[0] = {1'b0,layer_1_0[3511:3504]} - {1'b0, layer_0_0[3511:3504]};
      top_0[1] = {1'b0,layer_1_0[3519:3512]} - {1'b0, layer_0_0[3519:3512]};
      top_0[2] = {1'b0,layer_1_0[3527:3520]} - {1'b0, layer_0_0[3527:3520]};
      top_1[0] = {1'b0,layer_1_1[3511:3504]} - {1'b0, layer_0_1[3511:3504]};
      top_1[1] = {1'b0,layer_1_1[3519:3512]} - {1'b0, layer_0_1[3519:3512]};
      top_1[2] = {1'b0,layer_1_1[3527:3520]} - {1'b0, layer_0_1[3527:3520]};
      top_2[0] = {1'b0,layer_1_2[3511:3504]} - {1'b0, layer_0_2[3511:3504]};
      top_2[1] = {1'b0,layer_1_2[3519:3512]} - {1'b0, layer_0_2[3519:3512]};
      top_2[2] = {1'b0,layer_1_2[3527:3520]} - {1'b0, layer_0_2[3527:3520]};
      mid_0[0] = {1'b0,layer_2_0[3511:3504]} - {1'b0, layer_1_0[3511:3504]};
      mid_0[1] = {1'b0,layer_2_0[3519:3512]} - {1'b0, layer_1_0[3519:3512]};
      mid_0[2] = {1'b0,layer_2_0[3527:3520]} - {1'b0, layer_1_0[3527:3520]};
      mid_1[0] = {1'b0,layer_2_1[3511:3504]} - {1'b0, layer_1_1[3511:3504]};
      mid_1[1] = {1'b0,layer_2_1[3519:3512]} - {1'b0, layer_1_1[3519:3512]};
      mid_1[2] = {1'b0,layer_2_1[3527:3520]} - {1'b0, layer_1_1[3527:3520]};
      mid_2[0] = {1'b0,layer_2_2[3511:3504]} - {1'b0, layer_1_2[3511:3504]};
      mid_2[1] = {1'b0,layer_2_2[3519:3512]} - {1'b0, layer_1_2[3519:3512]};
      mid_2[2] = {1'b0,layer_2_2[3527:3520]} - {1'b0, layer_1_2[3527:3520]};
      btm_0[0] = {1'b0,layer_3_0[3511:3504]} - {1'b0, layer_2_0[3511:3504]};
      btm_0[1] = {1'b0,layer_3_0[3519:3512]} - {1'b0, layer_2_0[3519:3512]};
      btm_0[2] = {1'b0,layer_3_0[3527:3520]} - {1'b0, layer_2_0[3527:3520]};
      btm_1[0] = {1'b0,layer_3_1[3511:3504]} - {1'b0, layer_2_1[3511:3504]};
      btm_1[1] = {1'b0,layer_3_1[3519:3512]} - {1'b0, layer_2_1[3519:3512]};
      btm_1[2] = {1'b0,layer_3_1[3527:3520]} - {1'b0, layer_2_1[3527:3520]};
      btm_2[0] = {1'b0,layer_3_2[3511:3504]} - {1'b0, layer_2_2[3511:3504]};
      btm_2[1] = {1'b0,layer_3_2[3519:3512]} - {1'b0, layer_2_2[3519:3512]};
      btm_2[2] = {1'b0,layer_3_2[3527:3520]} - {1'b0, layer_2_2[3527:3520]};
    end
    'd440: begin
      top_0[0] = {1'b0,layer_1_0[3519:3512]} - {1'b0, layer_0_0[3519:3512]};
      top_0[1] = {1'b0,layer_1_0[3527:3520]} - {1'b0, layer_0_0[3527:3520]};
      top_0[2] = {1'b0,layer_1_0[3535:3528]} - {1'b0, layer_0_0[3535:3528]};
      top_1[0] = {1'b0,layer_1_1[3519:3512]} - {1'b0, layer_0_1[3519:3512]};
      top_1[1] = {1'b0,layer_1_1[3527:3520]} - {1'b0, layer_0_1[3527:3520]};
      top_1[2] = {1'b0,layer_1_1[3535:3528]} - {1'b0, layer_0_1[3535:3528]};
      top_2[0] = {1'b0,layer_1_2[3519:3512]} - {1'b0, layer_0_2[3519:3512]};
      top_2[1] = {1'b0,layer_1_2[3527:3520]} - {1'b0, layer_0_2[3527:3520]};
      top_2[2] = {1'b0,layer_1_2[3535:3528]} - {1'b0, layer_0_2[3535:3528]};
      mid_0[0] = {1'b0,layer_2_0[3519:3512]} - {1'b0, layer_1_0[3519:3512]};
      mid_0[1] = {1'b0,layer_2_0[3527:3520]} - {1'b0, layer_1_0[3527:3520]};
      mid_0[2] = {1'b0,layer_2_0[3535:3528]} - {1'b0, layer_1_0[3535:3528]};
      mid_1[0] = {1'b0,layer_2_1[3519:3512]} - {1'b0, layer_1_1[3519:3512]};
      mid_1[1] = {1'b0,layer_2_1[3527:3520]} - {1'b0, layer_1_1[3527:3520]};
      mid_1[2] = {1'b0,layer_2_1[3535:3528]} - {1'b0, layer_1_1[3535:3528]};
      mid_2[0] = {1'b0,layer_2_2[3519:3512]} - {1'b0, layer_1_2[3519:3512]};
      mid_2[1] = {1'b0,layer_2_2[3527:3520]} - {1'b0, layer_1_2[3527:3520]};
      mid_2[2] = {1'b0,layer_2_2[3535:3528]} - {1'b0, layer_1_2[3535:3528]};
      btm_0[0] = {1'b0,layer_3_0[3519:3512]} - {1'b0, layer_2_0[3519:3512]};
      btm_0[1] = {1'b0,layer_3_0[3527:3520]} - {1'b0, layer_2_0[3527:3520]};
      btm_0[2] = {1'b0,layer_3_0[3535:3528]} - {1'b0, layer_2_0[3535:3528]};
      btm_1[0] = {1'b0,layer_3_1[3519:3512]} - {1'b0, layer_2_1[3519:3512]};
      btm_1[1] = {1'b0,layer_3_1[3527:3520]} - {1'b0, layer_2_1[3527:3520]};
      btm_1[2] = {1'b0,layer_3_1[3535:3528]} - {1'b0, layer_2_1[3535:3528]};
      btm_2[0] = {1'b0,layer_3_2[3519:3512]} - {1'b0, layer_2_2[3519:3512]};
      btm_2[1] = {1'b0,layer_3_2[3527:3520]} - {1'b0, layer_2_2[3527:3520]};
      btm_2[2] = {1'b0,layer_3_2[3535:3528]} - {1'b0, layer_2_2[3535:3528]};
    end
    'd441: begin
      top_0[0] = {1'b0,layer_1_0[3527:3520]} - {1'b0, layer_0_0[3527:3520]};
      top_0[1] = {1'b0,layer_1_0[3535:3528]} - {1'b0, layer_0_0[3535:3528]};
      top_0[2] = {1'b0,layer_1_0[3543:3536]} - {1'b0, layer_0_0[3543:3536]};
      top_1[0] = {1'b0,layer_1_1[3527:3520]} - {1'b0, layer_0_1[3527:3520]};
      top_1[1] = {1'b0,layer_1_1[3535:3528]} - {1'b0, layer_0_1[3535:3528]};
      top_1[2] = {1'b0,layer_1_1[3543:3536]} - {1'b0, layer_0_1[3543:3536]};
      top_2[0] = {1'b0,layer_1_2[3527:3520]} - {1'b0, layer_0_2[3527:3520]};
      top_2[1] = {1'b0,layer_1_2[3535:3528]} - {1'b0, layer_0_2[3535:3528]};
      top_2[2] = {1'b0,layer_1_2[3543:3536]} - {1'b0, layer_0_2[3543:3536]};
      mid_0[0] = {1'b0,layer_2_0[3527:3520]} - {1'b0, layer_1_0[3527:3520]};
      mid_0[1] = {1'b0,layer_2_0[3535:3528]} - {1'b0, layer_1_0[3535:3528]};
      mid_0[2] = {1'b0,layer_2_0[3543:3536]} - {1'b0, layer_1_0[3543:3536]};
      mid_1[0] = {1'b0,layer_2_1[3527:3520]} - {1'b0, layer_1_1[3527:3520]};
      mid_1[1] = {1'b0,layer_2_1[3535:3528]} - {1'b0, layer_1_1[3535:3528]};
      mid_1[2] = {1'b0,layer_2_1[3543:3536]} - {1'b0, layer_1_1[3543:3536]};
      mid_2[0] = {1'b0,layer_2_2[3527:3520]} - {1'b0, layer_1_2[3527:3520]};
      mid_2[1] = {1'b0,layer_2_2[3535:3528]} - {1'b0, layer_1_2[3535:3528]};
      mid_2[2] = {1'b0,layer_2_2[3543:3536]} - {1'b0, layer_1_2[3543:3536]};
      btm_0[0] = {1'b0,layer_3_0[3527:3520]} - {1'b0, layer_2_0[3527:3520]};
      btm_0[1] = {1'b0,layer_3_0[3535:3528]} - {1'b0, layer_2_0[3535:3528]};
      btm_0[2] = {1'b0,layer_3_0[3543:3536]} - {1'b0, layer_2_0[3543:3536]};
      btm_1[0] = {1'b0,layer_3_1[3527:3520]} - {1'b0, layer_2_1[3527:3520]};
      btm_1[1] = {1'b0,layer_3_1[3535:3528]} - {1'b0, layer_2_1[3535:3528]};
      btm_1[2] = {1'b0,layer_3_1[3543:3536]} - {1'b0, layer_2_1[3543:3536]};
      btm_2[0] = {1'b0,layer_3_2[3527:3520]} - {1'b0, layer_2_2[3527:3520]};
      btm_2[1] = {1'b0,layer_3_2[3535:3528]} - {1'b0, layer_2_2[3535:3528]};
      btm_2[2] = {1'b0,layer_3_2[3543:3536]} - {1'b0, layer_2_2[3543:3536]};
    end
    'd442: begin
      top_0[0] = {1'b0,layer_1_0[3535:3528]} - {1'b0, layer_0_0[3535:3528]};
      top_0[1] = {1'b0,layer_1_0[3543:3536]} - {1'b0, layer_0_0[3543:3536]};
      top_0[2] = {1'b0,layer_1_0[3551:3544]} - {1'b0, layer_0_0[3551:3544]};
      top_1[0] = {1'b0,layer_1_1[3535:3528]} - {1'b0, layer_0_1[3535:3528]};
      top_1[1] = {1'b0,layer_1_1[3543:3536]} - {1'b0, layer_0_1[3543:3536]};
      top_1[2] = {1'b0,layer_1_1[3551:3544]} - {1'b0, layer_0_1[3551:3544]};
      top_2[0] = {1'b0,layer_1_2[3535:3528]} - {1'b0, layer_0_2[3535:3528]};
      top_2[1] = {1'b0,layer_1_2[3543:3536]} - {1'b0, layer_0_2[3543:3536]};
      top_2[2] = {1'b0,layer_1_2[3551:3544]} - {1'b0, layer_0_2[3551:3544]};
      mid_0[0] = {1'b0,layer_2_0[3535:3528]} - {1'b0, layer_1_0[3535:3528]};
      mid_0[1] = {1'b0,layer_2_0[3543:3536]} - {1'b0, layer_1_0[3543:3536]};
      mid_0[2] = {1'b0,layer_2_0[3551:3544]} - {1'b0, layer_1_0[3551:3544]};
      mid_1[0] = {1'b0,layer_2_1[3535:3528]} - {1'b0, layer_1_1[3535:3528]};
      mid_1[1] = {1'b0,layer_2_1[3543:3536]} - {1'b0, layer_1_1[3543:3536]};
      mid_1[2] = {1'b0,layer_2_1[3551:3544]} - {1'b0, layer_1_1[3551:3544]};
      mid_2[0] = {1'b0,layer_2_2[3535:3528]} - {1'b0, layer_1_2[3535:3528]};
      mid_2[1] = {1'b0,layer_2_2[3543:3536]} - {1'b0, layer_1_2[3543:3536]};
      mid_2[2] = {1'b0,layer_2_2[3551:3544]} - {1'b0, layer_1_2[3551:3544]};
      btm_0[0] = {1'b0,layer_3_0[3535:3528]} - {1'b0, layer_2_0[3535:3528]};
      btm_0[1] = {1'b0,layer_3_0[3543:3536]} - {1'b0, layer_2_0[3543:3536]};
      btm_0[2] = {1'b0,layer_3_0[3551:3544]} - {1'b0, layer_2_0[3551:3544]};
      btm_1[0] = {1'b0,layer_3_1[3535:3528]} - {1'b0, layer_2_1[3535:3528]};
      btm_1[1] = {1'b0,layer_3_1[3543:3536]} - {1'b0, layer_2_1[3543:3536]};
      btm_1[2] = {1'b0,layer_3_1[3551:3544]} - {1'b0, layer_2_1[3551:3544]};
      btm_2[0] = {1'b0,layer_3_2[3535:3528]} - {1'b0, layer_2_2[3535:3528]};
      btm_2[1] = {1'b0,layer_3_2[3543:3536]} - {1'b0, layer_2_2[3543:3536]};
      btm_2[2] = {1'b0,layer_3_2[3551:3544]} - {1'b0, layer_2_2[3551:3544]};
    end
    'd443: begin
      top_0[0] = {1'b0,layer_1_0[3543:3536]} - {1'b0, layer_0_0[3543:3536]};
      top_0[1] = {1'b0,layer_1_0[3551:3544]} - {1'b0, layer_0_0[3551:3544]};
      top_0[2] = {1'b0,layer_1_0[3559:3552]} - {1'b0, layer_0_0[3559:3552]};
      top_1[0] = {1'b0,layer_1_1[3543:3536]} - {1'b0, layer_0_1[3543:3536]};
      top_1[1] = {1'b0,layer_1_1[3551:3544]} - {1'b0, layer_0_1[3551:3544]};
      top_1[2] = {1'b0,layer_1_1[3559:3552]} - {1'b0, layer_0_1[3559:3552]};
      top_2[0] = {1'b0,layer_1_2[3543:3536]} - {1'b0, layer_0_2[3543:3536]};
      top_2[1] = {1'b0,layer_1_2[3551:3544]} - {1'b0, layer_0_2[3551:3544]};
      top_2[2] = {1'b0,layer_1_2[3559:3552]} - {1'b0, layer_0_2[3559:3552]};
      mid_0[0] = {1'b0,layer_2_0[3543:3536]} - {1'b0, layer_1_0[3543:3536]};
      mid_0[1] = {1'b0,layer_2_0[3551:3544]} - {1'b0, layer_1_0[3551:3544]};
      mid_0[2] = {1'b0,layer_2_0[3559:3552]} - {1'b0, layer_1_0[3559:3552]};
      mid_1[0] = {1'b0,layer_2_1[3543:3536]} - {1'b0, layer_1_1[3543:3536]};
      mid_1[1] = {1'b0,layer_2_1[3551:3544]} - {1'b0, layer_1_1[3551:3544]};
      mid_1[2] = {1'b0,layer_2_1[3559:3552]} - {1'b0, layer_1_1[3559:3552]};
      mid_2[0] = {1'b0,layer_2_2[3543:3536]} - {1'b0, layer_1_2[3543:3536]};
      mid_2[1] = {1'b0,layer_2_2[3551:3544]} - {1'b0, layer_1_2[3551:3544]};
      mid_2[2] = {1'b0,layer_2_2[3559:3552]} - {1'b0, layer_1_2[3559:3552]};
      btm_0[0] = {1'b0,layer_3_0[3543:3536]} - {1'b0, layer_2_0[3543:3536]};
      btm_0[1] = {1'b0,layer_3_0[3551:3544]} - {1'b0, layer_2_0[3551:3544]};
      btm_0[2] = {1'b0,layer_3_0[3559:3552]} - {1'b0, layer_2_0[3559:3552]};
      btm_1[0] = {1'b0,layer_3_1[3543:3536]} - {1'b0, layer_2_1[3543:3536]};
      btm_1[1] = {1'b0,layer_3_1[3551:3544]} - {1'b0, layer_2_1[3551:3544]};
      btm_1[2] = {1'b0,layer_3_1[3559:3552]} - {1'b0, layer_2_1[3559:3552]};
      btm_2[0] = {1'b0,layer_3_2[3543:3536]} - {1'b0, layer_2_2[3543:3536]};
      btm_2[1] = {1'b0,layer_3_2[3551:3544]} - {1'b0, layer_2_2[3551:3544]};
      btm_2[2] = {1'b0,layer_3_2[3559:3552]} - {1'b0, layer_2_2[3559:3552]};
    end
    'd444: begin
      top_0[0] = {1'b0,layer_1_0[3551:3544]} - {1'b0, layer_0_0[3551:3544]};
      top_0[1] = {1'b0,layer_1_0[3559:3552]} - {1'b0, layer_0_0[3559:3552]};
      top_0[2] = {1'b0,layer_1_0[3567:3560]} - {1'b0, layer_0_0[3567:3560]};
      top_1[0] = {1'b0,layer_1_1[3551:3544]} - {1'b0, layer_0_1[3551:3544]};
      top_1[1] = {1'b0,layer_1_1[3559:3552]} - {1'b0, layer_0_1[3559:3552]};
      top_1[2] = {1'b0,layer_1_1[3567:3560]} - {1'b0, layer_0_1[3567:3560]};
      top_2[0] = {1'b0,layer_1_2[3551:3544]} - {1'b0, layer_0_2[3551:3544]};
      top_2[1] = {1'b0,layer_1_2[3559:3552]} - {1'b0, layer_0_2[3559:3552]};
      top_2[2] = {1'b0,layer_1_2[3567:3560]} - {1'b0, layer_0_2[3567:3560]};
      mid_0[0] = {1'b0,layer_2_0[3551:3544]} - {1'b0, layer_1_0[3551:3544]};
      mid_0[1] = {1'b0,layer_2_0[3559:3552]} - {1'b0, layer_1_0[3559:3552]};
      mid_0[2] = {1'b0,layer_2_0[3567:3560]} - {1'b0, layer_1_0[3567:3560]};
      mid_1[0] = {1'b0,layer_2_1[3551:3544]} - {1'b0, layer_1_1[3551:3544]};
      mid_1[1] = {1'b0,layer_2_1[3559:3552]} - {1'b0, layer_1_1[3559:3552]};
      mid_1[2] = {1'b0,layer_2_1[3567:3560]} - {1'b0, layer_1_1[3567:3560]};
      mid_2[0] = {1'b0,layer_2_2[3551:3544]} - {1'b0, layer_1_2[3551:3544]};
      mid_2[1] = {1'b0,layer_2_2[3559:3552]} - {1'b0, layer_1_2[3559:3552]};
      mid_2[2] = {1'b0,layer_2_2[3567:3560]} - {1'b0, layer_1_2[3567:3560]};
      btm_0[0] = {1'b0,layer_3_0[3551:3544]} - {1'b0, layer_2_0[3551:3544]};
      btm_0[1] = {1'b0,layer_3_0[3559:3552]} - {1'b0, layer_2_0[3559:3552]};
      btm_0[2] = {1'b0,layer_3_0[3567:3560]} - {1'b0, layer_2_0[3567:3560]};
      btm_1[0] = {1'b0,layer_3_1[3551:3544]} - {1'b0, layer_2_1[3551:3544]};
      btm_1[1] = {1'b0,layer_3_1[3559:3552]} - {1'b0, layer_2_1[3559:3552]};
      btm_1[2] = {1'b0,layer_3_1[3567:3560]} - {1'b0, layer_2_1[3567:3560]};
      btm_2[0] = {1'b0,layer_3_2[3551:3544]} - {1'b0, layer_2_2[3551:3544]};
      btm_2[1] = {1'b0,layer_3_2[3559:3552]} - {1'b0, layer_2_2[3559:3552]};
      btm_2[2] = {1'b0,layer_3_2[3567:3560]} - {1'b0, layer_2_2[3567:3560]};
    end
    'd445: begin
      top_0[0] = {1'b0,layer_1_0[3559:3552]} - {1'b0, layer_0_0[3559:3552]};
      top_0[1] = {1'b0,layer_1_0[3567:3560]} - {1'b0, layer_0_0[3567:3560]};
      top_0[2] = {1'b0,layer_1_0[3575:3568]} - {1'b0, layer_0_0[3575:3568]};
      top_1[0] = {1'b0,layer_1_1[3559:3552]} - {1'b0, layer_0_1[3559:3552]};
      top_1[1] = {1'b0,layer_1_1[3567:3560]} - {1'b0, layer_0_1[3567:3560]};
      top_1[2] = {1'b0,layer_1_1[3575:3568]} - {1'b0, layer_0_1[3575:3568]};
      top_2[0] = {1'b0,layer_1_2[3559:3552]} - {1'b0, layer_0_2[3559:3552]};
      top_2[1] = {1'b0,layer_1_2[3567:3560]} - {1'b0, layer_0_2[3567:3560]};
      top_2[2] = {1'b0,layer_1_2[3575:3568]} - {1'b0, layer_0_2[3575:3568]};
      mid_0[0] = {1'b0,layer_2_0[3559:3552]} - {1'b0, layer_1_0[3559:3552]};
      mid_0[1] = {1'b0,layer_2_0[3567:3560]} - {1'b0, layer_1_0[3567:3560]};
      mid_0[2] = {1'b0,layer_2_0[3575:3568]} - {1'b0, layer_1_0[3575:3568]};
      mid_1[0] = {1'b0,layer_2_1[3559:3552]} - {1'b0, layer_1_1[3559:3552]};
      mid_1[1] = {1'b0,layer_2_1[3567:3560]} - {1'b0, layer_1_1[3567:3560]};
      mid_1[2] = {1'b0,layer_2_1[3575:3568]} - {1'b0, layer_1_1[3575:3568]};
      mid_2[0] = {1'b0,layer_2_2[3559:3552]} - {1'b0, layer_1_2[3559:3552]};
      mid_2[1] = {1'b0,layer_2_2[3567:3560]} - {1'b0, layer_1_2[3567:3560]};
      mid_2[2] = {1'b0,layer_2_2[3575:3568]} - {1'b0, layer_1_2[3575:3568]};
      btm_0[0] = {1'b0,layer_3_0[3559:3552]} - {1'b0, layer_2_0[3559:3552]};
      btm_0[1] = {1'b0,layer_3_0[3567:3560]} - {1'b0, layer_2_0[3567:3560]};
      btm_0[2] = {1'b0,layer_3_0[3575:3568]} - {1'b0, layer_2_0[3575:3568]};
      btm_1[0] = {1'b0,layer_3_1[3559:3552]} - {1'b0, layer_2_1[3559:3552]};
      btm_1[1] = {1'b0,layer_3_1[3567:3560]} - {1'b0, layer_2_1[3567:3560]};
      btm_1[2] = {1'b0,layer_3_1[3575:3568]} - {1'b0, layer_2_1[3575:3568]};
      btm_2[0] = {1'b0,layer_3_2[3559:3552]} - {1'b0, layer_2_2[3559:3552]};
      btm_2[1] = {1'b0,layer_3_2[3567:3560]} - {1'b0, layer_2_2[3567:3560]};
      btm_2[2] = {1'b0,layer_3_2[3575:3568]} - {1'b0, layer_2_2[3575:3568]};
    end
    'd446: begin
      top_0[0] = {1'b0,layer_1_0[3567:3560]} - {1'b0, layer_0_0[3567:3560]};
      top_0[1] = {1'b0,layer_1_0[3575:3568]} - {1'b0, layer_0_0[3575:3568]};
      top_0[2] = {1'b0,layer_1_0[3583:3576]} - {1'b0, layer_0_0[3583:3576]};
      top_1[0] = {1'b0,layer_1_1[3567:3560]} - {1'b0, layer_0_1[3567:3560]};
      top_1[1] = {1'b0,layer_1_1[3575:3568]} - {1'b0, layer_0_1[3575:3568]};
      top_1[2] = {1'b0,layer_1_1[3583:3576]} - {1'b0, layer_0_1[3583:3576]};
      top_2[0] = {1'b0,layer_1_2[3567:3560]} - {1'b0, layer_0_2[3567:3560]};
      top_2[1] = {1'b0,layer_1_2[3575:3568]} - {1'b0, layer_0_2[3575:3568]};
      top_2[2] = {1'b0,layer_1_2[3583:3576]} - {1'b0, layer_0_2[3583:3576]};
      mid_0[0] = {1'b0,layer_2_0[3567:3560]} - {1'b0, layer_1_0[3567:3560]};
      mid_0[1] = {1'b0,layer_2_0[3575:3568]} - {1'b0, layer_1_0[3575:3568]};
      mid_0[2] = {1'b0,layer_2_0[3583:3576]} - {1'b0, layer_1_0[3583:3576]};
      mid_1[0] = {1'b0,layer_2_1[3567:3560]} - {1'b0, layer_1_1[3567:3560]};
      mid_1[1] = {1'b0,layer_2_1[3575:3568]} - {1'b0, layer_1_1[3575:3568]};
      mid_1[2] = {1'b0,layer_2_1[3583:3576]} - {1'b0, layer_1_1[3583:3576]};
      mid_2[0] = {1'b0,layer_2_2[3567:3560]} - {1'b0, layer_1_2[3567:3560]};
      mid_2[1] = {1'b0,layer_2_2[3575:3568]} - {1'b0, layer_1_2[3575:3568]};
      mid_2[2] = {1'b0,layer_2_2[3583:3576]} - {1'b0, layer_1_2[3583:3576]};
      btm_0[0] = {1'b0,layer_3_0[3567:3560]} - {1'b0, layer_2_0[3567:3560]};
      btm_0[1] = {1'b0,layer_3_0[3575:3568]} - {1'b0, layer_2_0[3575:3568]};
      btm_0[2] = {1'b0,layer_3_0[3583:3576]} - {1'b0, layer_2_0[3583:3576]};
      btm_1[0] = {1'b0,layer_3_1[3567:3560]} - {1'b0, layer_2_1[3567:3560]};
      btm_1[1] = {1'b0,layer_3_1[3575:3568]} - {1'b0, layer_2_1[3575:3568]};
      btm_1[2] = {1'b0,layer_3_1[3583:3576]} - {1'b0, layer_2_1[3583:3576]};
      btm_2[0] = {1'b0,layer_3_2[3567:3560]} - {1'b0, layer_2_2[3567:3560]};
      btm_2[1] = {1'b0,layer_3_2[3575:3568]} - {1'b0, layer_2_2[3575:3568]};
      btm_2[2] = {1'b0,layer_3_2[3583:3576]} - {1'b0, layer_2_2[3583:3576]};
    end
    'd447: begin
      top_0[0] = {1'b0,layer_1_0[3575:3568]} - {1'b0, layer_0_0[3575:3568]};
      top_0[1] = {1'b0,layer_1_0[3583:3576]} - {1'b0, layer_0_0[3583:3576]};
      top_0[2] = {1'b0,layer_1_0[3591:3584]} - {1'b0, layer_0_0[3591:3584]};
      top_1[0] = {1'b0,layer_1_1[3575:3568]} - {1'b0, layer_0_1[3575:3568]};
      top_1[1] = {1'b0,layer_1_1[3583:3576]} - {1'b0, layer_0_1[3583:3576]};
      top_1[2] = {1'b0,layer_1_1[3591:3584]} - {1'b0, layer_0_1[3591:3584]};
      top_2[0] = {1'b0,layer_1_2[3575:3568]} - {1'b0, layer_0_2[3575:3568]};
      top_2[1] = {1'b0,layer_1_2[3583:3576]} - {1'b0, layer_0_2[3583:3576]};
      top_2[2] = {1'b0,layer_1_2[3591:3584]} - {1'b0, layer_0_2[3591:3584]};
      mid_0[0] = {1'b0,layer_2_0[3575:3568]} - {1'b0, layer_1_0[3575:3568]};
      mid_0[1] = {1'b0,layer_2_0[3583:3576]} - {1'b0, layer_1_0[3583:3576]};
      mid_0[2] = {1'b0,layer_2_0[3591:3584]} - {1'b0, layer_1_0[3591:3584]};
      mid_1[0] = {1'b0,layer_2_1[3575:3568]} - {1'b0, layer_1_1[3575:3568]};
      mid_1[1] = {1'b0,layer_2_1[3583:3576]} - {1'b0, layer_1_1[3583:3576]};
      mid_1[2] = {1'b0,layer_2_1[3591:3584]} - {1'b0, layer_1_1[3591:3584]};
      mid_2[0] = {1'b0,layer_2_2[3575:3568]} - {1'b0, layer_1_2[3575:3568]};
      mid_2[1] = {1'b0,layer_2_2[3583:3576]} - {1'b0, layer_1_2[3583:3576]};
      mid_2[2] = {1'b0,layer_2_2[3591:3584]} - {1'b0, layer_1_2[3591:3584]};
      btm_0[0] = {1'b0,layer_3_0[3575:3568]} - {1'b0, layer_2_0[3575:3568]};
      btm_0[1] = {1'b0,layer_3_0[3583:3576]} - {1'b0, layer_2_0[3583:3576]};
      btm_0[2] = {1'b0,layer_3_0[3591:3584]} - {1'b0, layer_2_0[3591:3584]};
      btm_1[0] = {1'b0,layer_3_1[3575:3568]} - {1'b0, layer_2_1[3575:3568]};
      btm_1[1] = {1'b0,layer_3_1[3583:3576]} - {1'b0, layer_2_1[3583:3576]};
      btm_1[2] = {1'b0,layer_3_1[3591:3584]} - {1'b0, layer_2_1[3591:3584]};
      btm_2[0] = {1'b0,layer_3_2[3575:3568]} - {1'b0, layer_2_2[3575:3568]};
      btm_2[1] = {1'b0,layer_3_2[3583:3576]} - {1'b0, layer_2_2[3583:3576]};
      btm_2[2] = {1'b0,layer_3_2[3591:3584]} - {1'b0, layer_2_2[3591:3584]};
    end
    'd448: begin
      top_0[0] = {1'b0,layer_1_0[3583:3576]} - {1'b0, layer_0_0[3583:3576]};
      top_0[1] = {1'b0,layer_1_0[3591:3584]} - {1'b0, layer_0_0[3591:3584]};
      top_0[2] = {1'b0,layer_1_0[3599:3592]} - {1'b0, layer_0_0[3599:3592]};
      top_1[0] = {1'b0,layer_1_1[3583:3576]} - {1'b0, layer_0_1[3583:3576]};
      top_1[1] = {1'b0,layer_1_1[3591:3584]} - {1'b0, layer_0_1[3591:3584]};
      top_1[2] = {1'b0,layer_1_1[3599:3592]} - {1'b0, layer_0_1[3599:3592]};
      top_2[0] = {1'b0,layer_1_2[3583:3576]} - {1'b0, layer_0_2[3583:3576]};
      top_2[1] = {1'b0,layer_1_2[3591:3584]} - {1'b0, layer_0_2[3591:3584]};
      top_2[2] = {1'b0,layer_1_2[3599:3592]} - {1'b0, layer_0_2[3599:3592]};
      mid_0[0] = {1'b0,layer_2_0[3583:3576]} - {1'b0, layer_1_0[3583:3576]};
      mid_0[1] = {1'b0,layer_2_0[3591:3584]} - {1'b0, layer_1_0[3591:3584]};
      mid_0[2] = {1'b0,layer_2_0[3599:3592]} - {1'b0, layer_1_0[3599:3592]};
      mid_1[0] = {1'b0,layer_2_1[3583:3576]} - {1'b0, layer_1_1[3583:3576]};
      mid_1[1] = {1'b0,layer_2_1[3591:3584]} - {1'b0, layer_1_1[3591:3584]};
      mid_1[2] = {1'b0,layer_2_1[3599:3592]} - {1'b0, layer_1_1[3599:3592]};
      mid_2[0] = {1'b0,layer_2_2[3583:3576]} - {1'b0, layer_1_2[3583:3576]};
      mid_2[1] = {1'b0,layer_2_2[3591:3584]} - {1'b0, layer_1_2[3591:3584]};
      mid_2[2] = {1'b0,layer_2_2[3599:3592]} - {1'b0, layer_1_2[3599:3592]};
      btm_0[0] = {1'b0,layer_3_0[3583:3576]} - {1'b0, layer_2_0[3583:3576]};
      btm_0[1] = {1'b0,layer_3_0[3591:3584]} - {1'b0, layer_2_0[3591:3584]};
      btm_0[2] = {1'b0,layer_3_0[3599:3592]} - {1'b0, layer_2_0[3599:3592]};
      btm_1[0] = {1'b0,layer_3_1[3583:3576]} - {1'b0, layer_2_1[3583:3576]};
      btm_1[1] = {1'b0,layer_3_1[3591:3584]} - {1'b0, layer_2_1[3591:3584]};
      btm_1[2] = {1'b0,layer_3_1[3599:3592]} - {1'b0, layer_2_1[3599:3592]};
      btm_2[0] = {1'b0,layer_3_2[3583:3576]} - {1'b0, layer_2_2[3583:3576]};
      btm_2[1] = {1'b0,layer_3_2[3591:3584]} - {1'b0, layer_2_2[3591:3584]};
      btm_2[2] = {1'b0,layer_3_2[3599:3592]} - {1'b0, layer_2_2[3599:3592]};
    end
    'd449: begin
      top_0[0] = {1'b0,layer_1_0[3591:3584]} - {1'b0, layer_0_0[3591:3584]};
      top_0[1] = {1'b0,layer_1_0[3599:3592]} - {1'b0, layer_0_0[3599:3592]};
      top_0[2] = {1'b0,layer_1_0[3607:3600]} - {1'b0, layer_0_0[3607:3600]};
      top_1[0] = {1'b0,layer_1_1[3591:3584]} - {1'b0, layer_0_1[3591:3584]};
      top_1[1] = {1'b0,layer_1_1[3599:3592]} - {1'b0, layer_0_1[3599:3592]};
      top_1[2] = {1'b0,layer_1_1[3607:3600]} - {1'b0, layer_0_1[3607:3600]};
      top_2[0] = {1'b0,layer_1_2[3591:3584]} - {1'b0, layer_0_2[3591:3584]};
      top_2[1] = {1'b0,layer_1_2[3599:3592]} - {1'b0, layer_0_2[3599:3592]};
      top_2[2] = {1'b0,layer_1_2[3607:3600]} - {1'b0, layer_0_2[3607:3600]};
      mid_0[0] = {1'b0,layer_2_0[3591:3584]} - {1'b0, layer_1_0[3591:3584]};
      mid_0[1] = {1'b0,layer_2_0[3599:3592]} - {1'b0, layer_1_0[3599:3592]};
      mid_0[2] = {1'b0,layer_2_0[3607:3600]} - {1'b0, layer_1_0[3607:3600]};
      mid_1[0] = {1'b0,layer_2_1[3591:3584]} - {1'b0, layer_1_1[3591:3584]};
      mid_1[1] = {1'b0,layer_2_1[3599:3592]} - {1'b0, layer_1_1[3599:3592]};
      mid_1[2] = {1'b0,layer_2_1[3607:3600]} - {1'b0, layer_1_1[3607:3600]};
      mid_2[0] = {1'b0,layer_2_2[3591:3584]} - {1'b0, layer_1_2[3591:3584]};
      mid_2[1] = {1'b0,layer_2_2[3599:3592]} - {1'b0, layer_1_2[3599:3592]};
      mid_2[2] = {1'b0,layer_2_2[3607:3600]} - {1'b0, layer_1_2[3607:3600]};
      btm_0[0] = {1'b0,layer_3_0[3591:3584]} - {1'b0, layer_2_0[3591:3584]};
      btm_0[1] = {1'b0,layer_3_0[3599:3592]} - {1'b0, layer_2_0[3599:3592]};
      btm_0[2] = {1'b0,layer_3_0[3607:3600]} - {1'b0, layer_2_0[3607:3600]};
      btm_1[0] = {1'b0,layer_3_1[3591:3584]} - {1'b0, layer_2_1[3591:3584]};
      btm_1[1] = {1'b0,layer_3_1[3599:3592]} - {1'b0, layer_2_1[3599:3592]};
      btm_1[2] = {1'b0,layer_3_1[3607:3600]} - {1'b0, layer_2_1[3607:3600]};
      btm_2[0] = {1'b0,layer_3_2[3591:3584]} - {1'b0, layer_2_2[3591:3584]};
      btm_2[1] = {1'b0,layer_3_2[3599:3592]} - {1'b0, layer_2_2[3599:3592]};
      btm_2[2] = {1'b0,layer_3_2[3607:3600]} - {1'b0, layer_2_2[3607:3600]};
    end
    'd450: begin
      top_0[0] = {1'b0,layer_1_0[3599:3592]} - {1'b0, layer_0_0[3599:3592]};
      top_0[1] = {1'b0,layer_1_0[3607:3600]} - {1'b0, layer_0_0[3607:3600]};
      top_0[2] = {1'b0,layer_1_0[3615:3608]} - {1'b0, layer_0_0[3615:3608]};
      top_1[0] = {1'b0,layer_1_1[3599:3592]} - {1'b0, layer_0_1[3599:3592]};
      top_1[1] = {1'b0,layer_1_1[3607:3600]} - {1'b0, layer_0_1[3607:3600]};
      top_1[2] = {1'b0,layer_1_1[3615:3608]} - {1'b0, layer_0_1[3615:3608]};
      top_2[0] = {1'b0,layer_1_2[3599:3592]} - {1'b0, layer_0_2[3599:3592]};
      top_2[1] = {1'b0,layer_1_2[3607:3600]} - {1'b0, layer_0_2[3607:3600]};
      top_2[2] = {1'b0,layer_1_2[3615:3608]} - {1'b0, layer_0_2[3615:3608]};
      mid_0[0] = {1'b0,layer_2_0[3599:3592]} - {1'b0, layer_1_0[3599:3592]};
      mid_0[1] = {1'b0,layer_2_0[3607:3600]} - {1'b0, layer_1_0[3607:3600]};
      mid_0[2] = {1'b0,layer_2_0[3615:3608]} - {1'b0, layer_1_0[3615:3608]};
      mid_1[0] = {1'b0,layer_2_1[3599:3592]} - {1'b0, layer_1_1[3599:3592]};
      mid_1[1] = {1'b0,layer_2_1[3607:3600]} - {1'b0, layer_1_1[3607:3600]};
      mid_1[2] = {1'b0,layer_2_1[3615:3608]} - {1'b0, layer_1_1[3615:3608]};
      mid_2[0] = {1'b0,layer_2_2[3599:3592]} - {1'b0, layer_1_2[3599:3592]};
      mid_2[1] = {1'b0,layer_2_2[3607:3600]} - {1'b0, layer_1_2[3607:3600]};
      mid_2[2] = {1'b0,layer_2_2[3615:3608]} - {1'b0, layer_1_2[3615:3608]};
      btm_0[0] = {1'b0,layer_3_0[3599:3592]} - {1'b0, layer_2_0[3599:3592]};
      btm_0[1] = {1'b0,layer_3_0[3607:3600]} - {1'b0, layer_2_0[3607:3600]};
      btm_0[2] = {1'b0,layer_3_0[3615:3608]} - {1'b0, layer_2_0[3615:3608]};
      btm_1[0] = {1'b0,layer_3_1[3599:3592]} - {1'b0, layer_2_1[3599:3592]};
      btm_1[1] = {1'b0,layer_3_1[3607:3600]} - {1'b0, layer_2_1[3607:3600]};
      btm_1[2] = {1'b0,layer_3_1[3615:3608]} - {1'b0, layer_2_1[3615:3608]};
      btm_2[0] = {1'b0,layer_3_2[3599:3592]} - {1'b0, layer_2_2[3599:3592]};
      btm_2[1] = {1'b0,layer_3_2[3607:3600]} - {1'b0, layer_2_2[3607:3600]};
      btm_2[2] = {1'b0,layer_3_2[3615:3608]} - {1'b0, layer_2_2[3615:3608]};
    end
    'd451: begin
      top_0[0] = {1'b0,layer_1_0[3607:3600]} - {1'b0, layer_0_0[3607:3600]};
      top_0[1] = {1'b0,layer_1_0[3615:3608]} - {1'b0, layer_0_0[3615:3608]};
      top_0[2] = {1'b0,layer_1_0[3623:3616]} - {1'b0, layer_0_0[3623:3616]};
      top_1[0] = {1'b0,layer_1_1[3607:3600]} - {1'b0, layer_0_1[3607:3600]};
      top_1[1] = {1'b0,layer_1_1[3615:3608]} - {1'b0, layer_0_1[3615:3608]};
      top_1[2] = {1'b0,layer_1_1[3623:3616]} - {1'b0, layer_0_1[3623:3616]};
      top_2[0] = {1'b0,layer_1_2[3607:3600]} - {1'b0, layer_0_2[3607:3600]};
      top_2[1] = {1'b0,layer_1_2[3615:3608]} - {1'b0, layer_0_2[3615:3608]};
      top_2[2] = {1'b0,layer_1_2[3623:3616]} - {1'b0, layer_0_2[3623:3616]};
      mid_0[0] = {1'b0,layer_2_0[3607:3600]} - {1'b0, layer_1_0[3607:3600]};
      mid_0[1] = {1'b0,layer_2_0[3615:3608]} - {1'b0, layer_1_0[3615:3608]};
      mid_0[2] = {1'b0,layer_2_0[3623:3616]} - {1'b0, layer_1_0[3623:3616]};
      mid_1[0] = {1'b0,layer_2_1[3607:3600]} - {1'b0, layer_1_1[3607:3600]};
      mid_1[1] = {1'b0,layer_2_1[3615:3608]} - {1'b0, layer_1_1[3615:3608]};
      mid_1[2] = {1'b0,layer_2_1[3623:3616]} - {1'b0, layer_1_1[3623:3616]};
      mid_2[0] = {1'b0,layer_2_2[3607:3600]} - {1'b0, layer_1_2[3607:3600]};
      mid_2[1] = {1'b0,layer_2_2[3615:3608]} - {1'b0, layer_1_2[3615:3608]};
      mid_2[2] = {1'b0,layer_2_2[3623:3616]} - {1'b0, layer_1_2[3623:3616]};
      btm_0[0] = {1'b0,layer_3_0[3607:3600]} - {1'b0, layer_2_0[3607:3600]};
      btm_0[1] = {1'b0,layer_3_0[3615:3608]} - {1'b0, layer_2_0[3615:3608]};
      btm_0[2] = {1'b0,layer_3_0[3623:3616]} - {1'b0, layer_2_0[3623:3616]};
      btm_1[0] = {1'b0,layer_3_1[3607:3600]} - {1'b0, layer_2_1[3607:3600]};
      btm_1[1] = {1'b0,layer_3_1[3615:3608]} - {1'b0, layer_2_1[3615:3608]};
      btm_1[2] = {1'b0,layer_3_1[3623:3616]} - {1'b0, layer_2_1[3623:3616]};
      btm_2[0] = {1'b0,layer_3_2[3607:3600]} - {1'b0, layer_2_2[3607:3600]};
      btm_2[1] = {1'b0,layer_3_2[3615:3608]} - {1'b0, layer_2_2[3615:3608]};
      btm_2[2] = {1'b0,layer_3_2[3623:3616]} - {1'b0, layer_2_2[3623:3616]};
    end
    'd452: begin
      top_0[0] = {1'b0,layer_1_0[3615:3608]} - {1'b0, layer_0_0[3615:3608]};
      top_0[1] = {1'b0,layer_1_0[3623:3616]} - {1'b0, layer_0_0[3623:3616]};
      top_0[2] = {1'b0,layer_1_0[3631:3624]} - {1'b0, layer_0_0[3631:3624]};
      top_1[0] = {1'b0,layer_1_1[3615:3608]} - {1'b0, layer_0_1[3615:3608]};
      top_1[1] = {1'b0,layer_1_1[3623:3616]} - {1'b0, layer_0_1[3623:3616]};
      top_1[2] = {1'b0,layer_1_1[3631:3624]} - {1'b0, layer_0_1[3631:3624]};
      top_2[0] = {1'b0,layer_1_2[3615:3608]} - {1'b0, layer_0_2[3615:3608]};
      top_2[1] = {1'b0,layer_1_2[3623:3616]} - {1'b0, layer_0_2[3623:3616]};
      top_2[2] = {1'b0,layer_1_2[3631:3624]} - {1'b0, layer_0_2[3631:3624]};
      mid_0[0] = {1'b0,layer_2_0[3615:3608]} - {1'b0, layer_1_0[3615:3608]};
      mid_0[1] = {1'b0,layer_2_0[3623:3616]} - {1'b0, layer_1_0[3623:3616]};
      mid_0[2] = {1'b0,layer_2_0[3631:3624]} - {1'b0, layer_1_0[3631:3624]};
      mid_1[0] = {1'b0,layer_2_1[3615:3608]} - {1'b0, layer_1_1[3615:3608]};
      mid_1[1] = {1'b0,layer_2_1[3623:3616]} - {1'b0, layer_1_1[3623:3616]};
      mid_1[2] = {1'b0,layer_2_1[3631:3624]} - {1'b0, layer_1_1[3631:3624]};
      mid_2[0] = {1'b0,layer_2_2[3615:3608]} - {1'b0, layer_1_2[3615:3608]};
      mid_2[1] = {1'b0,layer_2_2[3623:3616]} - {1'b0, layer_1_2[3623:3616]};
      mid_2[2] = {1'b0,layer_2_2[3631:3624]} - {1'b0, layer_1_2[3631:3624]};
      btm_0[0] = {1'b0,layer_3_0[3615:3608]} - {1'b0, layer_2_0[3615:3608]};
      btm_0[1] = {1'b0,layer_3_0[3623:3616]} - {1'b0, layer_2_0[3623:3616]};
      btm_0[2] = {1'b0,layer_3_0[3631:3624]} - {1'b0, layer_2_0[3631:3624]};
      btm_1[0] = {1'b0,layer_3_1[3615:3608]} - {1'b0, layer_2_1[3615:3608]};
      btm_1[1] = {1'b0,layer_3_1[3623:3616]} - {1'b0, layer_2_1[3623:3616]};
      btm_1[2] = {1'b0,layer_3_1[3631:3624]} - {1'b0, layer_2_1[3631:3624]};
      btm_2[0] = {1'b0,layer_3_2[3615:3608]} - {1'b0, layer_2_2[3615:3608]};
      btm_2[1] = {1'b0,layer_3_2[3623:3616]} - {1'b0, layer_2_2[3623:3616]};
      btm_2[2] = {1'b0,layer_3_2[3631:3624]} - {1'b0, layer_2_2[3631:3624]};
    end
    'd453: begin
      top_0[0] = {1'b0,layer_1_0[3623:3616]} - {1'b0, layer_0_0[3623:3616]};
      top_0[1] = {1'b0,layer_1_0[3631:3624]} - {1'b0, layer_0_0[3631:3624]};
      top_0[2] = {1'b0,layer_1_0[3639:3632]} - {1'b0, layer_0_0[3639:3632]};
      top_1[0] = {1'b0,layer_1_1[3623:3616]} - {1'b0, layer_0_1[3623:3616]};
      top_1[1] = {1'b0,layer_1_1[3631:3624]} - {1'b0, layer_0_1[3631:3624]};
      top_1[2] = {1'b0,layer_1_1[3639:3632]} - {1'b0, layer_0_1[3639:3632]};
      top_2[0] = {1'b0,layer_1_2[3623:3616]} - {1'b0, layer_0_2[3623:3616]};
      top_2[1] = {1'b0,layer_1_2[3631:3624]} - {1'b0, layer_0_2[3631:3624]};
      top_2[2] = {1'b0,layer_1_2[3639:3632]} - {1'b0, layer_0_2[3639:3632]};
      mid_0[0] = {1'b0,layer_2_0[3623:3616]} - {1'b0, layer_1_0[3623:3616]};
      mid_0[1] = {1'b0,layer_2_0[3631:3624]} - {1'b0, layer_1_0[3631:3624]};
      mid_0[2] = {1'b0,layer_2_0[3639:3632]} - {1'b0, layer_1_0[3639:3632]};
      mid_1[0] = {1'b0,layer_2_1[3623:3616]} - {1'b0, layer_1_1[3623:3616]};
      mid_1[1] = {1'b0,layer_2_1[3631:3624]} - {1'b0, layer_1_1[3631:3624]};
      mid_1[2] = {1'b0,layer_2_1[3639:3632]} - {1'b0, layer_1_1[3639:3632]};
      mid_2[0] = {1'b0,layer_2_2[3623:3616]} - {1'b0, layer_1_2[3623:3616]};
      mid_2[1] = {1'b0,layer_2_2[3631:3624]} - {1'b0, layer_1_2[3631:3624]};
      mid_2[2] = {1'b0,layer_2_2[3639:3632]} - {1'b0, layer_1_2[3639:3632]};
      btm_0[0] = {1'b0,layer_3_0[3623:3616]} - {1'b0, layer_2_0[3623:3616]};
      btm_0[1] = {1'b0,layer_3_0[3631:3624]} - {1'b0, layer_2_0[3631:3624]};
      btm_0[2] = {1'b0,layer_3_0[3639:3632]} - {1'b0, layer_2_0[3639:3632]};
      btm_1[0] = {1'b0,layer_3_1[3623:3616]} - {1'b0, layer_2_1[3623:3616]};
      btm_1[1] = {1'b0,layer_3_1[3631:3624]} - {1'b0, layer_2_1[3631:3624]};
      btm_1[2] = {1'b0,layer_3_1[3639:3632]} - {1'b0, layer_2_1[3639:3632]};
      btm_2[0] = {1'b0,layer_3_2[3623:3616]} - {1'b0, layer_2_2[3623:3616]};
      btm_2[1] = {1'b0,layer_3_2[3631:3624]} - {1'b0, layer_2_2[3631:3624]};
      btm_2[2] = {1'b0,layer_3_2[3639:3632]} - {1'b0, layer_2_2[3639:3632]};
    end
    'd454: begin
      top_0[0] = {1'b0,layer_1_0[3631:3624]} - {1'b0, layer_0_0[3631:3624]};
      top_0[1] = {1'b0,layer_1_0[3639:3632]} - {1'b0, layer_0_0[3639:3632]};
      top_0[2] = {1'b0,layer_1_0[3647:3640]} - {1'b0, layer_0_0[3647:3640]};
      top_1[0] = {1'b0,layer_1_1[3631:3624]} - {1'b0, layer_0_1[3631:3624]};
      top_1[1] = {1'b0,layer_1_1[3639:3632]} - {1'b0, layer_0_1[3639:3632]};
      top_1[2] = {1'b0,layer_1_1[3647:3640]} - {1'b0, layer_0_1[3647:3640]};
      top_2[0] = {1'b0,layer_1_2[3631:3624]} - {1'b0, layer_0_2[3631:3624]};
      top_2[1] = {1'b0,layer_1_2[3639:3632]} - {1'b0, layer_0_2[3639:3632]};
      top_2[2] = {1'b0,layer_1_2[3647:3640]} - {1'b0, layer_0_2[3647:3640]};
      mid_0[0] = {1'b0,layer_2_0[3631:3624]} - {1'b0, layer_1_0[3631:3624]};
      mid_0[1] = {1'b0,layer_2_0[3639:3632]} - {1'b0, layer_1_0[3639:3632]};
      mid_0[2] = {1'b0,layer_2_0[3647:3640]} - {1'b0, layer_1_0[3647:3640]};
      mid_1[0] = {1'b0,layer_2_1[3631:3624]} - {1'b0, layer_1_1[3631:3624]};
      mid_1[1] = {1'b0,layer_2_1[3639:3632]} - {1'b0, layer_1_1[3639:3632]};
      mid_1[2] = {1'b0,layer_2_1[3647:3640]} - {1'b0, layer_1_1[3647:3640]};
      mid_2[0] = {1'b0,layer_2_2[3631:3624]} - {1'b0, layer_1_2[3631:3624]};
      mid_2[1] = {1'b0,layer_2_2[3639:3632]} - {1'b0, layer_1_2[3639:3632]};
      mid_2[2] = {1'b0,layer_2_2[3647:3640]} - {1'b0, layer_1_2[3647:3640]};
      btm_0[0] = {1'b0,layer_3_0[3631:3624]} - {1'b0, layer_2_0[3631:3624]};
      btm_0[1] = {1'b0,layer_3_0[3639:3632]} - {1'b0, layer_2_0[3639:3632]};
      btm_0[2] = {1'b0,layer_3_0[3647:3640]} - {1'b0, layer_2_0[3647:3640]};
      btm_1[0] = {1'b0,layer_3_1[3631:3624]} - {1'b0, layer_2_1[3631:3624]};
      btm_1[1] = {1'b0,layer_3_1[3639:3632]} - {1'b0, layer_2_1[3639:3632]};
      btm_1[2] = {1'b0,layer_3_1[3647:3640]} - {1'b0, layer_2_1[3647:3640]};
      btm_2[0] = {1'b0,layer_3_2[3631:3624]} - {1'b0, layer_2_2[3631:3624]};
      btm_2[1] = {1'b0,layer_3_2[3639:3632]} - {1'b0, layer_2_2[3639:3632]};
      btm_2[2] = {1'b0,layer_3_2[3647:3640]} - {1'b0, layer_2_2[3647:3640]};
    end
    'd455: begin
      top_0[0] = {1'b0,layer_1_0[3639:3632]} - {1'b0, layer_0_0[3639:3632]};
      top_0[1] = {1'b0,layer_1_0[3647:3640]} - {1'b0, layer_0_0[3647:3640]};
      top_0[2] = {1'b0,layer_1_0[3655:3648]} - {1'b0, layer_0_0[3655:3648]};
      top_1[0] = {1'b0,layer_1_1[3639:3632]} - {1'b0, layer_0_1[3639:3632]};
      top_1[1] = {1'b0,layer_1_1[3647:3640]} - {1'b0, layer_0_1[3647:3640]};
      top_1[2] = {1'b0,layer_1_1[3655:3648]} - {1'b0, layer_0_1[3655:3648]};
      top_2[0] = {1'b0,layer_1_2[3639:3632]} - {1'b0, layer_0_2[3639:3632]};
      top_2[1] = {1'b0,layer_1_2[3647:3640]} - {1'b0, layer_0_2[3647:3640]};
      top_2[2] = {1'b0,layer_1_2[3655:3648]} - {1'b0, layer_0_2[3655:3648]};
      mid_0[0] = {1'b0,layer_2_0[3639:3632]} - {1'b0, layer_1_0[3639:3632]};
      mid_0[1] = {1'b0,layer_2_0[3647:3640]} - {1'b0, layer_1_0[3647:3640]};
      mid_0[2] = {1'b0,layer_2_0[3655:3648]} - {1'b0, layer_1_0[3655:3648]};
      mid_1[0] = {1'b0,layer_2_1[3639:3632]} - {1'b0, layer_1_1[3639:3632]};
      mid_1[1] = {1'b0,layer_2_1[3647:3640]} - {1'b0, layer_1_1[3647:3640]};
      mid_1[2] = {1'b0,layer_2_1[3655:3648]} - {1'b0, layer_1_1[3655:3648]};
      mid_2[0] = {1'b0,layer_2_2[3639:3632]} - {1'b0, layer_1_2[3639:3632]};
      mid_2[1] = {1'b0,layer_2_2[3647:3640]} - {1'b0, layer_1_2[3647:3640]};
      mid_2[2] = {1'b0,layer_2_2[3655:3648]} - {1'b0, layer_1_2[3655:3648]};
      btm_0[0] = {1'b0,layer_3_0[3639:3632]} - {1'b0, layer_2_0[3639:3632]};
      btm_0[1] = {1'b0,layer_3_0[3647:3640]} - {1'b0, layer_2_0[3647:3640]};
      btm_0[2] = {1'b0,layer_3_0[3655:3648]} - {1'b0, layer_2_0[3655:3648]};
      btm_1[0] = {1'b0,layer_3_1[3639:3632]} - {1'b0, layer_2_1[3639:3632]};
      btm_1[1] = {1'b0,layer_3_1[3647:3640]} - {1'b0, layer_2_1[3647:3640]};
      btm_1[2] = {1'b0,layer_3_1[3655:3648]} - {1'b0, layer_2_1[3655:3648]};
      btm_2[0] = {1'b0,layer_3_2[3639:3632]} - {1'b0, layer_2_2[3639:3632]};
      btm_2[1] = {1'b0,layer_3_2[3647:3640]} - {1'b0, layer_2_2[3647:3640]};
      btm_2[2] = {1'b0,layer_3_2[3655:3648]} - {1'b0, layer_2_2[3655:3648]};
    end
    'd456: begin
      top_0[0] = {1'b0,layer_1_0[3647:3640]} - {1'b0, layer_0_0[3647:3640]};
      top_0[1] = {1'b0,layer_1_0[3655:3648]} - {1'b0, layer_0_0[3655:3648]};
      top_0[2] = {1'b0,layer_1_0[3663:3656]} - {1'b0, layer_0_0[3663:3656]};
      top_1[0] = {1'b0,layer_1_1[3647:3640]} - {1'b0, layer_0_1[3647:3640]};
      top_1[1] = {1'b0,layer_1_1[3655:3648]} - {1'b0, layer_0_1[3655:3648]};
      top_1[2] = {1'b0,layer_1_1[3663:3656]} - {1'b0, layer_0_1[3663:3656]};
      top_2[0] = {1'b0,layer_1_2[3647:3640]} - {1'b0, layer_0_2[3647:3640]};
      top_2[1] = {1'b0,layer_1_2[3655:3648]} - {1'b0, layer_0_2[3655:3648]};
      top_2[2] = {1'b0,layer_1_2[3663:3656]} - {1'b0, layer_0_2[3663:3656]};
      mid_0[0] = {1'b0,layer_2_0[3647:3640]} - {1'b0, layer_1_0[3647:3640]};
      mid_0[1] = {1'b0,layer_2_0[3655:3648]} - {1'b0, layer_1_0[3655:3648]};
      mid_0[2] = {1'b0,layer_2_0[3663:3656]} - {1'b0, layer_1_0[3663:3656]};
      mid_1[0] = {1'b0,layer_2_1[3647:3640]} - {1'b0, layer_1_1[3647:3640]};
      mid_1[1] = {1'b0,layer_2_1[3655:3648]} - {1'b0, layer_1_1[3655:3648]};
      mid_1[2] = {1'b0,layer_2_1[3663:3656]} - {1'b0, layer_1_1[3663:3656]};
      mid_2[0] = {1'b0,layer_2_2[3647:3640]} - {1'b0, layer_1_2[3647:3640]};
      mid_2[1] = {1'b0,layer_2_2[3655:3648]} - {1'b0, layer_1_2[3655:3648]};
      mid_2[2] = {1'b0,layer_2_2[3663:3656]} - {1'b0, layer_1_2[3663:3656]};
      btm_0[0] = {1'b0,layer_3_0[3647:3640]} - {1'b0, layer_2_0[3647:3640]};
      btm_0[1] = {1'b0,layer_3_0[3655:3648]} - {1'b0, layer_2_0[3655:3648]};
      btm_0[2] = {1'b0,layer_3_0[3663:3656]} - {1'b0, layer_2_0[3663:3656]};
      btm_1[0] = {1'b0,layer_3_1[3647:3640]} - {1'b0, layer_2_1[3647:3640]};
      btm_1[1] = {1'b0,layer_3_1[3655:3648]} - {1'b0, layer_2_1[3655:3648]};
      btm_1[2] = {1'b0,layer_3_1[3663:3656]} - {1'b0, layer_2_1[3663:3656]};
      btm_2[0] = {1'b0,layer_3_2[3647:3640]} - {1'b0, layer_2_2[3647:3640]};
      btm_2[1] = {1'b0,layer_3_2[3655:3648]} - {1'b0, layer_2_2[3655:3648]};
      btm_2[2] = {1'b0,layer_3_2[3663:3656]} - {1'b0, layer_2_2[3663:3656]};
    end
    'd457: begin
      top_0[0] = {1'b0,layer_1_0[3655:3648]} - {1'b0, layer_0_0[3655:3648]};
      top_0[1] = {1'b0,layer_1_0[3663:3656]} - {1'b0, layer_0_0[3663:3656]};
      top_0[2] = {1'b0,layer_1_0[3671:3664]} - {1'b0, layer_0_0[3671:3664]};
      top_1[0] = {1'b0,layer_1_1[3655:3648]} - {1'b0, layer_0_1[3655:3648]};
      top_1[1] = {1'b0,layer_1_1[3663:3656]} - {1'b0, layer_0_1[3663:3656]};
      top_1[2] = {1'b0,layer_1_1[3671:3664]} - {1'b0, layer_0_1[3671:3664]};
      top_2[0] = {1'b0,layer_1_2[3655:3648]} - {1'b0, layer_0_2[3655:3648]};
      top_2[1] = {1'b0,layer_1_2[3663:3656]} - {1'b0, layer_0_2[3663:3656]};
      top_2[2] = {1'b0,layer_1_2[3671:3664]} - {1'b0, layer_0_2[3671:3664]};
      mid_0[0] = {1'b0,layer_2_0[3655:3648]} - {1'b0, layer_1_0[3655:3648]};
      mid_0[1] = {1'b0,layer_2_0[3663:3656]} - {1'b0, layer_1_0[3663:3656]};
      mid_0[2] = {1'b0,layer_2_0[3671:3664]} - {1'b0, layer_1_0[3671:3664]};
      mid_1[0] = {1'b0,layer_2_1[3655:3648]} - {1'b0, layer_1_1[3655:3648]};
      mid_1[1] = {1'b0,layer_2_1[3663:3656]} - {1'b0, layer_1_1[3663:3656]};
      mid_1[2] = {1'b0,layer_2_1[3671:3664]} - {1'b0, layer_1_1[3671:3664]};
      mid_2[0] = {1'b0,layer_2_2[3655:3648]} - {1'b0, layer_1_2[3655:3648]};
      mid_2[1] = {1'b0,layer_2_2[3663:3656]} - {1'b0, layer_1_2[3663:3656]};
      mid_2[2] = {1'b0,layer_2_2[3671:3664]} - {1'b0, layer_1_2[3671:3664]};
      btm_0[0] = {1'b0,layer_3_0[3655:3648]} - {1'b0, layer_2_0[3655:3648]};
      btm_0[1] = {1'b0,layer_3_0[3663:3656]} - {1'b0, layer_2_0[3663:3656]};
      btm_0[2] = {1'b0,layer_3_0[3671:3664]} - {1'b0, layer_2_0[3671:3664]};
      btm_1[0] = {1'b0,layer_3_1[3655:3648]} - {1'b0, layer_2_1[3655:3648]};
      btm_1[1] = {1'b0,layer_3_1[3663:3656]} - {1'b0, layer_2_1[3663:3656]};
      btm_1[2] = {1'b0,layer_3_1[3671:3664]} - {1'b0, layer_2_1[3671:3664]};
      btm_2[0] = {1'b0,layer_3_2[3655:3648]} - {1'b0, layer_2_2[3655:3648]};
      btm_2[1] = {1'b0,layer_3_2[3663:3656]} - {1'b0, layer_2_2[3663:3656]};
      btm_2[2] = {1'b0,layer_3_2[3671:3664]} - {1'b0, layer_2_2[3671:3664]};
    end
    'd458: begin
      top_0[0] = {1'b0,layer_1_0[3663:3656]} - {1'b0, layer_0_0[3663:3656]};
      top_0[1] = {1'b0,layer_1_0[3671:3664]} - {1'b0, layer_0_0[3671:3664]};
      top_0[2] = {1'b0,layer_1_0[3679:3672]} - {1'b0, layer_0_0[3679:3672]};
      top_1[0] = {1'b0,layer_1_1[3663:3656]} - {1'b0, layer_0_1[3663:3656]};
      top_1[1] = {1'b0,layer_1_1[3671:3664]} - {1'b0, layer_0_1[3671:3664]};
      top_1[2] = {1'b0,layer_1_1[3679:3672]} - {1'b0, layer_0_1[3679:3672]};
      top_2[0] = {1'b0,layer_1_2[3663:3656]} - {1'b0, layer_0_2[3663:3656]};
      top_2[1] = {1'b0,layer_1_2[3671:3664]} - {1'b0, layer_0_2[3671:3664]};
      top_2[2] = {1'b0,layer_1_2[3679:3672]} - {1'b0, layer_0_2[3679:3672]};
      mid_0[0] = {1'b0,layer_2_0[3663:3656]} - {1'b0, layer_1_0[3663:3656]};
      mid_0[1] = {1'b0,layer_2_0[3671:3664]} - {1'b0, layer_1_0[3671:3664]};
      mid_0[2] = {1'b0,layer_2_0[3679:3672]} - {1'b0, layer_1_0[3679:3672]};
      mid_1[0] = {1'b0,layer_2_1[3663:3656]} - {1'b0, layer_1_1[3663:3656]};
      mid_1[1] = {1'b0,layer_2_1[3671:3664]} - {1'b0, layer_1_1[3671:3664]};
      mid_1[2] = {1'b0,layer_2_1[3679:3672]} - {1'b0, layer_1_1[3679:3672]};
      mid_2[0] = {1'b0,layer_2_2[3663:3656]} - {1'b0, layer_1_2[3663:3656]};
      mid_2[1] = {1'b0,layer_2_2[3671:3664]} - {1'b0, layer_1_2[3671:3664]};
      mid_2[2] = {1'b0,layer_2_2[3679:3672]} - {1'b0, layer_1_2[3679:3672]};
      btm_0[0] = {1'b0,layer_3_0[3663:3656]} - {1'b0, layer_2_0[3663:3656]};
      btm_0[1] = {1'b0,layer_3_0[3671:3664]} - {1'b0, layer_2_0[3671:3664]};
      btm_0[2] = {1'b0,layer_3_0[3679:3672]} - {1'b0, layer_2_0[3679:3672]};
      btm_1[0] = {1'b0,layer_3_1[3663:3656]} - {1'b0, layer_2_1[3663:3656]};
      btm_1[1] = {1'b0,layer_3_1[3671:3664]} - {1'b0, layer_2_1[3671:3664]};
      btm_1[2] = {1'b0,layer_3_1[3679:3672]} - {1'b0, layer_2_1[3679:3672]};
      btm_2[0] = {1'b0,layer_3_2[3663:3656]} - {1'b0, layer_2_2[3663:3656]};
      btm_2[1] = {1'b0,layer_3_2[3671:3664]} - {1'b0, layer_2_2[3671:3664]};
      btm_2[2] = {1'b0,layer_3_2[3679:3672]} - {1'b0, layer_2_2[3679:3672]};
    end
    'd459: begin
      top_0[0] = {1'b0,layer_1_0[3671:3664]} - {1'b0, layer_0_0[3671:3664]};
      top_0[1] = {1'b0,layer_1_0[3679:3672]} - {1'b0, layer_0_0[3679:3672]};
      top_0[2] = {1'b0,layer_1_0[3687:3680]} - {1'b0, layer_0_0[3687:3680]};
      top_1[0] = {1'b0,layer_1_1[3671:3664]} - {1'b0, layer_0_1[3671:3664]};
      top_1[1] = {1'b0,layer_1_1[3679:3672]} - {1'b0, layer_0_1[3679:3672]};
      top_1[2] = {1'b0,layer_1_1[3687:3680]} - {1'b0, layer_0_1[3687:3680]};
      top_2[0] = {1'b0,layer_1_2[3671:3664]} - {1'b0, layer_0_2[3671:3664]};
      top_2[1] = {1'b0,layer_1_2[3679:3672]} - {1'b0, layer_0_2[3679:3672]};
      top_2[2] = {1'b0,layer_1_2[3687:3680]} - {1'b0, layer_0_2[3687:3680]};
      mid_0[0] = {1'b0,layer_2_0[3671:3664]} - {1'b0, layer_1_0[3671:3664]};
      mid_0[1] = {1'b0,layer_2_0[3679:3672]} - {1'b0, layer_1_0[3679:3672]};
      mid_0[2] = {1'b0,layer_2_0[3687:3680]} - {1'b0, layer_1_0[3687:3680]};
      mid_1[0] = {1'b0,layer_2_1[3671:3664]} - {1'b0, layer_1_1[3671:3664]};
      mid_1[1] = {1'b0,layer_2_1[3679:3672]} - {1'b0, layer_1_1[3679:3672]};
      mid_1[2] = {1'b0,layer_2_1[3687:3680]} - {1'b0, layer_1_1[3687:3680]};
      mid_2[0] = {1'b0,layer_2_2[3671:3664]} - {1'b0, layer_1_2[3671:3664]};
      mid_2[1] = {1'b0,layer_2_2[3679:3672]} - {1'b0, layer_1_2[3679:3672]};
      mid_2[2] = {1'b0,layer_2_2[3687:3680]} - {1'b0, layer_1_2[3687:3680]};
      btm_0[0] = {1'b0,layer_3_0[3671:3664]} - {1'b0, layer_2_0[3671:3664]};
      btm_0[1] = {1'b0,layer_3_0[3679:3672]} - {1'b0, layer_2_0[3679:3672]};
      btm_0[2] = {1'b0,layer_3_0[3687:3680]} - {1'b0, layer_2_0[3687:3680]};
      btm_1[0] = {1'b0,layer_3_1[3671:3664]} - {1'b0, layer_2_1[3671:3664]};
      btm_1[1] = {1'b0,layer_3_1[3679:3672]} - {1'b0, layer_2_1[3679:3672]};
      btm_1[2] = {1'b0,layer_3_1[3687:3680]} - {1'b0, layer_2_1[3687:3680]};
      btm_2[0] = {1'b0,layer_3_2[3671:3664]} - {1'b0, layer_2_2[3671:3664]};
      btm_2[1] = {1'b0,layer_3_2[3679:3672]} - {1'b0, layer_2_2[3679:3672]};
      btm_2[2] = {1'b0,layer_3_2[3687:3680]} - {1'b0, layer_2_2[3687:3680]};
    end
    'd460: begin
      top_0[0] = {1'b0,layer_1_0[3679:3672]} - {1'b0, layer_0_0[3679:3672]};
      top_0[1] = {1'b0,layer_1_0[3687:3680]} - {1'b0, layer_0_0[3687:3680]};
      top_0[2] = {1'b0,layer_1_0[3695:3688]} - {1'b0, layer_0_0[3695:3688]};
      top_1[0] = {1'b0,layer_1_1[3679:3672]} - {1'b0, layer_0_1[3679:3672]};
      top_1[1] = {1'b0,layer_1_1[3687:3680]} - {1'b0, layer_0_1[3687:3680]};
      top_1[2] = {1'b0,layer_1_1[3695:3688]} - {1'b0, layer_0_1[3695:3688]};
      top_2[0] = {1'b0,layer_1_2[3679:3672]} - {1'b0, layer_0_2[3679:3672]};
      top_2[1] = {1'b0,layer_1_2[3687:3680]} - {1'b0, layer_0_2[3687:3680]};
      top_2[2] = {1'b0,layer_1_2[3695:3688]} - {1'b0, layer_0_2[3695:3688]};
      mid_0[0] = {1'b0,layer_2_0[3679:3672]} - {1'b0, layer_1_0[3679:3672]};
      mid_0[1] = {1'b0,layer_2_0[3687:3680]} - {1'b0, layer_1_0[3687:3680]};
      mid_0[2] = {1'b0,layer_2_0[3695:3688]} - {1'b0, layer_1_0[3695:3688]};
      mid_1[0] = {1'b0,layer_2_1[3679:3672]} - {1'b0, layer_1_1[3679:3672]};
      mid_1[1] = {1'b0,layer_2_1[3687:3680]} - {1'b0, layer_1_1[3687:3680]};
      mid_1[2] = {1'b0,layer_2_1[3695:3688]} - {1'b0, layer_1_1[3695:3688]};
      mid_2[0] = {1'b0,layer_2_2[3679:3672]} - {1'b0, layer_1_2[3679:3672]};
      mid_2[1] = {1'b0,layer_2_2[3687:3680]} - {1'b0, layer_1_2[3687:3680]};
      mid_2[2] = {1'b0,layer_2_2[3695:3688]} - {1'b0, layer_1_2[3695:3688]};
      btm_0[0] = {1'b0,layer_3_0[3679:3672]} - {1'b0, layer_2_0[3679:3672]};
      btm_0[1] = {1'b0,layer_3_0[3687:3680]} - {1'b0, layer_2_0[3687:3680]};
      btm_0[2] = {1'b0,layer_3_0[3695:3688]} - {1'b0, layer_2_0[3695:3688]};
      btm_1[0] = {1'b0,layer_3_1[3679:3672]} - {1'b0, layer_2_1[3679:3672]};
      btm_1[1] = {1'b0,layer_3_1[3687:3680]} - {1'b0, layer_2_1[3687:3680]};
      btm_1[2] = {1'b0,layer_3_1[3695:3688]} - {1'b0, layer_2_1[3695:3688]};
      btm_2[0] = {1'b0,layer_3_2[3679:3672]} - {1'b0, layer_2_2[3679:3672]};
      btm_2[1] = {1'b0,layer_3_2[3687:3680]} - {1'b0, layer_2_2[3687:3680]};
      btm_2[2] = {1'b0,layer_3_2[3695:3688]} - {1'b0, layer_2_2[3695:3688]};
    end
    'd461: begin
      top_0[0] = {1'b0,layer_1_0[3687:3680]} - {1'b0, layer_0_0[3687:3680]};
      top_0[1] = {1'b0,layer_1_0[3695:3688]} - {1'b0, layer_0_0[3695:3688]};
      top_0[2] = {1'b0,layer_1_0[3703:3696]} - {1'b0, layer_0_0[3703:3696]};
      top_1[0] = {1'b0,layer_1_1[3687:3680]} - {1'b0, layer_0_1[3687:3680]};
      top_1[1] = {1'b0,layer_1_1[3695:3688]} - {1'b0, layer_0_1[3695:3688]};
      top_1[2] = {1'b0,layer_1_1[3703:3696]} - {1'b0, layer_0_1[3703:3696]};
      top_2[0] = {1'b0,layer_1_2[3687:3680]} - {1'b0, layer_0_2[3687:3680]};
      top_2[1] = {1'b0,layer_1_2[3695:3688]} - {1'b0, layer_0_2[3695:3688]};
      top_2[2] = {1'b0,layer_1_2[3703:3696]} - {1'b0, layer_0_2[3703:3696]};
      mid_0[0] = {1'b0,layer_2_0[3687:3680]} - {1'b0, layer_1_0[3687:3680]};
      mid_0[1] = {1'b0,layer_2_0[3695:3688]} - {1'b0, layer_1_0[3695:3688]};
      mid_0[2] = {1'b0,layer_2_0[3703:3696]} - {1'b0, layer_1_0[3703:3696]};
      mid_1[0] = {1'b0,layer_2_1[3687:3680]} - {1'b0, layer_1_1[3687:3680]};
      mid_1[1] = {1'b0,layer_2_1[3695:3688]} - {1'b0, layer_1_1[3695:3688]};
      mid_1[2] = {1'b0,layer_2_1[3703:3696]} - {1'b0, layer_1_1[3703:3696]};
      mid_2[0] = {1'b0,layer_2_2[3687:3680]} - {1'b0, layer_1_2[3687:3680]};
      mid_2[1] = {1'b0,layer_2_2[3695:3688]} - {1'b0, layer_1_2[3695:3688]};
      mid_2[2] = {1'b0,layer_2_2[3703:3696]} - {1'b0, layer_1_2[3703:3696]};
      btm_0[0] = {1'b0,layer_3_0[3687:3680]} - {1'b0, layer_2_0[3687:3680]};
      btm_0[1] = {1'b0,layer_3_0[3695:3688]} - {1'b0, layer_2_0[3695:3688]};
      btm_0[2] = {1'b0,layer_3_0[3703:3696]} - {1'b0, layer_2_0[3703:3696]};
      btm_1[0] = {1'b0,layer_3_1[3687:3680]} - {1'b0, layer_2_1[3687:3680]};
      btm_1[1] = {1'b0,layer_3_1[3695:3688]} - {1'b0, layer_2_1[3695:3688]};
      btm_1[2] = {1'b0,layer_3_1[3703:3696]} - {1'b0, layer_2_1[3703:3696]};
      btm_2[0] = {1'b0,layer_3_2[3687:3680]} - {1'b0, layer_2_2[3687:3680]};
      btm_2[1] = {1'b0,layer_3_2[3695:3688]} - {1'b0, layer_2_2[3695:3688]};
      btm_2[2] = {1'b0,layer_3_2[3703:3696]} - {1'b0, layer_2_2[3703:3696]};
    end
    'd462: begin
      top_0[0] = {1'b0,layer_1_0[3695:3688]} - {1'b0, layer_0_0[3695:3688]};
      top_0[1] = {1'b0,layer_1_0[3703:3696]} - {1'b0, layer_0_0[3703:3696]};
      top_0[2] = {1'b0,layer_1_0[3711:3704]} - {1'b0, layer_0_0[3711:3704]};
      top_1[0] = {1'b0,layer_1_1[3695:3688]} - {1'b0, layer_0_1[3695:3688]};
      top_1[1] = {1'b0,layer_1_1[3703:3696]} - {1'b0, layer_0_1[3703:3696]};
      top_1[2] = {1'b0,layer_1_1[3711:3704]} - {1'b0, layer_0_1[3711:3704]};
      top_2[0] = {1'b0,layer_1_2[3695:3688]} - {1'b0, layer_0_2[3695:3688]};
      top_2[1] = {1'b0,layer_1_2[3703:3696]} - {1'b0, layer_0_2[3703:3696]};
      top_2[2] = {1'b0,layer_1_2[3711:3704]} - {1'b0, layer_0_2[3711:3704]};
      mid_0[0] = {1'b0,layer_2_0[3695:3688]} - {1'b0, layer_1_0[3695:3688]};
      mid_0[1] = {1'b0,layer_2_0[3703:3696]} - {1'b0, layer_1_0[3703:3696]};
      mid_0[2] = {1'b0,layer_2_0[3711:3704]} - {1'b0, layer_1_0[3711:3704]};
      mid_1[0] = {1'b0,layer_2_1[3695:3688]} - {1'b0, layer_1_1[3695:3688]};
      mid_1[1] = {1'b0,layer_2_1[3703:3696]} - {1'b0, layer_1_1[3703:3696]};
      mid_1[2] = {1'b0,layer_2_1[3711:3704]} - {1'b0, layer_1_1[3711:3704]};
      mid_2[0] = {1'b0,layer_2_2[3695:3688]} - {1'b0, layer_1_2[3695:3688]};
      mid_2[1] = {1'b0,layer_2_2[3703:3696]} - {1'b0, layer_1_2[3703:3696]};
      mid_2[2] = {1'b0,layer_2_2[3711:3704]} - {1'b0, layer_1_2[3711:3704]};
      btm_0[0] = {1'b0,layer_3_0[3695:3688]} - {1'b0, layer_2_0[3695:3688]};
      btm_0[1] = {1'b0,layer_3_0[3703:3696]} - {1'b0, layer_2_0[3703:3696]};
      btm_0[2] = {1'b0,layer_3_0[3711:3704]} - {1'b0, layer_2_0[3711:3704]};
      btm_1[0] = {1'b0,layer_3_1[3695:3688]} - {1'b0, layer_2_1[3695:3688]};
      btm_1[1] = {1'b0,layer_3_1[3703:3696]} - {1'b0, layer_2_1[3703:3696]};
      btm_1[2] = {1'b0,layer_3_1[3711:3704]} - {1'b0, layer_2_1[3711:3704]};
      btm_2[0] = {1'b0,layer_3_2[3695:3688]} - {1'b0, layer_2_2[3695:3688]};
      btm_2[1] = {1'b0,layer_3_2[3703:3696]} - {1'b0, layer_2_2[3703:3696]};
      btm_2[2] = {1'b0,layer_3_2[3711:3704]} - {1'b0, layer_2_2[3711:3704]};
    end
    'd463: begin
      top_0[0] = {1'b0,layer_1_0[3703:3696]} - {1'b0, layer_0_0[3703:3696]};
      top_0[1] = {1'b0,layer_1_0[3711:3704]} - {1'b0, layer_0_0[3711:3704]};
      top_0[2] = {1'b0,layer_1_0[3719:3712]} - {1'b0, layer_0_0[3719:3712]};
      top_1[0] = {1'b0,layer_1_1[3703:3696]} - {1'b0, layer_0_1[3703:3696]};
      top_1[1] = {1'b0,layer_1_1[3711:3704]} - {1'b0, layer_0_1[3711:3704]};
      top_1[2] = {1'b0,layer_1_1[3719:3712]} - {1'b0, layer_0_1[3719:3712]};
      top_2[0] = {1'b0,layer_1_2[3703:3696]} - {1'b0, layer_0_2[3703:3696]};
      top_2[1] = {1'b0,layer_1_2[3711:3704]} - {1'b0, layer_0_2[3711:3704]};
      top_2[2] = {1'b0,layer_1_2[3719:3712]} - {1'b0, layer_0_2[3719:3712]};
      mid_0[0] = {1'b0,layer_2_0[3703:3696]} - {1'b0, layer_1_0[3703:3696]};
      mid_0[1] = {1'b0,layer_2_0[3711:3704]} - {1'b0, layer_1_0[3711:3704]};
      mid_0[2] = {1'b0,layer_2_0[3719:3712]} - {1'b0, layer_1_0[3719:3712]};
      mid_1[0] = {1'b0,layer_2_1[3703:3696]} - {1'b0, layer_1_1[3703:3696]};
      mid_1[1] = {1'b0,layer_2_1[3711:3704]} - {1'b0, layer_1_1[3711:3704]};
      mid_1[2] = {1'b0,layer_2_1[3719:3712]} - {1'b0, layer_1_1[3719:3712]};
      mid_2[0] = {1'b0,layer_2_2[3703:3696]} - {1'b0, layer_1_2[3703:3696]};
      mid_2[1] = {1'b0,layer_2_2[3711:3704]} - {1'b0, layer_1_2[3711:3704]};
      mid_2[2] = {1'b0,layer_2_2[3719:3712]} - {1'b0, layer_1_2[3719:3712]};
      btm_0[0] = {1'b0,layer_3_0[3703:3696]} - {1'b0, layer_2_0[3703:3696]};
      btm_0[1] = {1'b0,layer_3_0[3711:3704]} - {1'b0, layer_2_0[3711:3704]};
      btm_0[2] = {1'b0,layer_3_0[3719:3712]} - {1'b0, layer_2_0[3719:3712]};
      btm_1[0] = {1'b0,layer_3_1[3703:3696]} - {1'b0, layer_2_1[3703:3696]};
      btm_1[1] = {1'b0,layer_3_1[3711:3704]} - {1'b0, layer_2_1[3711:3704]};
      btm_1[2] = {1'b0,layer_3_1[3719:3712]} - {1'b0, layer_2_1[3719:3712]};
      btm_2[0] = {1'b0,layer_3_2[3703:3696]} - {1'b0, layer_2_2[3703:3696]};
      btm_2[1] = {1'b0,layer_3_2[3711:3704]} - {1'b0, layer_2_2[3711:3704]};
      btm_2[2] = {1'b0,layer_3_2[3719:3712]} - {1'b0, layer_2_2[3719:3712]};
    end
    'd464: begin
      top_0[0] = {1'b0,layer_1_0[3711:3704]} - {1'b0, layer_0_0[3711:3704]};
      top_0[1] = {1'b0,layer_1_0[3719:3712]} - {1'b0, layer_0_0[3719:3712]};
      top_0[2] = {1'b0,layer_1_0[3727:3720]} - {1'b0, layer_0_0[3727:3720]};
      top_1[0] = {1'b0,layer_1_1[3711:3704]} - {1'b0, layer_0_1[3711:3704]};
      top_1[1] = {1'b0,layer_1_1[3719:3712]} - {1'b0, layer_0_1[3719:3712]};
      top_1[2] = {1'b0,layer_1_1[3727:3720]} - {1'b0, layer_0_1[3727:3720]};
      top_2[0] = {1'b0,layer_1_2[3711:3704]} - {1'b0, layer_0_2[3711:3704]};
      top_2[1] = {1'b0,layer_1_2[3719:3712]} - {1'b0, layer_0_2[3719:3712]};
      top_2[2] = {1'b0,layer_1_2[3727:3720]} - {1'b0, layer_0_2[3727:3720]};
      mid_0[0] = {1'b0,layer_2_0[3711:3704]} - {1'b0, layer_1_0[3711:3704]};
      mid_0[1] = {1'b0,layer_2_0[3719:3712]} - {1'b0, layer_1_0[3719:3712]};
      mid_0[2] = {1'b0,layer_2_0[3727:3720]} - {1'b0, layer_1_0[3727:3720]};
      mid_1[0] = {1'b0,layer_2_1[3711:3704]} - {1'b0, layer_1_1[3711:3704]};
      mid_1[1] = {1'b0,layer_2_1[3719:3712]} - {1'b0, layer_1_1[3719:3712]};
      mid_1[2] = {1'b0,layer_2_1[3727:3720]} - {1'b0, layer_1_1[3727:3720]};
      mid_2[0] = {1'b0,layer_2_2[3711:3704]} - {1'b0, layer_1_2[3711:3704]};
      mid_2[1] = {1'b0,layer_2_2[3719:3712]} - {1'b0, layer_1_2[3719:3712]};
      mid_2[2] = {1'b0,layer_2_2[3727:3720]} - {1'b0, layer_1_2[3727:3720]};
      btm_0[0] = {1'b0,layer_3_0[3711:3704]} - {1'b0, layer_2_0[3711:3704]};
      btm_0[1] = {1'b0,layer_3_0[3719:3712]} - {1'b0, layer_2_0[3719:3712]};
      btm_0[2] = {1'b0,layer_3_0[3727:3720]} - {1'b0, layer_2_0[3727:3720]};
      btm_1[0] = {1'b0,layer_3_1[3711:3704]} - {1'b0, layer_2_1[3711:3704]};
      btm_1[1] = {1'b0,layer_3_1[3719:3712]} - {1'b0, layer_2_1[3719:3712]};
      btm_1[2] = {1'b0,layer_3_1[3727:3720]} - {1'b0, layer_2_1[3727:3720]};
      btm_2[0] = {1'b0,layer_3_2[3711:3704]} - {1'b0, layer_2_2[3711:3704]};
      btm_2[1] = {1'b0,layer_3_2[3719:3712]} - {1'b0, layer_2_2[3719:3712]};
      btm_2[2] = {1'b0,layer_3_2[3727:3720]} - {1'b0, layer_2_2[3727:3720]};
    end
    'd465: begin
      top_0[0] = {1'b0,layer_1_0[3719:3712]} - {1'b0, layer_0_0[3719:3712]};
      top_0[1] = {1'b0,layer_1_0[3727:3720]} - {1'b0, layer_0_0[3727:3720]};
      top_0[2] = {1'b0,layer_1_0[3735:3728]} - {1'b0, layer_0_0[3735:3728]};
      top_1[0] = {1'b0,layer_1_1[3719:3712]} - {1'b0, layer_0_1[3719:3712]};
      top_1[1] = {1'b0,layer_1_1[3727:3720]} - {1'b0, layer_0_1[3727:3720]};
      top_1[2] = {1'b0,layer_1_1[3735:3728]} - {1'b0, layer_0_1[3735:3728]};
      top_2[0] = {1'b0,layer_1_2[3719:3712]} - {1'b0, layer_0_2[3719:3712]};
      top_2[1] = {1'b0,layer_1_2[3727:3720]} - {1'b0, layer_0_2[3727:3720]};
      top_2[2] = {1'b0,layer_1_2[3735:3728]} - {1'b0, layer_0_2[3735:3728]};
      mid_0[0] = {1'b0,layer_2_0[3719:3712]} - {1'b0, layer_1_0[3719:3712]};
      mid_0[1] = {1'b0,layer_2_0[3727:3720]} - {1'b0, layer_1_0[3727:3720]};
      mid_0[2] = {1'b0,layer_2_0[3735:3728]} - {1'b0, layer_1_0[3735:3728]};
      mid_1[0] = {1'b0,layer_2_1[3719:3712]} - {1'b0, layer_1_1[3719:3712]};
      mid_1[1] = {1'b0,layer_2_1[3727:3720]} - {1'b0, layer_1_1[3727:3720]};
      mid_1[2] = {1'b0,layer_2_1[3735:3728]} - {1'b0, layer_1_1[3735:3728]};
      mid_2[0] = {1'b0,layer_2_2[3719:3712]} - {1'b0, layer_1_2[3719:3712]};
      mid_2[1] = {1'b0,layer_2_2[3727:3720]} - {1'b0, layer_1_2[3727:3720]};
      mid_2[2] = {1'b0,layer_2_2[3735:3728]} - {1'b0, layer_1_2[3735:3728]};
      btm_0[0] = {1'b0,layer_3_0[3719:3712]} - {1'b0, layer_2_0[3719:3712]};
      btm_0[1] = {1'b0,layer_3_0[3727:3720]} - {1'b0, layer_2_0[3727:3720]};
      btm_0[2] = {1'b0,layer_3_0[3735:3728]} - {1'b0, layer_2_0[3735:3728]};
      btm_1[0] = {1'b0,layer_3_1[3719:3712]} - {1'b0, layer_2_1[3719:3712]};
      btm_1[1] = {1'b0,layer_3_1[3727:3720]} - {1'b0, layer_2_1[3727:3720]};
      btm_1[2] = {1'b0,layer_3_1[3735:3728]} - {1'b0, layer_2_1[3735:3728]};
      btm_2[0] = {1'b0,layer_3_2[3719:3712]} - {1'b0, layer_2_2[3719:3712]};
      btm_2[1] = {1'b0,layer_3_2[3727:3720]} - {1'b0, layer_2_2[3727:3720]};
      btm_2[2] = {1'b0,layer_3_2[3735:3728]} - {1'b0, layer_2_2[3735:3728]};
    end
    'd466: begin
      top_0[0] = {1'b0,layer_1_0[3727:3720]} - {1'b0, layer_0_0[3727:3720]};
      top_0[1] = {1'b0,layer_1_0[3735:3728]} - {1'b0, layer_0_0[3735:3728]};
      top_0[2] = {1'b0,layer_1_0[3743:3736]} - {1'b0, layer_0_0[3743:3736]};
      top_1[0] = {1'b0,layer_1_1[3727:3720]} - {1'b0, layer_0_1[3727:3720]};
      top_1[1] = {1'b0,layer_1_1[3735:3728]} - {1'b0, layer_0_1[3735:3728]};
      top_1[2] = {1'b0,layer_1_1[3743:3736]} - {1'b0, layer_0_1[3743:3736]};
      top_2[0] = {1'b0,layer_1_2[3727:3720]} - {1'b0, layer_0_2[3727:3720]};
      top_2[1] = {1'b0,layer_1_2[3735:3728]} - {1'b0, layer_0_2[3735:3728]};
      top_2[2] = {1'b0,layer_1_2[3743:3736]} - {1'b0, layer_0_2[3743:3736]};
      mid_0[0] = {1'b0,layer_2_0[3727:3720]} - {1'b0, layer_1_0[3727:3720]};
      mid_0[1] = {1'b0,layer_2_0[3735:3728]} - {1'b0, layer_1_0[3735:3728]};
      mid_0[2] = {1'b0,layer_2_0[3743:3736]} - {1'b0, layer_1_0[3743:3736]};
      mid_1[0] = {1'b0,layer_2_1[3727:3720]} - {1'b0, layer_1_1[3727:3720]};
      mid_1[1] = {1'b0,layer_2_1[3735:3728]} - {1'b0, layer_1_1[3735:3728]};
      mid_1[2] = {1'b0,layer_2_1[3743:3736]} - {1'b0, layer_1_1[3743:3736]};
      mid_2[0] = {1'b0,layer_2_2[3727:3720]} - {1'b0, layer_1_2[3727:3720]};
      mid_2[1] = {1'b0,layer_2_2[3735:3728]} - {1'b0, layer_1_2[3735:3728]};
      mid_2[2] = {1'b0,layer_2_2[3743:3736]} - {1'b0, layer_1_2[3743:3736]};
      btm_0[0] = {1'b0,layer_3_0[3727:3720]} - {1'b0, layer_2_0[3727:3720]};
      btm_0[1] = {1'b0,layer_3_0[3735:3728]} - {1'b0, layer_2_0[3735:3728]};
      btm_0[2] = {1'b0,layer_3_0[3743:3736]} - {1'b0, layer_2_0[3743:3736]};
      btm_1[0] = {1'b0,layer_3_1[3727:3720]} - {1'b0, layer_2_1[3727:3720]};
      btm_1[1] = {1'b0,layer_3_1[3735:3728]} - {1'b0, layer_2_1[3735:3728]};
      btm_1[2] = {1'b0,layer_3_1[3743:3736]} - {1'b0, layer_2_1[3743:3736]};
      btm_2[0] = {1'b0,layer_3_2[3727:3720]} - {1'b0, layer_2_2[3727:3720]};
      btm_2[1] = {1'b0,layer_3_2[3735:3728]} - {1'b0, layer_2_2[3735:3728]};
      btm_2[2] = {1'b0,layer_3_2[3743:3736]} - {1'b0, layer_2_2[3743:3736]};
    end
    'd467: begin
      top_0[0] = {1'b0,layer_1_0[3735:3728]} - {1'b0, layer_0_0[3735:3728]};
      top_0[1] = {1'b0,layer_1_0[3743:3736]} - {1'b0, layer_0_0[3743:3736]};
      top_0[2] = {1'b0,layer_1_0[3751:3744]} - {1'b0, layer_0_0[3751:3744]};
      top_1[0] = {1'b0,layer_1_1[3735:3728]} - {1'b0, layer_0_1[3735:3728]};
      top_1[1] = {1'b0,layer_1_1[3743:3736]} - {1'b0, layer_0_1[3743:3736]};
      top_1[2] = {1'b0,layer_1_1[3751:3744]} - {1'b0, layer_0_1[3751:3744]};
      top_2[0] = {1'b0,layer_1_2[3735:3728]} - {1'b0, layer_0_2[3735:3728]};
      top_2[1] = {1'b0,layer_1_2[3743:3736]} - {1'b0, layer_0_2[3743:3736]};
      top_2[2] = {1'b0,layer_1_2[3751:3744]} - {1'b0, layer_0_2[3751:3744]};
      mid_0[0] = {1'b0,layer_2_0[3735:3728]} - {1'b0, layer_1_0[3735:3728]};
      mid_0[1] = {1'b0,layer_2_0[3743:3736]} - {1'b0, layer_1_0[3743:3736]};
      mid_0[2] = {1'b0,layer_2_0[3751:3744]} - {1'b0, layer_1_0[3751:3744]};
      mid_1[0] = {1'b0,layer_2_1[3735:3728]} - {1'b0, layer_1_1[3735:3728]};
      mid_1[1] = {1'b0,layer_2_1[3743:3736]} - {1'b0, layer_1_1[3743:3736]};
      mid_1[2] = {1'b0,layer_2_1[3751:3744]} - {1'b0, layer_1_1[3751:3744]};
      mid_2[0] = {1'b0,layer_2_2[3735:3728]} - {1'b0, layer_1_2[3735:3728]};
      mid_2[1] = {1'b0,layer_2_2[3743:3736]} - {1'b0, layer_1_2[3743:3736]};
      mid_2[2] = {1'b0,layer_2_2[3751:3744]} - {1'b0, layer_1_2[3751:3744]};
      btm_0[0] = {1'b0,layer_3_0[3735:3728]} - {1'b0, layer_2_0[3735:3728]};
      btm_0[1] = {1'b0,layer_3_0[3743:3736]} - {1'b0, layer_2_0[3743:3736]};
      btm_0[2] = {1'b0,layer_3_0[3751:3744]} - {1'b0, layer_2_0[3751:3744]};
      btm_1[0] = {1'b0,layer_3_1[3735:3728]} - {1'b0, layer_2_1[3735:3728]};
      btm_1[1] = {1'b0,layer_3_1[3743:3736]} - {1'b0, layer_2_1[3743:3736]};
      btm_1[2] = {1'b0,layer_3_1[3751:3744]} - {1'b0, layer_2_1[3751:3744]};
      btm_2[0] = {1'b0,layer_3_2[3735:3728]} - {1'b0, layer_2_2[3735:3728]};
      btm_2[1] = {1'b0,layer_3_2[3743:3736]} - {1'b0, layer_2_2[3743:3736]};
      btm_2[2] = {1'b0,layer_3_2[3751:3744]} - {1'b0, layer_2_2[3751:3744]};
    end
    'd468: begin
      top_0[0] = {1'b0,layer_1_0[3743:3736]} - {1'b0, layer_0_0[3743:3736]};
      top_0[1] = {1'b0,layer_1_0[3751:3744]} - {1'b0, layer_0_0[3751:3744]};
      top_0[2] = {1'b0,layer_1_0[3759:3752]} - {1'b0, layer_0_0[3759:3752]};
      top_1[0] = {1'b0,layer_1_1[3743:3736]} - {1'b0, layer_0_1[3743:3736]};
      top_1[1] = {1'b0,layer_1_1[3751:3744]} - {1'b0, layer_0_1[3751:3744]};
      top_1[2] = {1'b0,layer_1_1[3759:3752]} - {1'b0, layer_0_1[3759:3752]};
      top_2[0] = {1'b0,layer_1_2[3743:3736]} - {1'b0, layer_0_2[3743:3736]};
      top_2[1] = {1'b0,layer_1_2[3751:3744]} - {1'b0, layer_0_2[3751:3744]};
      top_2[2] = {1'b0,layer_1_2[3759:3752]} - {1'b0, layer_0_2[3759:3752]};
      mid_0[0] = {1'b0,layer_2_0[3743:3736]} - {1'b0, layer_1_0[3743:3736]};
      mid_0[1] = {1'b0,layer_2_0[3751:3744]} - {1'b0, layer_1_0[3751:3744]};
      mid_0[2] = {1'b0,layer_2_0[3759:3752]} - {1'b0, layer_1_0[3759:3752]};
      mid_1[0] = {1'b0,layer_2_1[3743:3736]} - {1'b0, layer_1_1[3743:3736]};
      mid_1[1] = {1'b0,layer_2_1[3751:3744]} - {1'b0, layer_1_1[3751:3744]};
      mid_1[2] = {1'b0,layer_2_1[3759:3752]} - {1'b0, layer_1_1[3759:3752]};
      mid_2[0] = {1'b0,layer_2_2[3743:3736]} - {1'b0, layer_1_2[3743:3736]};
      mid_2[1] = {1'b0,layer_2_2[3751:3744]} - {1'b0, layer_1_2[3751:3744]};
      mid_2[2] = {1'b0,layer_2_2[3759:3752]} - {1'b0, layer_1_2[3759:3752]};
      btm_0[0] = {1'b0,layer_3_0[3743:3736]} - {1'b0, layer_2_0[3743:3736]};
      btm_0[1] = {1'b0,layer_3_0[3751:3744]} - {1'b0, layer_2_0[3751:3744]};
      btm_0[2] = {1'b0,layer_3_0[3759:3752]} - {1'b0, layer_2_0[3759:3752]};
      btm_1[0] = {1'b0,layer_3_1[3743:3736]} - {1'b0, layer_2_1[3743:3736]};
      btm_1[1] = {1'b0,layer_3_1[3751:3744]} - {1'b0, layer_2_1[3751:3744]};
      btm_1[2] = {1'b0,layer_3_1[3759:3752]} - {1'b0, layer_2_1[3759:3752]};
      btm_2[0] = {1'b0,layer_3_2[3743:3736]} - {1'b0, layer_2_2[3743:3736]};
      btm_2[1] = {1'b0,layer_3_2[3751:3744]} - {1'b0, layer_2_2[3751:3744]};
      btm_2[2] = {1'b0,layer_3_2[3759:3752]} - {1'b0, layer_2_2[3759:3752]};
    end
    'd469: begin
      top_0[0] = {1'b0,layer_1_0[3751:3744]} - {1'b0, layer_0_0[3751:3744]};
      top_0[1] = {1'b0,layer_1_0[3759:3752]} - {1'b0, layer_0_0[3759:3752]};
      top_0[2] = {1'b0,layer_1_0[3767:3760]} - {1'b0, layer_0_0[3767:3760]};
      top_1[0] = {1'b0,layer_1_1[3751:3744]} - {1'b0, layer_0_1[3751:3744]};
      top_1[1] = {1'b0,layer_1_1[3759:3752]} - {1'b0, layer_0_1[3759:3752]};
      top_1[2] = {1'b0,layer_1_1[3767:3760]} - {1'b0, layer_0_1[3767:3760]};
      top_2[0] = {1'b0,layer_1_2[3751:3744]} - {1'b0, layer_0_2[3751:3744]};
      top_2[1] = {1'b0,layer_1_2[3759:3752]} - {1'b0, layer_0_2[3759:3752]};
      top_2[2] = {1'b0,layer_1_2[3767:3760]} - {1'b0, layer_0_2[3767:3760]};
      mid_0[0] = {1'b0,layer_2_0[3751:3744]} - {1'b0, layer_1_0[3751:3744]};
      mid_0[1] = {1'b0,layer_2_0[3759:3752]} - {1'b0, layer_1_0[3759:3752]};
      mid_0[2] = {1'b0,layer_2_0[3767:3760]} - {1'b0, layer_1_0[3767:3760]};
      mid_1[0] = {1'b0,layer_2_1[3751:3744]} - {1'b0, layer_1_1[3751:3744]};
      mid_1[1] = {1'b0,layer_2_1[3759:3752]} - {1'b0, layer_1_1[3759:3752]};
      mid_1[2] = {1'b0,layer_2_1[3767:3760]} - {1'b0, layer_1_1[3767:3760]};
      mid_2[0] = {1'b0,layer_2_2[3751:3744]} - {1'b0, layer_1_2[3751:3744]};
      mid_2[1] = {1'b0,layer_2_2[3759:3752]} - {1'b0, layer_1_2[3759:3752]};
      mid_2[2] = {1'b0,layer_2_2[3767:3760]} - {1'b0, layer_1_2[3767:3760]};
      btm_0[0] = {1'b0,layer_3_0[3751:3744]} - {1'b0, layer_2_0[3751:3744]};
      btm_0[1] = {1'b0,layer_3_0[3759:3752]} - {1'b0, layer_2_0[3759:3752]};
      btm_0[2] = {1'b0,layer_3_0[3767:3760]} - {1'b0, layer_2_0[3767:3760]};
      btm_1[0] = {1'b0,layer_3_1[3751:3744]} - {1'b0, layer_2_1[3751:3744]};
      btm_1[1] = {1'b0,layer_3_1[3759:3752]} - {1'b0, layer_2_1[3759:3752]};
      btm_1[2] = {1'b0,layer_3_1[3767:3760]} - {1'b0, layer_2_1[3767:3760]};
      btm_2[0] = {1'b0,layer_3_2[3751:3744]} - {1'b0, layer_2_2[3751:3744]};
      btm_2[1] = {1'b0,layer_3_2[3759:3752]} - {1'b0, layer_2_2[3759:3752]};
      btm_2[2] = {1'b0,layer_3_2[3767:3760]} - {1'b0, layer_2_2[3767:3760]};
    end
    'd470: begin
      top_0[0] = {1'b0,layer_1_0[3759:3752]} - {1'b0, layer_0_0[3759:3752]};
      top_0[1] = {1'b0,layer_1_0[3767:3760]} - {1'b0, layer_0_0[3767:3760]};
      top_0[2] = {1'b0,layer_1_0[3775:3768]} - {1'b0, layer_0_0[3775:3768]};
      top_1[0] = {1'b0,layer_1_1[3759:3752]} - {1'b0, layer_0_1[3759:3752]};
      top_1[1] = {1'b0,layer_1_1[3767:3760]} - {1'b0, layer_0_1[3767:3760]};
      top_1[2] = {1'b0,layer_1_1[3775:3768]} - {1'b0, layer_0_1[3775:3768]};
      top_2[0] = {1'b0,layer_1_2[3759:3752]} - {1'b0, layer_0_2[3759:3752]};
      top_2[1] = {1'b0,layer_1_2[3767:3760]} - {1'b0, layer_0_2[3767:3760]};
      top_2[2] = {1'b0,layer_1_2[3775:3768]} - {1'b0, layer_0_2[3775:3768]};
      mid_0[0] = {1'b0,layer_2_0[3759:3752]} - {1'b0, layer_1_0[3759:3752]};
      mid_0[1] = {1'b0,layer_2_0[3767:3760]} - {1'b0, layer_1_0[3767:3760]};
      mid_0[2] = {1'b0,layer_2_0[3775:3768]} - {1'b0, layer_1_0[3775:3768]};
      mid_1[0] = {1'b0,layer_2_1[3759:3752]} - {1'b0, layer_1_1[3759:3752]};
      mid_1[1] = {1'b0,layer_2_1[3767:3760]} - {1'b0, layer_1_1[3767:3760]};
      mid_1[2] = {1'b0,layer_2_1[3775:3768]} - {1'b0, layer_1_1[3775:3768]};
      mid_2[0] = {1'b0,layer_2_2[3759:3752]} - {1'b0, layer_1_2[3759:3752]};
      mid_2[1] = {1'b0,layer_2_2[3767:3760]} - {1'b0, layer_1_2[3767:3760]};
      mid_2[2] = {1'b0,layer_2_2[3775:3768]} - {1'b0, layer_1_2[3775:3768]};
      btm_0[0] = {1'b0,layer_3_0[3759:3752]} - {1'b0, layer_2_0[3759:3752]};
      btm_0[1] = {1'b0,layer_3_0[3767:3760]} - {1'b0, layer_2_0[3767:3760]};
      btm_0[2] = {1'b0,layer_3_0[3775:3768]} - {1'b0, layer_2_0[3775:3768]};
      btm_1[0] = {1'b0,layer_3_1[3759:3752]} - {1'b0, layer_2_1[3759:3752]};
      btm_1[1] = {1'b0,layer_3_1[3767:3760]} - {1'b0, layer_2_1[3767:3760]};
      btm_1[2] = {1'b0,layer_3_1[3775:3768]} - {1'b0, layer_2_1[3775:3768]};
      btm_2[0] = {1'b0,layer_3_2[3759:3752]} - {1'b0, layer_2_2[3759:3752]};
      btm_2[1] = {1'b0,layer_3_2[3767:3760]} - {1'b0, layer_2_2[3767:3760]};
      btm_2[2] = {1'b0,layer_3_2[3775:3768]} - {1'b0, layer_2_2[3775:3768]};
    end
    'd471: begin
      top_0[0] = {1'b0,layer_1_0[3767:3760]} - {1'b0, layer_0_0[3767:3760]};
      top_0[1] = {1'b0,layer_1_0[3775:3768]} - {1'b0, layer_0_0[3775:3768]};
      top_0[2] = {1'b0,layer_1_0[3783:3776]} - {1'b0, layer_0_0[3783:3776]};
      top_1[0] = {1'b0,layer_1_1[3767:3760]} - {1'b0, layer_0_1[3767:3760]};
      top_1[1] = {1'b0,layer_1_1[3775:3768]} - {1'b0, layer_0_1[3775:3768]};
      top_1[2] = {1'b0,layer_1_1[3783:3776]} - {1'b0, layer_0_1[3783:3776]};
      top_2[0] = {1'b0,layer_1_2[3767:3760]} - {1'b0, layer_0_2[3767:3760]};
      top_2[1] = {1'b0,layer_1_2[3775:3768]} - {1'b0, layer_0_2[3775:3768]};
      top_2[2] = {1'b0,layer_1_2[3783:3776]} - {1'b0, layer_0_2[3783:3776]};
      mid_0[0] = {1'b0,layer_2_0[3767:3760]} - {1'b0, layer_1_0[3767:3760]};
      mid_0[1] = {1'b0,layer_2_0[3775:3768]} - {1'b0, layer_1_0[3775:3768]};
      mid_0[2] = {1'b0,layer_2_0[3783:3776]} - {1'b0, layer_1_0[3783:3776]};
      mid_1[0] = {1'b0,layer_2_1[3767:3760]} - {1'b0, layer_1_1[3767:3760]};
      mid_1[1] = {1'b0,layer_2_1[3775:3768]} - {1'b0, layer_1_1[3775:3768]};
      mid_1[2] = {1'b0,layer_2_1[3783:3776]} - {1'b0, layer_1_1[3783:3776]};
      mid_2[0] = {1'b0,layer_2_2[3767:3760]} - {1'b0, layer_1_2[3767:3760]};
      mid_2[1] = {1'b0,layer_2_2[3775:3768]} - {1'b0, layer_1_2[3775:3768]};
      mid_2[2] = {1'b0,layer_2_2[3783:3776]} - {1'b0, layer_1_2[3783:3776]};
      btm_0[0] = {1'b0,layer_3_0[3767:3760]} - {1'b0, layer_2_0[3767:3760]};
      btm_0[1] = {1'b0,layer_3_0[3775:3768]} - {1'b0, layer_2_0[3775:3768]};
      btm_0[2] = {1'b0,layer_3_0[3783:3776]} - {1'b0, layer_2_0[3783:3776]};
      btm_1[0] = {1'b0,layer_3_1[3767:3760]} - {1'b0, layer_2_1[3767:3760]};
      btm_1[1] = {1'b0,layer_3_1[3775:3768]} - {1'b0, layer_2_1[3775:3768]};
      btm_1[2] = {1'b0,layer_3_1[3783:3776]} - {1'b0, layer_2_1[3783:3776]};
      btm_2[0] = {1'b0,layer_3_2[3767:3760]} - {1'b0, layer_2_2[3767:3760]};
      btm_2[1] = {1'b0,layer_3_2[3775:3768]} - {1'b0, layer_2_2[3775:3768]};
      btm_2[2] = {1'b0,layer_3_2[3783:3776]} - {1'b0, layer_2_2[3783:3776]};
    end
    'd472: begin
      top_0[0] = {1'b0,layer_1_0[3775:3768]} - {1'b0, layer_0_0[3775:3768]};
      top_0[1] = {1'b0,layer_1_0[3783:3776]} - {1'b0, layer_0_0[3783:3776]};
      top_0[2] = {1'b0,layer_1_0[3791:3784]} - {1'b0, layer_0_0[3791:3784]};
      top_1[0] = {1'b0,layer_1_1[3775:3768]} - {1'b0, layer_0_1[3775:3768]};
      top_1[1] = {1'b0,layer_1_1[3783:3776]} - {1'b0, layer_0_1[3783:3776]};
      top_1[2] = {1'b0,layer_1_1[3791:3784]} - {1'b0, layer_0_1[3791:3784]};
      top_2[0] = {1'b0,layer_1_2[3775:3768]} - {1'b0, layer_0_2[3775:3768]};
      top_2[1] = {1'b0,layer_1_2[3783:3776]} - {1'b0, layer_0_2[3783:3776]};
      top_2[2] = {1'b0,layer_1_2[3791:3784]} - {1'b0, layer_0_2[3791:3784]};
      mid_0[0] = {1'b0,layer_2_0[3775:3768]} - {1'b0, layer_1_0[3775:3768]};
      mid_0[1] = {1'b0,layer_2_0[3783:3776]} - {1'b0, layer_1_0[3783:3776]};
      mid_0[2] = {1'b0,layer_2_0[3791:3784]} - {1'b0, layer_1_0[3791:3784]};
      mid_1[0] = {1'b0,layer_2_1[3775:3768]} - {1'b0, layer_1_1[3775:3768]};
      mid_1[1] = {1'b0,layer_2_1[3783:3776]} - {1'b0, layer_1_1[3783:3776]};
      mid_1[2] = {1'b0,layer_2_1[3791:3784]} - {1'b0, layer_1_1[3791:3784]};
      mid_2[0] = {1'b0,layer_2_2[3775:3768]} - {1'b0, layer_1_2[3775:3768]};
      mid_2[1] = {1'b0,layer_2_2[3783:3776]} - {1'b0, layer_1_2[3783:3776]};
      mid_2[2] = {1'b0,layer_2_2[3791:3784]} - {1'b0, layer_1_2[3791:3784]};
      btm_0[0] = {1'b0,layer_3_0[3775:3768]} - {1'b0, layer_2_0[3775:3768]};
      btm_0[1] = {1'b0,layer_3_0[3783:3776]} - {1'b0, layer_2_0[3783:3776]};
      btm_0[2] = {1'b0,layer_3_0[3791:3784]} - {1'b0, layer_2_0[3791:3784]};
      btm_1[0] = {1'b0,layer_3_1[3775:3768]} - {1'b0, layer_2_1[3775:3768]};
      btm_1[1] = {1'b0,layer_3_1[3783:3776]} - {1'b0, layer_2_1[3783:3776]};
      btm_1[2] = {1'b0,layer_3_1[3791:3784]} - {1'b0, layer_2_1[3791:3784]};
      btm_2[0] = {1'b0,layer_3_2[3775:3768]} - {1'b0, layer_2_2[3775:3768]};
      btm_2[1] = {1'b0,layer_3_2[3783:3776]} - {1'b0, layer_2_2[3783:3776]};
      btm_2[2] = {1'b0,layer_3_2[3791:3784]} - {1'b0, layer_2_2[3791:3784]};
    end
    'd473: begin
      top_0[0] = {1'b0,layer_1_0[3783:3776]} - {1'b0, layer_0_0[3783:3776]};
      top_0[1] = {1'b0,layer_1_0[3791:3784]} - {1'b0, layer_0_0[3791:3784]};
      top_0[2] = {1'b0,layer_1_0[3799:3792]} - {1'b0, layer_0_0[3799:3792]};
      top_1[0] = {1'b0,layer_1_1[3783:3776]} - {1'b0, layer_0_1[3783:3776]};
      top_1[1] = {1'b0,layer_1_1[3791:3784]} - {1'b0, layer_0_1[3791:3784]};
      top_1[2] = {1'b0,layer_1_1[3799:3792]} - {1'b0, layer_0_1[3799:3792]};
      top_2[0] = {1'b0,layer_1_2[3783:3776]} - {1'b0, layer_0_2[3783:3776]};
      top_2[1] = {1'b0,layer_1_2[3791:3784]} - {1'b0, layer_0_2[3791:3784]};
      top_2[2] = {1'b0,layer_1_2[3799:3792]} - {1'b0, layer_0_2[3799:3792]};
      mid_0[0] = {1'b0,layer_2_0[3783:3776]} - {1'b0, layer_1_0[3783:3776]};
      mid_0[1] = {1'b0,layer_2_0[3791:3784]} - {1'b0, layer_1_0[3791:3784]};
      mid_0[2] = {1'b0,layer_2_0[3799:3792]} - {1'b0, layer_1_0[3799:3792]};
      mid_1[0] = {1'b0,layer_2_1[3783:3776]} - {1'b0, layer_1_1[3783:3776]};
      mid_1[1] = {1'b0,layer_2_1[3791:3784]} - {1'b0, layer_1_1[3791:3784]};
      mid_1[2] = {1'b0,layer_2_1[3799:3792]} - {1'b0, layer_1_1[3799:3792]};
      mid_2[0] = {1'b0,layer_2_2[3783:3776]} - {1'b0, layer_1_2[3783:3776]};
      mid_2[1] = {1'b0,layer_2_2[3791:3784]} - {1'b0, layer_1_2[3791:3784]};
      mid_2[2] = {1'b0,layer_2_2[3799:3792]} - {1'b0, layer_1_2[3799:3792]};
      btm_0[0] = {1'b0,layer_3_0[3783:3776]} - {1'b0, layer_2_0[3783:3776]};
      btm_0[1] = {1'b0,layer_3_0[3791:3784]} - {1'b0, layer_2_0[3791:3784]};
      btm_0[2] = {1'b0,layer_3_0[3799:3792]} - {1'b0, layer_2_0[3799:3792]};
      btm_1[0] = {1'b0,layer_3_1[3783:3776]} - {1'b0, layer_2_1[3783:3776]};
      btm_1[1] = {1'b0,layer_3_1[3791:3784]} - {1'b0, layer_2_1[3791:3784]};
      btm_1[2] = {1'b0,layer_3_1[3799:3792]} - {1'b0, layer_2_1[3799:3792]};
      btm_2[0] = {1'b0,layer_3_2[3783:3776]} - {1'b0, layer_2_2[3783:3776]};
      btm_2[1] = {1'b0,layer_3_2[3791:3784]} - {1'b0, layer_2_2[3791:3784]};
      btm_2[2] = {1'b0,layer_3_2[3799:3792]} - {1'b0, layer_2_2[3799:3792]};
    end
    'd474: begin
      top_0[0] = {1'b0,layer_1_0[3791:3784]} - {1'b0, layer_0_0[3791:3784]};
      top_0[1] = {1'b0,layer_1_0[3799:3792]} - {1'b0, layer_0_0[3799:3792]};
      top_0[2] = {1'b0,layer_1_0[3807:3800]} - {1'b0, layer_0_0[3807:3800]};
      top_1[0] = {1'b0,layer_1_1[3791:3784]} - {1'b0, layer_0_1[3791:3784]};
      top_1[1] = {1'b0,layer_1_1[3799:3792]} - {1'b0, layer_0_1[3799:3792]};
      top_1[2] = {1'b0,layer_1_1[3807:3800]} - {1'b0, layer_0_1[3807:3800]};
      top_2[0] = {1'b0,layer_1_2[3791:3784]} - {1'b0, layer_0_2[3791:3784]};
      top_2[1] = {1'b0,layer_1_2[3799:3792]} - {1'b0, layer_0_2[3799:3792]};
      top_2[2] = {1'b0,layer_1_2[3807:3800]} - {1'b0, layer_0_2[3807:3800]};
      mid_0[0] = {1'b0,layer_2_0[3791:3784]} - {1'b0, layer_1_0[3791:3784]};
      mid_0[1] = {1'b0,layer_2_0[3799:3792]} - {1'b0, layer_1_0[3799:3792]};
      mid_0[2] = {1'b0,layer_2_0[3807:3800]} - {1'b0, layer_1_0[3807:3800]};
      mid_1[0] = {1'b0,layer_2_1[3791:3784]} - {1'b0, layer_1_1[3791:3784]};
      mid_1[1] = {1'b0,layer_2_1[3799:3792]} - {1'b0, layer_1_1[3799:3792]};
      mid_1[2] = {1'b0,layer_2_1[3807:3800]} - {1'b0, layer_1_1[3807:3800]};
      mid_2[0] = {1'b0,layer_2_2[3791:3784]} - {1'b0, layer_1_2[3791:3784]};
      mid_2[1] = {1'b0,layer_2_2[3799:3792]} - {1'b0, layer_1_2[3799:3792]};
      mid_2[2] = {1'b0,layer_2_2[3807:3800]} - {1'b0, layer_1_2[3807:3800]};
      btm_0[0] = {1'b0,layer_3_0[3791:3784]} - {1'b0, layer_2_0[3791:3784]};
      btm_0[1] = {1'b0,layer_3_0[3799:3792]} - {1'b0, layer_2_0[3799:3792]};
      btm_0[2] = {1'b0,layer_3_0[3807:3800]} - {1'b0, layer_2_0[3807:3800]};
      btm_1[0] = {1'b0,layer_3_1[3791:3784]} - {1'b0, layer_2_1[3791:3784]};
      btm_1[1] = {1'b0,layer_3_1[3799:3792]} - {1'b0, layer_2_1[3799:3792]};
      btm_1[2] = {1'b0,layer_3_1[3807:3800]} - {1'b0, layer_2_1[3807:3800]};
      btm_2[0] = {1'b0,layer_3_2[3791:3784]} - {1'b0, layer_2_2[3791:3784]};
      btm_2[1] = {1'b0,layer_3_2[3799:3792]} - {1'b0, layer_2_2[3799:3792]};
      btm_2[2] = {1'b0,layer_3_2[3807:3800]} - {1'b0, layer_2_2[3807:3800]};
    end
    'd475: begin
      top_0[0] = {1'b0,layer_1_0[3799:3792]} - {1'b0, layer_0_0[3799:3792]};
      top_0[1] = {1'b0,layer_1_0[3807:3800]} - {1'b0, layer_0_0[3807:3800]};
      top_0[2] = {1'b0,layer_1_0[3815:3808]} - {1'b0, layer_0_0[3815:3808]};
      top_1[0] = {1'b0,layer_1_1[3799:3792]} - {1'b0, layer_0_1[3799:3792]};
      top_1[1] = {1'b0,layer_1_1[3807:3800]} - {1'b0, layer_0_1[3807:3800]};
      top_1[2] = {1'b0,layer_1_1[3815:3808]} - {1'b0, layer_0_1[3815:3808]};
      top_2[0] = {1'b0,layer_1_2[3799:3792]} - {1'b0, layer_0_2[3799:3792]};
      top_2[1] = {1'b0,layer_1_2[3807:3800]} - {1'b0, layer_0_2[3807:3800]};
      top_2[2] = {1'b0,layer_1_2[3815:3808]} - {1'b0, layer_0_2[3815:3808]};
      mid_0[0] = {1'b0,layer_2_0[3799:3792]} - {1'b0, layer_1_0[3799:3792]};
      mid_0[1] = {1'b0,layer_2_0[3807:3800]} - {1'b0, layer_1_0[3807:3800]};
      mid_0[2] = {1'b0,layer_2_0[3815:3808]} - {1'b0, layer_1_0[3815:3808]};
      mid_1[0] = {1'b0,layer_2_1[3799:3792]} - {1'b0, layer_1_1[3799:3792]};
      mid_1[1] = {1'b0,layer_2_1[3807:3800]} - {1'b0, layer_1_1[3807:3800]};
      mid_1[2] = {1'b0,layer_2_1[3815:3808]} - {1'b0, layer_1_1[3815:3808]};
      mid_2[0] = {1'b0,layer_2_2[3799:3792]} - {1'b0, layer_1_2[3799:3792]};
      mid_2[1] = {1'b0,layer_2_2[3807:3800]} - {1'b0, layer_1_2[3807:3800]};
      mid_2[2] = {1'b0,layer_2_2[3815:3808]} - {1'b0, layer_1_2[3815:3808]};
      btm_0[0] = {1'b0,layer_3_0[3799:3792]} - {1'b0, layer_2_0[3799:3792]};
      btm_0[1] = {1'b0,layer_3_0[3807:3800]} - {1'b0, layer_2_0[3807:3800]};
      btm_0[2] = {1'b0,layer_3_0[3815:3808]} - {1'b0, layer_2_0[3815:3808]};
      btm_1[0] = {1'b0,layer_3_1[3799:3792]} - {1'b0, layer_2_1[3799:3792]};
      btm_1[1] = {1'b0,layer_3_1[3807:3800]} - {1'b0, layer_2_1[3807:3800]};
      btm_1[2] = {1'b0,layer_3_1[3815:3808]} - {1'b0, layer_2_1[3815:3808]};
      btm_2[0] = {1'b0,layer_3_2[3799:3792]} - {1'b0, layer_2_2[3799:3792]};
      btm_2[1] = {1'b0,layer_3_2[3807:3800]} - {1'b0, layer_2_2[3807:3800]};
      btm_2[2] = {1'b0,layer_3_2[3815:3808]} - {1'b0, layer_2_2[3815:3808]};
    end
    'd476: begin
      top_0[0] = {1'b0,layer_1_0[3807:3800]} - {1'b0, layer_0_0[3807:3800]};
      top_0[1] = {1'b0,layer_1_0[3815:3808]} - {1'b0, layer_0_0[3815:3808]};
      top_0[2] = {1'b0,layer_1_0[3823:3816]} - {1'b0, layer_0_0[3823:3816]};
      top_1[0] = {1'b0,layer_1_1[3807:3800]} - {1'b0, layer_0_1[3807:3800]};
      top_1[1] = {1'b0,layer_1_1[3815:3808]} - {1'b0, layer_0_1[3815:3808]};
      top_1[2] = {1'b0,layer_1_1[3823:3816]} - {1'b0, layer_0_1[3823:3816]};
      top_2[0] = {1'b0,layer_1_2[3807:3800]} - {1'b0, layer_0_2[3807:3800]};
      top_2[1] = {1'b0,layer_1_2[3815:3808]} - {1'b0, layer_0_2[3815:3808]};
      top_2[2] = {1'b0,layer_1_2[3823:3816]} - {1'b0, layer_0_2[3823:3816]};
      mid_0[0] = {1'b0,layer_2_0[3807:3800]} - {1'b0, layer_1_0[3807:3800]};
      mid_0[1] = {1'b0,layer_2_0[3815:3808]} - {1'b0, layer_1_0[3815:3808]};
      mid_0[2] = {1'b0,layer_2_0[3823:3816]} - {1'b0, layer_1_0[3823:3816]};
      mid_1[0] = {1'b0,layer_2_1[3807:3800]} - {1'b0, layer_1_1[3807:3800]};
      mid_1[1] = {1'b0,layer_2_1[3815:3808]} - {1'b0, layer_1_1[3815:3808]};
      mid_1[2] = {1'b0,layer_2_1[3823:3816]} - {1'b0, layer_1_1[3823:3816]};
      mid_2[0] = {1'b0,layer_2_2[3807:3800]} - {1'b0, layer_1_2[3807:3800]};
      mid_2[1] = {1'b0,layer_2_2[3815:3808]} - {1'b0, layer_1_2[3815:3808]};
      mid_2[2] = {1'b0,layer_2_2[3823:3816]} - {1'b0, layer_1_2[3823:3816]};
      btm_0[0] = {1'b0,layer_3_0[3807:3800]} - {1'b0, layer_2_0[3807:3800]};
      btm_0[1] = {1'b0,layer_3_0[3815:3808]} - {1'b0, layer_2_0[3815:3808]};
      btm_0[2] = {1'b0,layer_3_0[3823:3816]} - {1'b0, layer_2_0[3823:3816]};
      btm_1[0] = {1'b0,layer_3_1[3807:3800]} - {1'b0, layer_2_1[3807:3800]};
      btm_1[1] = {1'b0,layer_3_1[3815:3808]} - {1'b0, layer_2_1[3815:3808]};
      btm_1[2] = {1'b0,layer_3_1[3823:3816]} - {1'b0, layer_2_1[3823:3816]};
      btm_2[0] = {1'b0,layer_3_2[3807:3800]} - {1'b0, layer_2_2[3807:3800]};
      btm_2[1] = {1'b0,layer_3_2[3815:3808]} - {1'b0, layer_2_2[3815:3808]};
      btm_2[2] = {1'b0,layer_3_2[3823:3816]} - {1'b0, layer_2_2[3823:3816]};
    end
    'd477: begin
      top_0[0] = {1'b0,layer_1_0[3815:3808]} - {1'b0, layer_0_0[3815:3808]};
      top_0[1] = {1'b0,layer_1_0[3823:3816]} - {1'b0, layer_0_0[3823:3816]};
      top_0[2] = {1'b0,layer_1_0[3831:3824]} - {1'b0, layer_0_0[3831:3824]};
      top_1[0] = {1'b0,layer_1_1[3815:3808]} - {1'b0, layer_0_1[3815:3808]};
      top_1[1] = {1'b0,layer_1_1[3823:3816]} - {1'b0, layer_0_1[3823:3816]};
      top_1[2] = {1'b0,layer_1_1[3831:3824]} - {1'b0, layer_0_1[3831:3824]};
      top_2[0] = {1'b0,layer_1_2[3815:3808]} - {1'b0, layer_0_2[3815:3808]};
      top_2[1] = {1'b0,layer_1_2[3823:3816]} - {1'b0, layer_0_2[3823:3816]};
      top_2[2] = {1'b0,layer_1_2[3831:3824]} - {1'b0, layer_0_2[3831:3824]};
      mid_0[0] = {1'b0,layer_2_0[3815:3808]} - {1'b0, layer_1_0[3815:3808]};
      mid_0[1] = {1'b0,layer_2_0[3823:3816]} - {1'b0, layer_1_0[3823:3816]};
      mid_0[2] = {1'b0,layer_2_0[3831:3824]} - {1'b0, layer_1_0[3831:3824]};
      mid_1[0] = {1'b0,layer_2_1[3815:3808]} - {1'b0, layer_1_1[3815:3808]};
      mid_1[1] = {1'b0,layer_2_1[3823:3816]} - {1'b0, layer_1_1[3823:3816]};
      mid_1[2] = {1'b0,layer_2_1[3831:3824]} - {1'b0, layer_1_1[3831:3824]};
      mid_2[0] = {1'b0,layer_2_2[3815:3808]} - {1'b0, layer_1_2[3815:3808]};
      mid_2[1] = {1'b0,layer_2_2[3823:3816]} - {1'b0, layer_1_2[3823:3816]};
      mid_2[2] = {1'b0,layer_2_2[3831:3824]} - {1'b0, layer_1_2[3831:3824]};
      btm_0[0] = {1'b0,layer_3_0[3815:3808]} - {1'b0, layer_2_0[3815:3808]};
      btm_0[1] = {1'b0,layer_3_0[3823:3816]} - {1'b0, layer_2_0[3823:3816]};
      btm_0[2] = {1'b0,layer_3_0[3831:3824]} - {1'b0, layer_2_0[3831:3824]};
      btm_1[0] = {1'b0,layer_3_1[3815:3808]} - {1'b0, layer_2_1[3815:3808]};
      btm_1[1] = {1'b0,layer_3_1[3823:3816]} - {1'b0, layer_2_1[3823:3816]};
      btm_1[2] = {1'b0,layer_3_1[3831:3824]} - {1'b0, layer_2_1[3831:3824]};
      btm_2[0] = {1'b0,layer_3_2[3815:3808]} - {1'b0, layer_2_2[3815:3808]};
      btm_2[1] = {1'b0,layer_3_2[3823:3816]} - {1'b0, layer_2_2[3823:3816]};
      btm_2[2] = {1'b0,layer_3_2[3831:3824]} - {1'b0, layer_2_2[3831:3824]};
    end
    'd478: begin
      top_0[0] = {1'b0,layer_1_0[3823:3816]} - {1'b0, layer_0_0[3823:3816]};
      top_0[1] = {1'b0,layer_1_0[3831:3824]} - {1'b0, layer_0_0[3831:3824]};
      top_0[2] = {1'b0,layer_1_0[3839:3832]} - {1'b0, layer_0_0[3839:3832]};
      top_1[0] = {1'b0,layer_1_1[3823:3816]} - {1'b0, layer_0_1[3823:3816]};
      top_1[1] = {1'b0,layer_1_1[3831:3824]} - {1'b0, layer_0_1[3831:3824]};
      top_1[2] = {1'b0,layer_1_1[3839:3832]} - {1'b0, layer_0_1[3839:3832]};
      top_2[0] = {1'b0,layer_1_2[3823:3816]} - {1'b0, layer_0_2[3823:3816]};
      top_2[1] = {1'b0,layer_1_2[3831:3824]} - {1'b0, layer_0_2[3831:3824]};
      top_2[2] = {1'b0,layer_1_2[3839:3832]} - {1'b0, layer_0_2[3839:3832]};
      mid_0[0] = {1'b0,layer_2_0[3823:3816]} - {1'b0, layer_1_0[3823:3816]};
      mid_0[1] = {1'b0,layer_2_0[3831:3824]} - {1'b0, layer_1_0[3831:3824]};
      mid_0[2] = {1'b0,layer_2_0[3839:3832]} - {1'b0, layer_1_0[3839:3832]};
      mid_1[0] = {1'b0,layer_2_1[3823:3816]} - {1'b0, layer_1_1[3823:3816]};
      mid_1[1] = {1'b0,layer_2_1[3831:3824]} - {1'b0, layer_1_1[3831:3824]};
      mid_1[2] = {1'b0,layer_2_1[3839:3832]} - {1'b0, layer_1_1[3839:3832]};
      mid_2[0] = {1'b0,layer_2_2[3823:3816]} - {1'b0, layer_1_2[3823:3816]};
      mid_2[1] = {1'b0,layer_2_2[3831:3824]} - {1'b0, layer_1_2[3831:3824]};
      mid_2[2] = {1'b0,layer_2_2[3839:3832]} - {1'b0, layer_1_2[3839:3832]};
      btm_0[0] = {1'b0,layer_3_0[3823:3816]} - {1'b0, layer_2_0[3823:3816]};
      btm_0[1] = {1'b0,layer_3_0[3831:3824]} - {1'b0, layer_2_0[3831:3824]};
      btm_0[2] = {1'b0,layer_3_0[3839:3832]} - {1'b0, layer_2_0[3839:3832]};
      btm_1[0] = {1'b0,layer_3_1[3823:3816]} - {1'b0, layer_2_1[3823:3816]};
      btm_1[1] = {1'b0,layer_3_1[3831:3824]} - {1'b0, layer_2_1[3831:3824]};
      btm_1[2] = {1'b0,layer_3_1[3839:3832]} - {1'b0, layer_2_1[3839:3832]};
      btm_2[0] = {1'b0,layer_3_2[3823:3816]} - {1'b0, layer_2_2[3823:3816]};
      btm_2[1] = {1'b0,layer_3_2[3831:3824]} - {1'b0, layer_2_2[3831:3824]};
      btm_2[2] = {1'b0,layer_3_2[3839:3832]} - {1'b0, layer_2_2[3839:3832]};
    end
    'd479: begin
      top_0[0] = {1'b0,layer_1_0[3831:3824]} - {1'b0, layer_0_0[3831:3824]};
      top_0[1] = {1'b0,layer_1_0[3839:3832]} - {1'b0, layer_0_0[3839:3832]};
      top_0[2] = {1'b0,layer_1_0[3847:3840]} - {1'b0, layer_0_0[3847:3840]};
      top_1[0] = {1'b0,layer_1_1[3831:3824]} - {1'b0, layer_0_1[3831:3824]};
      top_1[1] = {1'b0,layer_1_1[3839:3832]} - {1'b0, layer_0_1[3839:3832]};
      top_1[2] = {1'b0,layer_1_1[3847:3840]} - {1'b0, layer_0_1[3847:3840]};
      top_2[0] = {1'b0,layer_1_2[3831:3824]} - {1'b0, layer_0_2[3831:3824]};
      top_2[1] = {1'b0,layer_1_2[3839:3832]} - {1'b0, layer_0_2[3839:3832]};
      top_2[2] = {1'b0,layer_1_2[3847:3840]} - {1'b0, layer_0_2[3847:3840]};
      mid_0[0] = {1'b0,layer_2_0[3831:3824]} - {1'b0, layer_1_0[3831:3824]};
      mid_0[1] = {1'b0,layer_2_0[3839:3832]} - {1'b0, layer_1_0[3839:3832]};
      mid_0[2] = {1'b0,layer_2_0[3847:3840]} - {1'b0, layer_1_0[3847:3840]};
      mid_1[0] = {1'b0,layer_2_1[3831:3824]} - {1'b0, layer_1_1[3831:3824]};
      mid_1[1] = {1'b0,layer_2_1[3839:3832]} - {1'b0, layer_1_1[3839:3832]};
      mid_1[2] = {1'b0,layer_2_1[3847:3840]} - {1'b0, layer_1_1[3847:3840]};
      mid_2[0] = {1'b0,layer_2_2[3831:3824]} - {1'b0, layer_1_2[3831:3824]};
      mid_2[1] = {1'b0,layer_2_2[3839:3832]} - {1'b0, layer_1_2[3839:3832]};
      mid_2[2] = {1'b0,layer_2_2[3847:3840]} - {1'b0, layer_1_2[3847:3840]};
      btm_0[0] = {1'b0,layer_3_0[3831:3824]} - {1'b0, layer_2_0[3831:3824]};
      btm_0[1] = {1'b0,layer_3_0[3839:3832]} - {1'b0, layer_2_0[3839:3832]};
      btm_0[2] = {1'b0,layer_3_0[3847:3840]} - {1'b0, layer_2_0[3847:3840]};
      btm_1[0] = {1'b0,layer_3_1[3831:3824]} - {1'b0, layer_2_1[3831:3824]};
      btm_1[1] = {1'b0,layer_3_1[3839:3832]} - {1'b0, layer_2_1[3839:3832]};
      btm_1[2] = {1'b0,layer_3_1[3847:3840]} - {1'b0, layer_2_1[3847:3840]};
      btm_2[0] = {1'b0,layer_3_2[3831:3824]} - {1'b0, layer_2_2[3831:3824]};
      btm_2[1] = {1'b0,layer_3_2[3839:3832]} - {1'b0, layer_2_2[3839:3832]};
      btm_2[2] = {1'b0,layer_3_2[3847:3840]} - {1'b0, layer_2_2[3847:3840]};
    end
    'd480: begin
      top_0[0] = {1'b0,layer_1_0[3839:3832]} - {1'b0, layer_0_0[3839:3832]};
      top_0[1] = {1'b0,layer_1_0[3847:3840]} - {1'b0, layer_0_0[3847:3840]};
      top_0[2] = {1'b0,layer_1_0[3855:3848]} - {1'b0, layer_0_0[3855:3848]};
      top_1[0] = {1'b0,layer_1_1[3839:3832]} - {1'b0, layer_0_1[3839:3832]};
      top_1[1] = {1'b0,layer_1_1[3847:3840]} - {1'b0, layer_0_1[3847:3840]};
      top_1[2] = {1'b0,layer_1_1[3855:3848]} - {1'b0, layer_0_1[3855:3848]};
      top_2[0] = {1'b0,layer_1_2[3839:3832]} - {1'b0, layer_0_2[3839:3832]};
      top_2[1] = {1'b0,layer_1_2[3847:3840]} - {1'b0, layer_0_2[3847:3840]};
      top_2[2] = {1'b0,layer_1_2[3855:3848]} - {1'b0, layer_0_2[3855:3848]};
      mid_0[0] = {1'b0,layer_2_0[3839:3832]} - {1'b0, layer_1_0[3839:3832]};
      mid_0[1] = {1'b0,layer_2_0[3847:3840]} - {1'b0, layer_1_0[3847:3840]};
      mid_0[2] = {1'b0,layer_2_0[3855:3848]} - {1'b0, layer_1_0[3855:3848]};
      mid_1[0] = {1'b0,layer_2_1[3839:3832]} - {1'b0, layer_1_1[3839:3832]};
      mid_1[1] = {1'b0,layer_2_1[3847:3840]} - {1'b0, layer_1_1[3847:3840]};
      mid_1[2] = {1'b0,layer_2_1[3855:3848]} - {1'b0, layer_1_1[3855:3848]};
      mid_2[0] = {1'b0,layer_2_2[3839:3832]} - {1'b0, layer_1_2[3839:3832]};
      mid_2[1] = {1'b0,layer_2_2[3847:3840]} - {1'b0, layer_1_2[3847:3840]};
      mid_2[2] = {1'b0,layer_2_2[3855:3848]} - {1'b0, layer_1_2[3855:3848]};
      btm_0[0] = {1'b0,layer_3_0[3839:3832]} - {1'b0, layer_2_0[3839:3832]};
      btm_0[1] = {1'b0,layer_3_0[3847:3840]} - {1'b0, layer_2_0[3847:3840]};
      btm_0[2] = {1'b0,layer_3_0[3855:3848]} - {1'b0, layer_2_0[3855:3848]};
      btm_1[0] = {1'b0,layer_3_1[3839:3832]} - {1'b0, layer_2_1[3839:3832]};
      btm_1[1] = {1'b0,layer_3_1[3847:3840]} - {1'b0, layer_2_1[3847:3840]};
      btm_1[2] = {1'b0,layer_3_1[3855:3848]} - {1'b0, layer_2_1[3855:3848]};
      btm_2[0] = {1'b0,layer_3_2[3839:3832]} - {1'b0, layer_2_2[3839:3832]};
      btm_2[1] = {1'b0,layer_3_2[3847:3840]} - {1'b0, layer_2_2[3847:3840]};
      btm_2[2] = {1'b0,layer_3_2[3855:3848]} - {1'b0, layer_2_2[3855:3848]};
    end
    'd481: begin
      top_0[0] = {1'b0,layer_1_0[3847:3840]} - {1'b0, layer_0_0[3847:3840]};
      top_0[1] = {1'b0,layer_1_0[3855:3848]} - {1'b0, layer_0_0[3855:3848]};
      top_0[2] = {1'b0,layer_1_0[3863:3856]} - {1'b0, layer_0_0[3863:3856]};
      top_1[0] = {1'b0,layer_1_1[3847:3840]} - {1'b0, layer_0_1[3847:3840]};
      top_1[1] = {1'b0,layer_1_1[3855:3848]} - {1'b0, layer_0_1[3855:3848]};
      top_1[2] = {1'b0,layer_1_1[3863:3856]} - {1'b0, layer_0_1[3863:3856]};
      top_2[0] = {1'b0,layer_1_2[3847:3840]} - {1'b0, layer_0_2[3847:3840]};
      top_2[1] = {1'b0,layer_1_2[3855:3848]} - {1'b0, layer_0_2[3855:3848]};
      top_2[2] = {1'b0,layer_1_2[3863:3856]} - {1'b0, layer_0_2[3863:3856]};
      mid_0[0] = {1'b0,layer_2_0[3847:3840]} - {1'b0, layer_1_0[3847:3840]};
      mid_0[1] = {1'b0,layer_2_0[3855:3848]} - {1'b0, layer_1_0[3855:3848]};
      mid_0[2] = {1'b0,layer_2_0[3863:3856]} - {1'b0, layer_1_0[3863:3856]};
      mid_1[0] = {1'b0,layer_2_1[3847:3840]} - {1'b0, layer_1_1[3847:3840]};
      mid_1[1] = {1'b0,layer_2_1[3855:3848]} - {1'b0, layer_1_1[3855:3848]};
      mid_1[2] = {1'b0,layer_2_1[3863:3856]} - {1'b0, layer_1_1[3863:3856]};
      mid_2[0] = {1'b0,layer_2_2[3847:3840]} - {1'b0, layer_1_2[3847:3840]};
      mid_2[1] = {1'b0,layer_2_2[3855:3848]} - {1'b0, layer_1_2[3855:3848]};
      mid_2[2] = {1'b0,layer_2_2[3863:3856]} - {1'b0, layer_1_2[3863:3856]};
      btm_0[0] = {1'b0,layer_3_0[3847:3840]} - {1'b0, layer_2_0[3847:3840]};
      btm_0[1] = {1'b0,layer_3_0[3855:3848]} - {1'b0, layer_2_0[3855:3848]};
      btm_0[2] = {1'b0,layer_3_0[3863:3856]} - {1'b0, layer_2_0[3863:3856]};
      btm_1[0] = {1'b0,layer_3_1[3847:3840]} - {1'b0, layer_2_1[3847:3840]};
      btm_1[1] = {1'b0,layer_3_1[3855:3848]} - {1'b0, layer_2_1[3855:3848]};
      btm_1[2] = {1'b0,layer_3_1[3863:3856]} - {1'b0, layer_2_1[3863:3856]};
      btm_2[0] = {1'b0,layer_3_2[3847:3840]} - {1'b0, layer_2_2[3847:3840]};
      btm_2[1] = {1'b0,layer_3_2[3855:3848]} - {1'b0, layer_2_2[3855:3848]};
      btm_2[2] = {1'b0,layer_3_2[3863:3856]} - {1'b0, layer_2_2[3863:3856]};
    end
    'd482: begin
      top_0[0] = {1'b0,layer_1_0[3855:3848]} - {1'b0, layer_0_0[3855:3848]};
      top_0[1] = {1'b0,layer_1_0[3863:3856]} - {1'b0, layer_0_0[3863:3856]};
      top_0[2] = {1'b0,layer_1_0[3871:3864]} - {1'b0, layer_0_0[3871:3864]};
      top_1[0] = {1'b0,layer_1_1[3855:3848]} - {1'b0, layer_0_1[3855:3848]};
      top_1[1] = {1'b0,layer_1_1[3863:3856]} - {1'b0, layer_0_1[3863:3856]};
      top_1[2] = {1'b0,layer_1_1[3871:3864]} - {1'b0, layer_0_1[3871:3864]};
      top_2[0] = {1'b0,layer_1_2[3855:3848]} - {1'b0, layer_0_2[3855:3848]};
      top_2[1] = {1'b0,layer_1_2[3863:3856]} - {1'b0, layer_0_2[3863:3856]};
      top_2[2] = {1'b0,layer_1_2[3871:3864]} - {1'b0, layer_0_2[3871:3864]};
      mid_0[0] = {1'b0,layer_2_0[3855:3848]} - {1'b0, layer_1_0[3855:3848]};
      mid_0[1] = {1'b0,layer_2_0[3863:3856]} - {1'b0, layer_1_0[3863:3856]};
      mid_0[2] = {1'b0,layer_2_0[3871:3864]} - {1'b0, layer_1_0[3871:3864]};
      mid_1[0] = {1'b0,layer_2_1[3855:3848]} - {1'b0, layer_1_1[3855:3848]};
      mid_1[1] = {1'b0,layer_2_1[3863:3856]} - {1'b0, layer_1_1[3863:3856]};
      mid_1[2] = {1'b0,layer_2_1[3871:3864]} - {1'b0, layer_1_1[3871:3864]};
      mid_2[0] = {1'b0,layer_2_2[3855:3848]} - {1'b0, layer_1_2[3855:3848]};
      mid_2[1] = {1'b0,layer_2_2[3863:3856]} - {1'b0, layer_1_2[3863:3856]};
      mid_2[2] = {1'b0,layer_2_2[3871:3864]} - {1'b0, layer_1_2[3871:3864]};
      btm_0[0] = {1'b0,layer_3_0[3855:3848]} - {1'b0, layer_2_0[3855:3848]};
      btm_0[1] = {1'b0,layer_3_0[3863:3856]} - {1'b0, layer_2_0[3863:3856]};
      btm_0[2] = {1'b0,layer_3_0[3871:3864]} - {1'b0, layer_2_0[3871:3864]};
      btm_1[0] = {1'b0,layer_3_1[3855:3848]} - {1'b0, layer_2_1[3855:3848]};
      btm_1[1] = {1'b0,layer_3_1[3863:3856]} - {1'b0, layer_2_1[3863:3856]};
      btm_1[2] = {1'b0,layer_3_1[3871:3864]} - {1'b0, layer_2_1[3871:3864]};
      btm_2[0] = {1'b0,layer_3_2[3855:3848]} - {1'b0, layer_2_2[3855:3848]};
      btm_2[1] = {1'b0,layer_3_2[3863:3856]} - {1'b0, layer_2_2[3863:3856]};
      btm_2[2] = {1'b0,layer_3_2[3871:3864]} - {1'b0, layer_2_2[3871:3864]};
    end
    'd483: begin
      top_0[0] = {1'b0,layer_1_0[3863:3856]} - {1'b0, layer_0_0[3863:3856]};
      top_0[1] = {1'b0,layer_1_0[3871:3864]} - {1'b0, layer_0_0[3871:3864]};
      top_0[2] = {1'b0,layer_1_0[3879:3872]} - {1'b0, layer_0_0[3879:3872]};
      top_1[0] = {1'b0,layer_1_1[3863:3856]} - {1'b0, layer_0_1[3863:3856]};
      top_1[1] = {1'b0,layer_1_1[3871:3864]} - {1'b0, layer_0_1[3871:3864]};
      top_1[2] = {1'b0,layer_1_1[3879:3872]} - {1'b0, layer_0_1[3879:3872]};
      top_2[0] = {1'b0,layer_1_2[3863:3856]} - {1'b0, layer_0_2[3863:3856]};
      top_2[1] = {1'b0,layer_1_2[3871:3864]} - {1'b0, layer_0_2[3871:3864]};
      top_2[2] = {1'b0,layer_1_2[3879:3872]} - {1'b0, layer_0_2[3879:3872]};
      mid_0[0] = {1'b0,layer_2_0[3863:3856]} - {1'b0, layer_1_0[3863:3856]};
      mid_0[1] = {1'b0,layer_2_0[3871:3864]} - {1'b0, layer_1_0[3871:3864]};
      mid_0[2] = {1'b0,layer_2_0[3879:3872]} - {1'b0, layer_1_0[3879:3872]};
      mid_1[0] = {1'b0,layer_2_1[3863:3856]} - {1'b0, layer_1_1[3863:3856]};
      mid_1[1] = {1'b0,layer_2_1[3871:3864]} - {1'b0, layer_1_1[3871:3864]};
      mid_1[2] = {1'b0,layer_2_1[3879:3872]} - {1'b0, layer_1_1[3879:3872]};
      mid_2[0] = {1'b0,layer_2_2[3863:3856]} - {1'b0, layer_1_2[3863:3856]};
      mid_2[1] = {1'b0,layer_2_2[3871:3864]} - {1'b0, layer_1_2[3871:3864]};
      mid_2[2] = {1'b0,layer_2_2[3879:3872]} - {1'b0, layer_1_2[3879:3872]};
      btm_0[0] = {1'b0,layer_3_0[3863:3856]} - {1'b0, layer_2_0[3863:3856]};
      btm_0[1] = {1'b0,layer_3_0[3871:3864]} - {1'b0, layer_2_0[3871:3864]};
      btm_0[2] = {1'b0,layer_3_0[3879:3872]} - {1'b0, layer_2_0[3879:3872]};
      btm_1[0] = {1'b0,layer_3_1[3863:3856]} - {1'b0, layer_2_1[3863:3856]};
      btm_1[1] = {1'b0,layer_3_1[3871:3864]} - {1'b0, layer_2_1[3871:3864]};
      btm_1[2] = {1'b0,layer_3_1[3879:3872]} - {1'b0, layer_2_1[3879:3872]};
      btm_2[0] = {1'b0,layer_3_2[3863:3856]} - {1'b0, layer_2_2[3863:3856]};
      btm_2[1] = {1'b0,layer_3_2[3871:3864]} - {1'b0, layer_2_2[3871:3864]};
      btm_2[2] = {1'b0,layer_3_2[3879:3872]} - {1'b0, layer_2_2[3879:3872]};
    end
    'd484: begin
      top_0[0] = {1'b0,layer_1_0[3871:3864]} - {1'b0, layer_0_0[3871:3864]};
      top_0[1] = {1'b0,layer_1_0[3879:3872]} - {1'b0, layer_0_0[3879:3872]};
      top_0[2] = {1'b0,layer_1_0[3887:3880]} - {1'b0, layer_0_0[3887:3880]};
      top_1[0] = {1'b0,layer_1_1[3871:3864]} - {1'b0, layer_0_1[3871:3864]};
      top_1[1] = {1'b0,layer_1_1[3879:3872]} - {1'b0, layer_0_1[3879:3872]};
      top_1[2] = {1'b0,layer_1_1[3887:3880]} - {1'b0, layer_0_1[3887:3880]};
      top_2[0] = {1'b0,layer_1_2[3871:3864]} - {1'b0, layer_0_2[3871:3864]};
      top_2[1] = {1'b0,layer_1_2[3879:3872]} - {1'b0, layer_0_2[3879:3872]};
      top_2[2] = {1'b0,layer_1_2[3887:3880]} - {1'b0, layer_0_2[3887:3880]};
      mid_0[0] = {1'b0,layer_2_0[3871:3864]} - {1'b0, layer_1_0[3871:3864]};
      mid_0[1] = {1'b0,layer_2_0[3879:3872]} - {1'b0, layer_1_0[3879:3872]};
      mid_0[2] = {1'b0,layer_2_0[3887:3880]} - {1'b0, layer_1_0[3887:3880]};
      mid_1[0] = {1'b0,layer_2_1[3871:3864]} - {1'b0, layer_1_1[3871:3864]};
      mid_1[1] = {1'b0,layer_2_1[3879:3872]} - {1'b0, layer_1_1[3879:3872]};
      mid_1[2] = {1'b0,layer_2_1[3887:3880]} - {1'b0, layer_1_1[3887:3880]};
      mid_2[0] = {1'b0,layer_2_2[3871:3864]} - {1'b0, layer_1_2[3871:3864]};
      mid_2[1] = {1'b0,layer_2_2[3879:3872]} - {1'b0, layer_1_2[3879:3872]};
      mid_2[2] = {1'b0,layer_2_2[3887:3880]} - {1'b0, layer_1_2[3887:3880]};
      btm_0[0] = {1'b0,layer_3_0[3871:3864]} - {1'b0, layer_2_0[3871:3864]};
      btm_0[1] = {1'b0,layer_3_0[3879:3872]} - {1'b0, layer_2_0[3879:3872]};
      btm_0[2] = {1'b0,layer_3_0[3887:3880]} - {1'b0, layer_2_0[3887:3880]};
      btm_1[0] = {1'b0,layer_3_1[3871:3864]} - {1'b0, layer_2_1[3871:3864]};
      btm_1[1] = {1'b0,layer_3_1[3879:3872]} - {1'b0, layer_2_1[3879:3872]};
      btm_1[2] = {1'b0,layer_3_1[3887:3880]} - {1'b0, layer_2_1[3887:3880]};
      btm_2[0] = {1'b0,layer_3_2[3871:3864]} - {1'b0, layer_2_2[3871:3864]};
      btm_2[1] = {1'b0,layer_3_2[3879:3872]} - {1'b0, layer_2_2[3879:3872]};
      btm_2[2] = {1'b0,layer_3_2[3887:3880]} - {1'b0, layer_2_2[3887:3880]};
    end
    'd485: begin
      top_0[0] = {1'b0,layer_1_0[3879:3872]} - {1'b0, layer_0_0[3879:3872]};
      top_0[1] = {1'b0,layer_1_0[3887:3880]} - {1'b0, layer_0_0[3887:3880]};
      top_0[2] = {1'b0,layer_1_0[3895:3888]} - {1'b0, layer_0_0[3895:3888]};
      top_1[0] = {1'b0,layer_1_1[3879:3872]} - {1'b0, layer_0_1[3879:3872]};
      top_1[1] = {1'b0,layer_1_1[3887:3880]} - {1'b0, layer_0_1[3887:3880]};
      top_1[2] = {1'b0,layer_1_1[3895:3888]} - {1'b0, layer_0_1[3895:3888]};
      top_2[0] = {1'b0,layer_1_2[3879:3872]} - {1'b0, layer_0_2[3879:3872]};
      top_2[1] = {1'b0,layer_1_2[3887:3880]} - {1'b0, layer_0_2[3887:3880]};
      top_2[2] = {1'b0,layer_1_2[3895:3888]} - {1'b0, layer_0_2[3895:3888]};
      mid_0[0] = {1'b0,layer_2_0[3879:3872]} - {1'b0, layer_1_0[3879:3872]};
      mid_0[1] = {1'b0,layer_2_0[3887:3880]} - {1'b0, layer_1_0[3887:3880]};
      mid_0[2] = {1'b0,layer_2_0[3895:3888]} - {1'b0, layer_1_0[3895:3888]};
      mid_1[0] = {1'b0,layer_2_1[3879:3872]} - {1'b0, layer_1_1[3879:3872]};
      mid_1[1] = {1'b0,layer_2_1[3887:3880]} - {1'b0, layer_1_1[3887:3880]};
      mid_1[2] = {1'b0,layer_2_1[3895:3888]} - {1'b0, layer_1_1[3895:3888]};
      mid_2[0] = {1'b0,layer_2_2[3879:3872]} - {1'b0, layer_1_2[3879:3872]};
      mid_2[1] = {1'b0,layer_2_2[3887:3880]} - {1'b0, layer_1_2[3887:3880]};
      mid_2[2] = {1'b0,layer_2_2[3895:3888]} - {1'b0, layer_1_2[3895:3888]};
      btm_0[0] = {1'b0,layer_3_0[3879:3872]} - {1'b0, layer_2_0[3879:3872]};
      btm_0[1] = {1'b0,layer_3_0[3887:3880]} - {1'b0, layer_2_0[3887:3880]};
      btm_0[2] = {1'b0,layer_3_0[3895:3888]} - {1'b0, layer_2_0[3895:3888]};
      btm_1[0] = {1'b0,layer_3_1[3879:3872]} - {1'b0, layer_2_1[3879:3872]};
      btm_1[1] = {1'b0,layer_3_1[3887:3880]} - {1'b0, layer_2_1[3887:3880]};
      btm_1[2] = {1'b0,layer_3_1[3895:3888]} - {1'b0, layer_2_1[3895:3888]};
      btm_2[0] = {1'b0,layer_3_2[3879:3872]} - {1'b0, layer_2_2[3879:3872]};
      btm_2[1] = {1'b0,layer_3_2[3887:3880]} - {1'b0, layer_2_2[3887:3880]};
      btm_2[2] = {1'b0,layer_3_2[3895:3888]} - {1'b0, layer_2_2[3895:3888]};
    end
    'd486: begin
      top_0[0] = {1'b0,layer_1_0[3887:3880]} - {1'b0, layer_0_0[3887:3880]};
      top_0[1] = {1'b0,layer_1_0[3895:3888]} - {1'b0, layer_0_0[3895:3888]};
      top_0[2] = {1'b0,layer_1_0[3903:3896]} - {1'b0, layer_0_0[3903:3896]};
      top_1[0] = {1'b0,layer_1_1[3887:3880]} - {1'b0, layer_0_1[3887:3880]};
      top_1[1] = {1'b0,layer_1_1[3895:3888]} - {1'b0, layer_0_1[3895:3888]};
      top_1[2] = {1'b0,layer_1_1[3903:3896]} - {1'b0, layer_0_1[3903:3896]};
      top_2[0] = {1'b0,layer_1_2[3887:3880]} - {1'b0, layer_0_2[3887:3880]};
      top_2[1] = {1'b0,layer_1_2[3895:3888]} - {1'b0, layer_0_2[3895:3888]};
      top_2[2] = {1'b0,layer_1_2[3903:3896]} - {1'b0, layer_0_2[3903:3896]};
      mid_0[0] = {1'b0,layer_2_0[3887:3880]} - {1'b0, layer_1_0[3887:3880]};
      mid_0[1] = {1'b0,layer_2_0[3895:3888]} - {1'b0, layer_1_0[3895:3888]};
      mid_0[2] = {1'b0,layer_2_0[3903:3896]} - {1'b0, layer_1_0[3903:3896]};
      mid_1[0] = {1'b0,layer_2_1[3887:3880]} - {1'b0, layer_1_1[3887:3880]};
      mid_1[1] = {1'b0,layer_2_1[3895:3888]} - {1'b0, layer_1_1[3895:3888]};
      mid_1[2] = {1'b0,layer_2_1[3903:3896]} - {1'b0, layer_1_1[3903:3896]};
      mid_2[0] = {1'b0,layer_2_2[3887:3880]} - {1'b0, layer_1_2[3887:3880]};
      mid_2[1] = {1'b0,layer_2_2[3895:3888]} - {1'b0, layer_1_2[3895:3888]};
      mid_2[2] = {1'b0,layer_2_2[3903:3896]} - {1'b0, layer_1_2[3903:3896]};
      btm_0[0] = {1'b0,layer_3_0[3887:3880]} - {1'b0, layer_2_0[3887:3880]};
      btm_0[1] = {1'b0,layer_3_0[3895:3888]} - {1'b0, layer_2_0[3895:3888]};
      btm_0[2] = {1'b0,layer_3_0[3903:3896]} - {1'b0, layer_2_0[3903:3896]};
      btm_1[0] = {1'b0,layer_3_1[3887:3880]} - {1'b0, layer_2_1[3887:3880]};
      btm_1[1] = {1'b0,layer_3_1[3895:3888]} - {1'b0, layer_2_1[3895:3888]};
      btm_1[2] = {1'b0,layer_3_1[3903:3896]} - {1'b0, layer_2_1[3903:3896]};
      btm_2[0] = {1'b0,layer_3_2[3887:3880]} - {1'b0, layer_2_2[3887:3880]};
      btm_2[1] = {1'b0,layer_3_2[3895:3888]} - {1'b0, layer_2_2[3895:3888]};
      btm_2[2] = {1'b0,layer_3_2[3903:3896]} - {1'b0, layer_2_2[3903:3896]};
    end
    'd487: begin
      top_0[0] = {1'b0,layer_1_0[3895:3888]} - {1'b0, layer_0_0[3895:3888]};
      top_0[1] = {1'b0,layer_1_0[3903:3896]} - {1'b0, layer_0_0[3903:3896]};
      top_0[2] = {1'b0,layer_1_0[3911:3904]} - {1'b0, layer_0_0[3911:3904]};
      top_1[0] = {1'b0,layer_1_1[3895:3888]} - {1'b0, layer_0_1[3895:3888]};
      top_1[1] = {1'b0,layer_1_1[3903:3896]} - {1'b0, layer_0_1[3903:3896]};
      top_1[2] = {1'b0,layer_1_1[3911:3904]} - {1'b0, layer_0_1[3911:3904]};
      top_2[0] = {1'b0,layer_1_2[3895:3888]} - {1'b0, layer_0_2[3895:3888]};
      top_2[1] = {1'b0,layer_1_2[3903:3896]} - {1'b0, layer_0_2[3903:3896]};
      top_2[2] = {1'b0,layer_1_2[3911:3904]} - {1'b0, layer_0_2[3911:3904]};
      mid_0[0] = {1'b0,layer_2_0[3895:3888]} - {1'b0, layer_1_0[3895:3888]};
      mid_0[1] = {1'b0,layer_2_0[3903:3896]} - {1'b0, layer_1_0[3903:3896]};
      mid_0[2] = {1'b0,layer_2_0[3911:3904]} - {1'b0, layer_1_0[3911:3904]};
      mid_1[0] = {1'b0,layer_2_1[3895:3888]} - {1'b0, layer_1_1[3895:3888]};
      mid_1[1] = {1'b0,layer_2_1[3903:3896]} - {1'b0, layer_1_1[3903:3896]};
      mid_1[2] = {1'b0,layer_2_1[3911:3904]} - {1'b0, layer_1_1[3911:3904]};
      mid_2[0] = {1'b0,layer_2_2[3895:3888]} - {1'b0, layer_1_2[3895:3888]};
      mid_2[1] = {1'b0,layer_2_2[3903:3896]} - {1'b0, layer_1_2[3903:3896]};
      mid_2[2] = {1'b0,layer_2_2[3911:3904]} - {1'b0, layer_1_2[3911:3904]};
      btm_0[0] = {1'b0,layer_3_0[3895:3888]} - {1'b0, layer_2_0[3895:3888]};
      btm_0[1] = {1'b0,layer_3_0[3903:3896]} - {1'b0, layer_2_0[3903:3896]};
      btm_0[2] = {1'b0,layer_3_0[3911:3904]} - {1'b0, layer_2_0[3911:3904]};
      btm_1[0] = {1'b0,layer_3_1[3895:3888]} - {1'b0, layer_2_1[3895:3888]};
      btm_1[1] = {1'b0,layer_3_1[3903:3896]} - {1'b0, layer_2_1[3903:3896]};
      btm_1[2] = {1'b0,layer_3_1[3911:3904]} - {1'b0, layer_2_1[3911:3904]};
      btm_2[0] = {1'b0,layer_3_2[3895:3888]} - {1'b0, layer_2_2[3895:3888]};
      btm_2[1] = {1'b0,layer_3_2[3903:3896]} - {1'b0, layer_2_2[3903:3896]};
      btm_2[2] = {1'b0,layer_3_2[3911:3904]} - {1'b0, layer_2_2[3911:3904]};
    end
    'd488: begin
      top_0[0] = {1'b0,layer_1_0[3903:3896]} - {1'b0, layer_0_0[3903:3896]};
      top_0[1] = {1'b0,layer_1_0[3911:3904]} - {1'b0, layer_0_0[3911:3904]};
      top_0[2] = {1'b0,layer_1_0[3919:3912]} - {1'b0, layer_0_0[3919:3912]};
      top_1[0] = {1'b0,layer_1_1[3903:3896]} - {1'b0, layer_0_1[3903:3896]};
      top_1[1] = {1'b0,layer_1_1[3911:3904]} - {1'b0, layer_0_1[3911:3904]};
      top_1[2] = {1'b0,layer_1_1[3919:3912]} - {1'b0, layer_0_1[3919:3912]};
      top_2[0] = {1'b0,layer_1_2[3903:3896]} - {1'b0, layer_0_2[3903:3896]};
      top_2[1] = {1'b0,layer_1_2[3911:3904]} - {1'b0, layer_0_2[3911:3904]};
      top_2[2] = {1'b0,layer_1_2[3919:3912]} - {1'b0, layer_0_2[3919:3912]};
      mid_0[0] = {1'b0,layer_2_0[3903:3896]} - {1'b0, layer_1_0[3903:3896]};
      mid_0[1] = {1'b0,layer_2_0[3911:3904]} - {1'b0, layer_1_0[3911:3904]};
      mid_0[2] = {1'b0,layer_2_0[3919:3912]} - {1'b0, layer_1_0[3919:3912]};
      mid_1[0] = {1'b0,layer_2_1[3903:3896]} - {1'b0, layer_1_1[3903:3896]};
      mid_1[1] = {1'b0,layer_2_1[3911:3904]} - {1'b0, layer_1_1[3911:3904]};
      mid_1[2] = {1'b0,layer_2_1[3919:3912]} - {1'b0, layer_1_1[3919:3912]};
      mid_2[0] = {1'b0,layer_2_2[3903:3896]} - {1'b0, layer_1_2[3903:3896]};
      mid_2[1] = {1'b0,layer_2_2[3911:3904]} - {1'b0, layer_1_2[3911:3904]};
      mid_2[2] = {1'b0,layer_2_2[3919:3912]} - {1'b0, layer_1_2[3919:3912]};
      btm_0[0] = {1'b0,layer_3_0[3903:3896]} - {1'b0, layer_2_0[3903:3896]};
      btm_0[1] = {1'b0,layer_3_0[3911:3904]} - {1'b0, layer_2_0[3911:3904]};
      btm_0[2] = {1'b0,layer_3_0[3919:3912]} - {1'b0, layer_2_0[3919:3912]};
      btm_1[0] = {1'b0,layer_3_1[3903:3896]} - {1'b0, layer_2_1[3903:3896]};
      btm_1[1] = {1'b0,layer_3_1[3911:3904]} - {1'b0, layer_2_1[3911:3904]};
      btm_1[2] = {1'b0,layer_3_1[3919:3912]} - {1'b0, layer_2_1[3919:3912]};
      btm_2[0] = {1'b0,layer_3_2[3903:3896]} - {1'b0, layer_2_2[3903:3896]};
      btm_2[1] = {1'b0,layer_3_2[3911:3904]} - {1'b0, layer_2_2[3911:3904]};
      btm_2[2] = {1'b0,layer_3_2[3919:3912]} - {1'b0, layer_2_2[3919:3912]};
    end
    'd489: begin
      top_0[0] = {1'b0,layer_1_0[3911:3904]} - {1'b0, layer_0_0[3911:3904]};
      top_0[1] = {1'b0,layer_1_0[3919:3912]} - {1'b0, layer_0_0[3919:3912]};
      top_0[2] = {1'b0,layer_1_0[3927:3920]} - {1'b0, layer_0_0[3927:3920]};
      top_1[0] = {1'b0,layer_1_1[3911:3904]} - {1'b0, layer_0_1[3911:3904]};
      top_1[1] = {1'b0,layer_1_1[3919:3912]} - {1'b0, layer_0_1[3919:3912]};
      top_1[2] = {1'b0,layer_1_1[3927:3920]} - {1'b0, layer_0_1[3927:3920]};
      top_2[0] = {1'b0,layer_1_2[3911:3904]} - {1'b0, layer_0_2[3911:3904]};
      top_2[1] = {1'b0,layer_1_2[3919:3912]} - {1'b0, layer_0_2[3919:3912]};
      top_2[2] = {1'b0,layer_1_2[3927:3920]} - {1'b0, layer_0_2[3927:3920]};
      mid_0[0] = {1'b0,layer_2_0[3911:3904]} - {1'b0, layer_1_0[3911:3904]};
      mid_0[1] = {1'b0,layer_2_0[3919:3912]} - {1'b0, layer_1_0[3919:3912]};
      mid_0[2] = {1'b0,layer_2_0[3927:3920]} - {1'b0, layer_1_0[3927:3920]};
      mid_1[0] = {1'b0,layer_2_1[3911:3904]} - {1'b0, layer_1_1[3911:3904]};
      mid_1[1] = {1'b0,layer_2_1[3919:3912]} - {1'b0, layer_1_1[3919:3912]};
      mid_1[2] = {1'b0,layer_2_1[3927:3920]} - {1'b0, layer_1_1[3927:3920]};
      mid_2[0] = {1'b0,layer_2_2[3911:3904]} - {1'b0, layer_1_2[3911:3904]};
      mid_2[1] = {1'b0,layer_2_2[3919:3912]} - {1'b0, layer_1_2[3919:3912]};
      mid_2[2] = {1'b0,layer_2_2[3927:3920]} - {1'b0, layer_1_2[3927:3920]};
      btm_0[0] = {1'b0,layer_3_0[3911:3904]} - {1'b0, layer_2_0[3911:3904]};
      btm_0[1] = {1'b0,layer_3_0[3919:3912]} - {1'b0, layer_2_0[3919:3912]};
      btm_0[2] = {1'b0,layer_3_0[3927:3920]} - {1'b0, layer_2_0[3927:3920]};
      btm_1[0] = {1'b0,layer_3_1[3911:3904]} - {1'b0, layer_2_1[3911:3904]};
      btm_1[1] = {1'b0,layer_3_1[3919:3912]} - {1'b0, layer_2_1[3919:3912]};
      btm_1[2] = {1'b0,layer_3_1[3927:3920]} - {1'b0, layer_2_1[3927:3920]};
      btm_2[0] = {1'b0,layer_3_2[3911:3904]} - {1'b0, layer_2_2[3911:3904]};
      btm_2[1] = {1'b0,layer_3_2[3919:3912]} - {1'b0, layer_2_2[3919:3912]};
      btm_2[2] = {1'b0,layer_3_2[3927:3920]} - {1'b0, layer_2_2[3927:3920]};
    end
    'd490: begin
      top_0[0] = {1'b0,layer_1_0[3919:3912]} - {1'b0, layer_0_0[3919:3912]};
      top_0[1] = {1'b0,layer_1_0[3927:3920]} - {1'b0, layer_0_0[3927:3920]};
      top_0[2] = {1'b0,layer_1_0[3935:3928]} - {1'b0, layer_0_0[3935:3928]};
      top_1[0] = {1'b0,layer_1_1[3919:3912]} - {1'b0, layer_0_1[3919:3912]};
      top_1[1] = {1'b0,layer_1_1[3927:3920]} - {1'b0, layer_0_1[3927:3920]};
      top_1[2] = {1'b0,layer_1_1[3935:3928]} - {1'b0, layer_0_1[3935:3928]};
      top_2[0] = {1'b0,layer_1_2[3919:3912]} - {1'b0, layer_0_2[3919:3912]};
      top_2[1] = {1'b0,layer_1_2[3927:3920]} - {1'b0, layer_0_2[3927:3920]};
      top_2[2] = {1'b0,layer_1_2[3935:3928]} - {1'b0, layer_0_2[3935:3928]};
      mid_0[0] = {1'b0,layer_2_0[3919:3912]} - {1'b0, layer_1_0[3919:3912]};
      mid_0[1] = {1'b0,layer_2_0[3927:3920]} - {1'b0, layer_1_0[3927:3920]};
      mid_0[2] = {1'b0,layer_2_0[3935:3928]} - {1'b0, layer_1_0[3935:3928]};
      mid_1[0] = {1'b0,layer_2_1[3919:3912]} - {1'b0, layer_1_1[3919:3912]};
      mid_1[1] = {1'b0,layer_2_1[3927:3920]} - {1'b0, layer_1_1[3927:3920]};
      mid_1[2] = {1'b0,layer_2_1[3935:3928]} - {1'b0, layer_1_1[3935:3928]};
      mid_2[0] = {1'b0,layer_2_2[3919:3912]} - {1'b0, layer_1_2[3919:3912]};
      mid_2[1] = {1'b0,layer_2_2[3927:3920]} - {1'b0, layer_1_2[3927:3920]};
      mid_2[2] = {1'b0,layer_2_2[3935:3928]} - {1'b0, layer_1_2[3935:3928]};
      btm_0[0] = {1'b0,layer_3_0[3919:3912]} - {1'b0, layer_2_0[3919:3912]};
      btm_0[1] = {1'b0,layer_3_0[3927:3920]} - {1'b0, layer_2_0[3927:3920]};
      btm_0[2] = {1'b0,layer_3_0[3935:3928]} - {1'b0, layer_2_0[3935:3928]};
      btm_1[0] = {1'b0,layer_3_1[3919:3912]} - {1'b0, layer_2_1[3919:3912]};
      btm_1[1] = {1'b0,layer_3_1[3927:3920]} - {1'b0, layer_2_1[3927:3920]};
      btm_1[2] = {1'b0,layer_3_1[3935:3928]} - {1'b0, layer_2_1[3935:3928]};
      btm_2[0] = {1'b0,layer_3_2[3919:3912]} - {1'b0, layer_2_2[3919:3912]};
      btm_2[1] = {1'b0,layer_3_2[3927:3920]} - {1'b0, layer_2_2[3927:3920]};
      btm_2[2] = {1'b0,layer_3_2[3935:3928]} - {1'b0, layer_2_2[3935:3928]};
    end
    'd491: begin
      top_0[0] = {1'b0,layer_1_0[3927:3920]} - {1'b0, layer_0_0[3927:3920]};
      top_0[1] = {1'b0,layer_1_0[3935:3928]} - {1'b0, layer_0_0[3935:3928]};
      top_0[2] = {1'b0,layer_1_0[3943:3936]} - {1'b0, layer_0_0[3943:3936]};
      top_1[0] = {1'b0,layer_1_1[3927:3920]} - {1'b0, layer_0_1[3927:3920]};
      top_1[1] = {1'b0,layer_1_1[3935:3928]} - {1'b0, layer_0_1[3935:3928]};
      top_1[2] = {1'b0,layer_1_1[3943:3936]} - {1'b0, layer_0_1[3943:3936]};
      top_2[0] = {1'b0,layer_1_2[3927:3920]} - {1'b0, layer_0_2[3927:3920]};
      top_2[1] = {1'b0,layer_1_2[3935:3928]} - {1'b0, layer_0_2[3935:3928]};
      top_2[2] = {1'b0,layer_1_2[3943:3936]} - {1'b0, layer_0_2[3943:3936]};
      mid_0[0] = {1'b0,layer_2_0[3927:3920]} - {1'b0, layer_1_0[3927:3920]};
      mid_0[1] = {1'b0,layer_2_0[3935:3928]} - {1'b0, layer_1_0[3935:3928]};
      mid_0[2] = {1'b0,layer_2_0[3943:3936]} - {1'b0, layer_1_0[3943:3936]};
      mid_1[0] = {1'b0,layer_2_1[3927:3920]} - {1'b0, layer_1_1[3927:3920]};
      mid_1[1] = {1'b0,layer_2_1[3935:3928]} - {1'b0, layer_1_1[3935:3928]};
      mid_1[2] = {1'b0,layer_2_1[3943:3936]} - {1'b0, layer_1_1[3943:3936]};
      mid_2[0] = {1'b0,layer_2_2[3927:3920]} - {1'b0, layer_1_2[3927:3920]};
      mid_2[1] = {1'b0,layer_2_2[3935:3928]} - {1'b0, layer_1_2[3935:3928]};
      mid_2[2] = {1'b0,layer_2_2[3943:3936]} - {1'b0, layer_1_2[3943:3936]};
      btm_0[0] = {1'b0,layer_3_0[3927:3920]} - {1'b0, layer_2_0[3927:3920]};
      btm_0[1] = {1'b0,layer_3_0[3935:3928]} - {1'b0, layer_2_0[3935:3928]};
      btm_0[2] = {1'b0,layer_3_0[3943:3936]} - {1'b0, layer_2_0[3943:3936]};
      btm_1[0] = {1'b0,layer_3_1[3927:3920]} - {1'b0, layer_2_1[3927:3920]};
      btm_1[1] = {1'b0,layer_3_1[3935:3928]} - {1'b0, layer_2_1[3935:3928]};
      btm_1[2] = {1'b0,layer_3_1[3943:3936]} - {1'b0, layer_2_1[3943:3936]};
      btm_2[0] = {1'b0,layer_3_2[3927:3920]} - {1'b0, layer_2_2[3927:3920]};
      btm_2[1] = {1'b0,layer_3_2[3935:3928]} - {1'b0, layer_2_2[3935:3928]};
      btm_2[2] = {1'b0,layer_3_2[3943:3936]} - {1'b0, layer_2_2[3943:3936]};
    end
    'd492: begin
      top_0[0] = {1'b0,layer_1_0[3935:3928]} - {1'b0, layer_0_0[3935:3928]};
      top_0[1] = {1'b0,layer_1_0[3943:3936]} - {1'b0, layer_0_0[3943:3936]};
      top_0[2] = {1'b0,layer_1_0[3951:3944]} - {1'b0, layer_0_0[3951:3944]};
      top_1[0] = {1'b0,layer_1_1[3935:3928]} - {1'b0, layer_0_1[3935:3928]};
      top_1[1] = {1'b0,layer_1_1[3943:3936]} - {1'b0, layer_0_1[3943:3936]};
      top_1[2] = {1'b0,layer_1_1[3951:3944]} - {1'b0, layer_0_1[3951:3944]};
      top_2[0] = {1'b0,layer_1_2[3935:3928]} - {1'b0, layer_0_2[3935:3928]};
      top_2[1] = {1'b0,layer_1_2[3943:3936]} - {1'b0, layer_0_2[3943:3936]};
      top_2[2] = {1'b0,layer_1_2[3951:3944]} - {1'b0, layer_0_2[3951:3944]};
      mid_0[0] = {1'b0,layer_2_0[3935:3928]} - {1'b0, layer_1_0[3935:3928]};
      mid_0[1] = {1'b0,layer_2_0[3943:3936]} - {1'b0, layer_1_0[3943:3936]};
      mid_0[2] = {1'b0,layer_2_0[3951:3944]} - {1'b0, layer_1_0[3951:3944]};
      mid_1[0] = {1'b0,layer_2_1[3935:3928]} - {1'b0, layer_1_1[3935:3928]};
      mid_1[1] = {1'b0,layer_2_1[3943:3936]} - {1'b0, layer_1_1[3943:3936]};
      mid_1[2] = {1'b0,layer_2_1[3951:3944]} - {1'b0, layer_1_1[3951:3944]};
      mid_2[0] = {1'b0,layer_2_2[3935:3928]} - {1'b0, layer_1_2[3935:3928]};
      mid_2[1] = {1'b0,layer_2_2[3943:3936]} - {1'b0, layer_1_2[3943:3936]};
      mid_2[2] = {1'b0,layer_2_2[3951:3944]} - {1'b0, layer_1_2[3951:3944]};
      btm_0[0] = {1'b0,layer_3_0[3935:3928]} - {1'b0, layer_2_0[3935:3928]};
      btm_0[1] = {1'b0,layer_3_0[3943:3936]} - {1'b0, layer_2_0[3943:3936]};
      btm_0[2] = {1'b0,layer_3_0[3951:3944]} - {1'b0, layer_2_0[3951:3944]};
      btm_1[0] = {1'b0,layer_3_1[3935:3928]} - {1'b0, layer_2_1[3935:3928]};
      btm_1[1] = {1'b0,layer_3_1[3943:3936]} - {1'b0, layer_2_1[3943:3936]};
      btm_1[2] = {1'b0,layer_3_1[3951:3944]} - {1'b0, layer_2_1[3951:3944]};
      btm_2[0] = {1'b0,layer_3_2[3935:3928]} - {1'b0, layer_2_2[3935:3928]};
      btm_2[1] = {1'b0,layer_3_2[3943:3936]} - {1'b0, layer_2_2[3943:3936]};
      btm_2[2] = {1'b0,layer_3_2[3951:3944]} - {1'b0, layer_2_2[3951:3944]};
    end
    'd493: begin
      top_0[0] = {1'b0,layer_1_0[3943:3936]} - {1'b0, layer_0_0[3943:3936]};
      top_0[1] = {1'b0,layer_1_0[3951:3944]} - {1'b0, layer_0_0[3951:3944]};
      top_0[2] = {1'b0,layer_1_0[3959:3952]} - {1'b0, layer_0_0[3959:3952]};
      top_1[0] = {1'b0,layer_1_1[3943:3936]} - {1'b0, layer_0_1[3943:3936]};
      top_1[1] = {1'b0,layer_1_1[3951:3944]} - {1'b0, layer_0_1[3951:3944]};
      top_1[2] = {1'b0,layer_1_1[3959:3952]} - {1'b0, layer_0_1[3959:3952]};
      top_2[0] = {1'b0,layer_1_2[3943:3936]} - {1'b0, layer_0_2[3943:3936]};
      top_2[1] = {1'b0,layer_1_2[3951:3944]} - {1'b0, layer_0_2[3951:3944]};
      top_2[2] = {1'b0,layer_1_2[3959:3952]} - {1'b0, layer_0_2[3959:3952]};
      mid_0[0] = {1'b0,layer_2_0[3943:3936]} - {1'b0, layer_1_0[3943:3936]};
      mid_0[1] = {1'b0,layer_2_0[3951:3944]} - {1'b0, layer_1_0[3951:3944]};
      mid_0[2] = {1'b0,layer_2_0[3959:3952]} - {1'b0, layer_1_0[3959:3952]};
      mid_1[0] = {1'b0,layer_2_1[3943:3936]} - {1'b0, layer_1_1[3943:3936]};
      mid_1[1] = {1'b0,layer_2_1[3951:3944]} - {1'b0, layer_1_1[3951:3944]};
      mid_1[2] = {1'b0,layer_2_1[3959:3952]} - {1'b0, layer_1_1[3959:3952]};
      mid_2[0] = {1'b0,layer_2_2[3943:3936]} - {1'b0, layer_1_2[3943:3936]};
      mid_2[1] = {1'b0,layer_2_2[3951:3944]} - {1'b0, layer_1_2[3951:3944]};
      mid_2[2] = {1'b0,layer_2_2[3959:3952]} - {1'b0, layer_1_2[3959:3952]};
      btm_0[0] = {1'b0,layer_3_0[3943:3936]} - {1'b0, layer_2_0[3943:3936]};
      btm_0[1] = {1'b0,layer_3_0[3951:3944]} - {1'b0, layer_2_0[3951:3944]};
      btm_0[2] = {1'b0,layer_3_0[3959:3952]} - {1'b0, layer_2_0[3959:3952]};
      btm_1[0] = {1'b0,layer_3_1[3943:3936]} - {1'b0, layer_2_1[3943:3936]};
      btm_1[1] = {1'b0,layer_3_1[3951:3944]} - {1'b0, layer_2_1[3951:3944]};
      btm_1[2] = {1'b0,layer_3_1[3959:3952]} - {1'b0, layer_2_1[3959:3952]};
      btm_2[0] = {1'b0,layer_3_2[3943:3936]} - {1'b0, layer_2_2[3943:3936]};
      btm_2[1] = {1'b0,layer_3_2[3951:3944]} - {1'b0, layer_2_2[3951:3944]};
      btm_2[2] = {1'b0,layer_3_2[3959:3952]} - {1'b0, layer_2_2[3959:3952]};
    end
    'd494: begin
      top_0[0] = {1'b0,layer_1_0[3951:3944]} - {1'b0, layer_0_0[3951:3944]};
      top_0[1] = {1'b0,layer_1_0[3959:3952]} - {1'b0, layer_0_0[3959:3952]};
      top_0[2] = {1'b0,layer_1_0[3967:3960]} - {1'b0, layer_0_0[3967:3960]};
      top_1[0] = {1'b0,layer_1_1[3951:3944]} - {1'b0, layer_0_1[3951:3944]};
      top_1[1] = {1'b0,layer_1_1[3959:3952]} - {1'b0, layer_0_1[3959:3952]};
      top_1[2] = {1'b0,layer_1_1[3967:3960]} - {1'b0, layer_0_1[3967:3960]};
      top_2[0] = {1'b0,layer_1_2[3951:3944]} - {1'b0, layer_0_2[3951:3944]};
      top_2[1] = {1'b0,layer_1_2[3959:3952]} - {1'b0, layer_0_2[3959:3952]};
      top_2[2] = {1'b0,layer_1_2[3967:3960]} - {1'b0, layer_0_2[3967:3960]};
      mid_0[0] = {1'b0,layer_2_0[3951:3944]} - {1'b0, layer_1_0[3951:3944]};
      mid_0[1] = {1'b0,layer_2_0[3959:3952]} - {1'b0, layer_1_0[3959:3952]};
      mid_0[2] = {1'b0,layer_2_0[3967:3960]} - {1'b0, layer_1_0[3967:3960]};
      mid_1[0] = {1'b0,layer_2_1[3951:3944]} - {1'b0, layer_1_1[3951:3944]};
      mid_1[1] = {1'b0,layer_2_1[3959:3952]} - {1'b0, layer_1_1[3959:3952]};
      mid_1[2] = {1'b0,layer_2_1[3967:3960]} - {1'b0, layer_1_1[3967:3960]};
      mid_2[0] = {1'b0,layer_2_2[3951:3944]} - {1'b0, layer_1_2[3951:3944]};
      mid_2[1] = {1'b0,layer_2_2[3959:3952]} - {1'b0, layer_1_2[3959:3952]};
      mid_2[2] = {1'b0,layer_2_2[3967:3960]} - {1'b0, layer_1_2[3967:3960]};
      btm_0[0] = {1'b0,layer_3_0[3951:3944]} - {1'b0, layer_2_0[3951:3944]};
      btm_0[1] = {1'b0,layer_3_0[3959:3952]} - {1'b0, layer_2_0[3959:3952]};
      btm_0[2] = {1'b0,layer_3_0[3967:3960]} - {1'b0, layer_2_0[3967:3960]};
      btm_1[0] = {1'b0,layer_3_1[3951:3944]} - {1'b0, layer_2_1[3951:3944]};
      btm_1[1] = {1'b0,layer_3_1[3959:3952]} - {1'b0, layer_2_1[3959:3952]};
      btm_1[2] = {1'b0,layer_3_1[3967:3960]} - {1'b0, layer_2_1[3967:3960]};
      btm_2[0] = {1'b0,layer_3_2[3951:3944]} - {1'b0, layer_2_2[3951:3944]};
      btm_2[1] = {1'b0,layer_3_2[3959:3952]} - {1'b0, layer_2_2[3959:3952]};
      btm_2[2] = {1'b0,layer_3_2[3967:3960]} - {1'b0, layer_2_2[3967:3960]};
    end
    'd495: begin
      top_0[0] = {1'b0,layer_1_0[3959:3952]} - {1'b0, layer_0_0[3959:3952]};
      top_0[1] = {1'b0,layer_1_0[3967:3960]} - {1'b0, layer_0_0[3967:3960]};
      top_0[2] = {1'b0,layer_1_0[3975:3968]} - {1'b0, layer_0_0[3975:3968]};
      top_1[0] = {1'b0,layer_1_1[3959:3952]} - {1'b0, layer_0_1[3959:3952]};
      top_1[1] = {1'b0,layer_1_1[3967:3960]} - {1'b0, layer_0_1[3967:3960]};
      top_1[2] = {1'b0,layer_1_1[3975:3968]} - {1'b0, layer_0_1[3975:3968]};
      top_2[0] = {1'b0,layer_1_2[3959:3952]} - {1'b0, layer_0_2[3959:3952]};
      top_2[1] = {1'b0,layer_1_2[3967:3960]} - {1'b0, layer_0_2[3967:3960]};
      top_2[2] = {1'b0,layer_1_2[3975:3968]} - {1'b0, layer_0_2[3975:3968]};
      mid_0[0] = {1'b0,layer_2_0[3959:3952]} - {1'b0, layer_1_0[3959:3952]};
      mid_0[1] = {1'b0,layer_2_0[3967:3960]} - {1'b0, layer_1_0[3967:3960]};
      mid_0[2] = {1'b0,layer_2_0[3975:3968]} - {1'b0, layer_1_0[3975:3968]};
      mid_1[0] = {1'b0,layer_2_1[3959:3952]} - {1'b0, layer_1_1[3959:3952]};
      mid_1[1] = {1'b0,layer_2_1[3967:3960]} - {1'b0, layer_1_1[3967:3960]};
      mid_1[2] = {1'b0,layer_2_1[3975:3968]} - {1'b0, layer_1_1[3975:3968]};
      mid_2[0] = {1'b0,layer_2_2[3959:3952]} - {1'b0, layer_1_2[3959:3952]};
      mid_2[1] = {1'b0,layer_2_2[3967:3960]} - {1'b0, layer_1_2[3967:3960]};
      mid_2[2] = {1'b0,layer_2_2[3975:3968]} - {1'b0, layer_1_2[3975:3968]};
      btm_0[0] = {1'b0,layer_3_0[3959:3952]} - {1'b0, layer_2_0[3959:3952]};
      btm_0[1] = {1'b0,layer_3_0[3967:3960]} - {1'b0, layer_2_0[3967:3960]};
      btm_0[2] = {1'b0,layer_3_0[3975:3968]} - {1'b0, layer_2_0[3975:3968]};
      btm_1[0] = {1'b0,layer_3_1[3959:3952]} - {1'b0, layer_2_1[3959:3952]};
      btm_1[1] = {1'b0,layer_3_1[3967:3960]} - {1'b0, layer_2_1[3967:3960]};
      btm_1[2] = {1'b0,layer_3_1[3975:3968]} - {1'b0, layer_2_1[3975:3968]};
      btm_2[0] = {1'b0,layer_3_2[3959:3952]} - {1'b0, layer_2_2[3959:3952]};
      btm_2[1] = {1'b0,layer_3_2[3967:3960]} - {1'b0, layer_2_2[3967:3960]};
      btm_2[2] = {1'b0,layer_3_2[3975:3968]} - {1'b0, layer_2_2[3975:3968]};
    end
    'd496: begin
      top_0[0] = {1'b0,layer_1_0[3967:3960]} - {1'b0, layer_0_0[3967:3960]};
      top_0[1] = {1'b0,layer_1_0[3975:3968]} - {1'b0, layer_0_0[3975:3968]};
      top_0[2] = {1'b0,layer_1_0[3983:3976]} - {1'b0, layer_0_0[3983:3976]};
      top_1[0] = {1'b0,layer_1_1[3967:3960]} - {1'b0, layer_0_1[3967:3960]};
      top_1[1] = {1'b0,layer_1_1[3975:3968]} - {1'b0, layer_0_1[3975:3968]};
      top_1[2] = {1'b0,layer_1_1[3983:3976]} - {1'b0, layer_0_1[3983:3976]};
      top_2[0] = {1'b0,layer_1_2[3967:3960]} - {1'b0, layer_0_2[3967:3960]};
      top_2[1] = {1'b0,layer_1_2[3975:3968]} - {1'b0, layer_0_2[3975:3968]};
      top_2[2] = {1'b0,layer_1_2[3983:3976]} - {1'b0, layer_0_2[3983:3976]};
      mid_0[0] = {1'b0,layer_2_0[3967:3960]} - {1'b0, layer_1_0[3967:3960]};
      mid_0[1] = {1'b0,layer_2_0[3975:3968]} - {1'b0, layer_1_0[3975:3968]};
      mid_0[2] = {1'b0,layer_2_0[3983:3976]} - {1'b0, layer_1_0[3983:3976]};
      mid_1[0] = {1'b0,layer_2_1[3967:3960]} - {1'b0, layer_1_1[3967:3960]};
      mid_1[1] = {1'b0,layer_2_1[3975:3968]} - {1'b0, layer_1_1[3975:3968]};
      mid_1[2] = {1'b0,layer_2_1[3983:3976]} - {1'b0, layer_1_1[3983:3976]};
      mid_2[0] = {1'b0,layer_2_2[3967:3960]} - {1'b0, layer_1_2[3967:3960]};
      mid_2[1] = {1'b0,layer_2_2[3975:3968]} - {1'b0, layer_1_2[3975:3968]};
      mid_2[2] = {1'b0,layer_2_2[3983:3976]} - {1'b0, layer_1_2[3983:3976]};
      btm_0[0] = {1'b0,layer_3_0[3967:3960]} - {1'b0, layer_2_0[3967:3960]};
      btm_0[1] = {1'b0,layer_3_0[3975:3968]} - {1'b0, layer_2_0[3975:3968]};
      btm_0[2] = {1'b0,layer_3_0[3983:3976]} - {1'b0, layer_2_0[3983:3976]};
      btm_1[0] = {1'b0,layer_3_1[3967:3960]} - {1'b0, layer_2_1[3967:3960]};
      btm_1[1] = {1'b0,layer_3_1[3975:3968]} - {1'b0, layer_2_1[3975:3968]};
      btm_1[2] = {1'b0,layer_3_1[3983:3976]} - {1'b0, layer_2_1[3983:3976]};
      btm_2[0] = {1'b0,layer_3_2[3967:3960]} - {1'b0, layer_2_2[3967:3960]};
      btm_2[1] = {1'b0,layer_3_2[3975:3968]} - {1'b0, layer_2_2[3975:3968]};
      btm_2[2] = {1'b0,layer_3_2[3983:3976]} - {1'b0, layer_2_2[3983:3976]};
    end
    'd497: begin
      top_0[0] = {1'b0,layer_1_0[3975:3968]} - {1'b0, layer_0_0[3975:3968]};
      top_0[1] = {1'b0,layer_1_0[3983:3976]} - {1'b0, layer_0_0[3983:3976]};
      top_0[2] = {1'b0,layer_1_0[3991:3984]} - {1'b0, layer_0_0[3991:3984]};
      top_1[0] = {1'b0,layer_1_1[3975:3968]} - {1'b0, layer_0_1[3975:3968]};
      top_1[1] = {1'b0,layer_1_1[3983:3976]} - {1'b0, layer_0_1[3983:3976]};
      top_1[2] = {1'b0,layer_1_1[3991:3984]} - {1'b0, layer_0_1[3991:3984]};
      top_2[0] = {1'b0,layer_1_2[3975:3968]} - {1'b0, layer_0_2[3975:3968]};
      top_2[1] = {1'b0,layer_1_2[3983:3976]} - {1'b0, layer_0_2[3983:3976]};
      top_2[2] = {1'b0,layer_1_2[3991:3984]} - {1'b0, layer_0_2[3991:3984]};
      mid_0[0] = {1'b0,layer_2_0[3975:3968]} - {1'b0, layer_1_0[3975:3968]};
      mid_0[1] = {1'b0,layer_2_0[3983:3976]} - {1'b0, layer_1_0[3983:3976]};
      mid_0[2] = {1'b0,layer_2_0[3991:3984]} - {1'b0, layer_1_0[3991:3984]};
      mid_1[0] = {1'b0,layer_2_1[3975:3968]} - {1'b0, layer_1_1[3975:3968]};
      mid_1[1] = {1'b0,layer_2_1[3983:3976]} - {1'b0, layer_1_1[3983:3976]};
      mid_1[2] = {1'b0,layer_2_1[3991:3984]} - {1'b0, layer_1_1[3991:3984]};
      mid_2[0] = {1'b0,layer_2_2[3975:3968]} - {1'b0, layer_1_2[3975:3968]};
      mid_2[1] = {1'b0,layer_2_2[3983:3976]} - {1'b0, layer_1_2[3983:3976]};
      mid_2[2] = {1'b0,layer_2_2[3991:3984]} - {1'b0, layer_1_2[3991:3984]};
      btm_0[0] = {1'b0,layer_3_0[3975:3968]} - {1'b0, layer_2_0[3975:3968]};
      btm_0[1] = {1'b0,layer_3_0[3983:3976]} - {1'b0, layer_2_0[3983:3976]};
      btm_0[2] = {1'b0,layer_3_0[3991:3984]} - {1'b0, layer_2_0[3991:3984]};
      btm_1[0] = {1'b0,layer_3_1[3975:3968]} - {1'b0, layer_2_1[3975:3968]};
      btm_1[1] = {1'b0,layer_3_1[3983:3976]} - {1'b0, layer_2_1[3983:3976]};
      btm_1[2] = {1'b0,layer_3_1[3991:3984]} - {1'b0, layer_2_1[3991:3984]};
      btm_2[0] = {1'b0,layer_3_2[3975:3968]} - {1'b0, layer_2_2[3975:3968]};
      btm_2[1] = {1'b0,layer_3_2[3983:3976]} - {1'b0, layer_2_2[3983:3976]};
      btm_2[2] = {1'b0,layer_3_2[3991:3984]} - {1'b0, layer_2_2[3991:3984]};
    end
    'd498: begin
      top_0[0] = {1'b0,layer_1_0[3983:3976]} - {1'b0, layer_0_0[3983:3976]};
      top_0[1] = {1'b0,layer_1_0[3991:3984]} - {1'b0, layer_0_0[3991:3984]};
      top_0[2] = {1'b0,layer_1_0[3999:3992]} - {1'b0, layer_0_0[3999:3992]};
      top_1[0] = {1'b0,layer_1_1[3983:3976]} - {1'b0, layer_0_1[3983:3976]};
      top_1[1] = {1'b0,layer_1_1[3991:3984]} - {1'b0, layer_0_1[3991:3984]};
      top_1[2] = {1'b0,layer_1_1[3999:3992]} - {1'b0, layer_0_1[3999:3992]};
      top_2[0] = {1'b0,layer_1_2[3983:3976]} - {1'b0, layer_0_2[3983:3976]};
      top_2[1] = {1'b0,layer_1_2[3991:3984]} - {1'b0, layer_0_2[3991:3984]};
      top_2[2] = {1'b0,layer_1_2[3999:3992]} - {1'b0, layer_0_2[3999:3992]};
      mid_0[0] = {1'b0,layer_2_0[3983:3976]} - {1'b0, layer_1_0[3983:3976]};
      mid_0[1] = {1'b0,layer_2_0[3991:3984]} - {1'b0, layer_1_0[3991:3984]};
      mid_0[2] = {1'b0,layer_2_0[3999:3992]} - {1'b0, layer_1_0[3999:3992]};
      mid_1[0] = {1'b0,layer_2_1[3983:3976]} - {1'b0, layer_1_1[3983:3976]};
      mid_1[1] = {1'b0,layer_2_1[3991:3984]} - {1'b0, layer_1_1[3991:3984]};
      mid_1[2] = {1'b0,layer_2_1[3999:3992]} - {1'b0, layer_1_1[3999:3992]};
      mid_2[0] = {1'b0,layer_2_2[3983:3976]} - {1'b0, layer_1_2[3983:3976]};
      mid_2[1] = {1'b0,layer_2_2[3991:3984]} - {1'b0, layer_1_2[3991:3984]};
      mid_2[2] = {1'b0,layer_2_2[3999:3992]} - {1'b0, layer_1_2[3999:3992]};
      btm_0[0] = {1'b0,layer_3_0[3983:3976]} - {1'b0, layer_2_0[3983:3976]};
      btm_0[1] = {1'b0,layer_3_0[3991:3984]} - {1'b0, layer_2_0[3991:3984]};
      btm_0[2] = {1'b0,layer_3_0[3999:3992]} - {1'b0, layer_2_0[3999:3992]};
      btm_1[0] = {1'b0,layer_3_1[3983:3976]} - {1'b0, layer_2_1[3983:3976]};
      btm_1[1] = {1'b0,layer_3_1[3991:3984]} - {1'b0, layer_2_1[3991:3984]};
      btm_1[2] = {1'b0,layer_3_1[3999:3992]} - {1'b0, layer_2_1[3999:3992]};
      btm_2[0] = {1'b0,layer_3_2[3983:3976]} - {1'b0, layer_2_2[3983:3976]};
      btm_2[1] = {1'b0,layer_3_2[3991:3984]} - {1'b0, layer_2_2[3991:3984]};
      btm_2[2] = {1'b0,layer_3_2[3999:3992]} - {1'b0, layer_2_2[3999:3992]};
    end
    'd499: begin
      top_0[0] = {1'b0,layer_1_0[3991:3984]} - {1'b0, layer_0_0[3991:3984]};
      top_0[1] = {1'b0,layer_1_0[3999:3992]} - {1'b0, layer_0_0[3999:3992]};
      top_0[2] = {1'b0,layer_1_0[4007:4000]} - {1'b0, layer_0_0[4007:4000]};
      top_1[0] = {1'b0,layer_1_1[3991:3984]} - {1'b0, layer_0_1[3991:3984]};
      top_1[1] = {1'b0,layer_1_1[3999:3992]} - {1'b0, layer_0_1[3999:3992]};
      top_1[2] = {1'b0,layer_1_1[4007:4000]} - {1'b0, layer_0_1[4007:4000]};
      top_2[0] = {1'b0,layer_1_2[3991:3984]} - {1'b0, layer_0_2[3991:3984]};
      top_2[1] = {1'b0,layer_1_2[3999:3992]} - {1'b0, layer_0_2[3999:3992]};
      top_2[2] = {1'b0,layer_1_2[4007:4000]} - {1'b0, layer_0_2[4007:4000]};
      mid_0[0] = {1'b0,layer_2_0[3991:3984]} - {1'b0, layer_1_0[3991:3984]};
      mid_0[1] = {1'b0,layer_2_0[3999:3992]} - {1'b0, layer_1_0[3999:3992]};
      mid_0[2] = {1'b0,layer_2_0[4007:4000]} - {1'b0, layer_1_0[4007:4000]};
      mid_1[0] = {1'b0,layer_2_1[3991:3984]} - {1'b0, layer_1_1[3991:3984]};
      mid_1[1] = {1'b0,layer_2_1[3999:3992]} - {1'b0, layer_1_1[3999:3992]};
      mid_1[2] = {1'b0,layer_2_1[4007:4000]} - {1'b0, layer_1_1[4007:4000]};
      mid_2[0] = {1'b0,layer_2_2[3991:3984]} - {1'b0, layer_1_2[3991:3984]};
      mid_2[1] = {1'b0,layer_2_2[3999:3992]} - {1'b0, layer_1_2[3999:3992]};
      mid_2[2] = {1'b0,layer_2_2[4007:4000]} - {1'b0, layer_1_2[4007:4000]};
      btm_0[0] = {1'b0,layer_3_0[3991:3984]} - {1'b0, layer_2_0[3991:3984]};
      btm_0[1] = {1'b0,layer_3_0[3999:3992]} - {1'b0, layer_2_0[3999:3992]};
      btm_0[2] = {1'b0,layer_3_0[4007:4000]} - {1'b0, layer_2_0[4007:4000]};
      btm_1[0] = {1'b0,layer_3_1[3991:3984]} - {1'b0, layer_2_1[3991:3984]};
      btm_1[1] = {1'b0,layer_3_1[3999:3992]} - {1'b0, layer_2_1[3999:3992]};
      btm_1[2] = {1'b0,layer_3_1[4007:4000]} - {1'b0, layer_2_1[4007:4000]};
      btm_2[0] = {1'b0,layer_3_2[3991:3984]} - {1'b0, layer_2_2[3991:3984]};
      btm_2[1] = {1'b0,layer_3_2[3999:3992]} - {1'b0, layer_2_2[3999:3992]};
      btm_2[2] = {1'b0,layer_3_2[4007:4000]} - {1'b0, layer_2_2[4007:4000]};
    end
    'd500: begin
      top_0[0] = {1'b0,layer_1_0[3999:3992]} - {1'b0, layer_0_0[3999:3992]};
      top_0[1] = {1'b0,layer_1_0[4007:4000]} - {1'b0, layer_0_0[4007:4000]};
      top_0[2] = {1'b0,layer_1_0[4015:4008]} - {1'b0, layer_0_0[4015:4008]};
      top_1[0] = {1'b0,layer_1_1[3999:3992]} - {1'b0, layer_0_1[3999:3992]};
      top_1[1] = {1'b0,layer_1_1[4007:4000]} - {1'b0, layer_0_1[4007:4000]};
      top_1[2] = {1'b0,layer_1_1[4015:4008]} - {1'b0, layer_0_1[4015:4008]};
      top_2[0] = {1'b0,layer_1_2[3999:3992]} - {1'b0, layer_0_2[3999:3992]};
      top_2[1] = {1'b0,layer_1_2[4007:4000]} - {1'b0, layer_0_2[4007:4000]};
      top_2[2] = {1'b0,layer_1_2[4015:4008]} - {1'b0, layer_0_2[4015:4008]};
      mid_0[0] = {1'b0,layer_2_0[3999:3992]} - {1'b0, layer_1_0[3999:3992]};
      mid_0[1] = {1'b0,layer_2_0[4007:4000]} - {1'b0, layer_1_0[4007:4000]};
      mid_0[2] = {1'b0,layer_2_0[4015:4008]} - {1'b0, layer_1_0[4015:4008]};
      mid_1[0] = {1'b0,layer_2_1[3999:3992]} - {1'b0, layer_1_1[3999:3992]};
      mid_1[1] = {1'b0,layer_2_1[4007:4000]} - {1'b0, layer_1_1[4007:4000]};
      mid_1[2] = {1'b0,layer_2_1[4015:4008]} - {1'b0, layer_1_1[4015:4008]};
      mid_2[0] = {1'b0,layer_2_2[3999:3992]} - {1'b0, layer_1_2[3999:3992]};
      mid_2[1] = {1'b0,layer_2_2[4007:4000]} - {1'b0, layer_1_2[4007:4000]};
      mid_2[2] = {1'b0,layer_2_2[4015:4008]} - {1'b0, layer_1_2[4015:4008]};
      btm_0[0] = {1'b0,layer_3_0[3999:3992]} - {1'b0, layer_2_0[3999:3992]};
      btm_0[1] = {1'b0,layer_3_0[4007:4000]} - {1'b0, layer_2_0[4007:4000]};
      btm_0[2] = {1'b0,layer_3_0[4015:4008]} - {1'b0, layer_2_0[4015:4008]};
      btm_1[0] = {1'b0,layer_3_1[3999:3992]} - {1'b0, layer_2_1[3999:3992]};
      btm_1[1] = {1'b0,layer_3_1[4007:4000]} - {1'b0, layer_2_1[4007:4000]};
      btm_1[2] = {1'b0,layer_3_1[4015:4008]} - {1'b0, layer_2_1[4015:4008]};
      btm_2[0] = {1'b0,layer_3_2[3999:3992]} - {1'b0, layer_2_2[3999:3992]};
      btm_2[1] = {1'b0,layer_3_2[4007:4000]} - {1'b0, layer_2_2[4007:4000]};
      btm_2[2] = {1'b0,layer_3_2[4015:4008]} - {1'b0, layer_2_2[4015:4008]};
    end
    'd501: begin
      top_0[0] = {1'b0,layer_1_0[4007:4000]} - {1'b0, layer_0_0[4007:4000]};
      top_0[1] = {1'b0,layer_1_0[4015:4008]} - {1'b0, layer_0_0[4015:4008]};
      top_0[2] = {1'b0,layer_1_0[4023:4016]} - {1'b0, layer_0_0[4023:4016]};
      top_1[0] = {1'b0,layer_1_1[4007:4000]} - {1'b0, layer_0_1[4007:4000]};
      top_1[1] = {1'b0,layer_1_1[4015:4008]} - {1'b0, layer_0_1[4015:4008]};
      top_1[2] = {1'b0,layer_1_1[4023:4016]} - {1'b0, layer_0_1[4023:4016]};
      top_2[0] = {1'b0,layer_1_2[4007:4000]} - {1'b0, layer_0_2[4007:4000]};
      top_2[1] = {1'b0,layer_1_2[4015:4008]} - {1'b0, layer_0_2[4015:4008]};
      top_2[2] = {1'b0,layer_1_2[4023:4016]} - {1'b0, layer_0_2[4023:4016]};
      mid_0[0] = {1'b0,layer_2_0[4007:4000]} - {1'b0, layer_1_0[4007:4000]};
      mid_0[1] = {1'b0,layer_2_0[4015:4008]} - {1'b0, layer_1_0[4015:4008]};
      mid_0[2] = {1'b0,layer_2_0[4023:4016]} - {1'b0, layer_1_0[4023:4016]};
      mid_1[0] = {1'b0,layer_2_1[4007:4000]} - {1'b0, layer_1_1[4007:4000]};
      mid_1[1] = {1'b0,layer_2_1[4015:4008]} - {1'b0, layer_1_1[4015:4008]};
      mid_1[2] = {1'b0,layer_2_1[4023:4016]} - {1'b0, layer_1_1[4023:4016]};
      mid_2[0] = {1'b0,layer_2_2[4007:4000]} - {1'b0, layer_1_2[4007:4000]};
      mid_2[1] = {1'b0,layer_2_2[4015:4008]} - {1'b0, layer_1_2[4015:4008]};
      mid_2[2] = {1'b0,layer_2_2[4023:4016]} - {1'b0, layer_1_2[4023:4016]};
      btm_0[0] = {1'b0,layer_3_0[4007:4000]} - {1'b0, layer_2_0[4007:4000]};
      btm_0[1] = {1'b0,layer_3_0[4015:4008]} - {1'b0, layer_2_0[4015:4008]};
      btm_0[2] = {1'b0,layer_3_0[4023:4016]} - {1'b0, layer_2_0[4023:4016]};
      btm_1[0] = {1'b0,layer_3_1[4007:4000]} - {1'b0, layer_2_1[4007:4000]};
      btm_1[1] = {1'b0,layer_3_1[4015:4008]} - {1'b0, layer_2_1[4015:4008]};
      btm_1[2] = {1'b0,layer_3_1[4023:4016]} - {1'b0, layer_2_1[4023:4016]};
      btm_2[0] = {1'b0,layer_3_2[4007:4000]} - {1'b0, layer_2_2[4007:4000]};
      btm_2[1] = {1'b0,layer_3_2[4015:4008]} - {1'b0, layer_2_2[4015:4008]};
      btm_2[2] = {1'b0,layer_3_2[4023:4016]} - {1'b0, layer_2_2[4023:4016]};
    end
    'd502: begin
      top_0[0] = {1'b0,layer_1_0[4015:4008]} - {1'b0, layer_0_0[4015:4008]};
      top_0[1] = {1'b0,layer_1_0[4023:4016]} - {1'b0, layer_0_0[4023:4016]};
      top_0[2] = {1'b0,layer_1_0[4031:4024]} - {1'b0, layer_0_0[4031:4024]};
      top_1[0] = {1'b0,layer_1_1[4015:4008]} - {1'b0, layer_0_1[4015:4008]};
      top_1[1] = {1'b0,layer_1_1[4023:4016]} - {1'b0, layer_0_1[4023:4016]};
      top_1[2] = {1'b0,layer_1_1[4031:4024]} - {1'b0, layer_0_1[4031:4024]};
      top_2[0] = {1'b0,layer_1_2[4015:4008]} - {1'b0, layer_0_2[4015:4008]};
      top_2[1] = {1'b0,layer_1_2[4023:4016]} - {1'b0, layer_0_2[4023:4016]};
      top_2[2] = {1'b0,layer_1_2[4031:4024]} - {1'b0, layer_0_2[4031:4024]};
      mid_0[0] = {1'b0,layer_2_0[4015:4008]} - {1'b0, layer_1_0[4015:4008]};
      mid_0[1] = {1'b0,layer_2_0[4023:4016]} - {1'b0, layer_1_0[4023:4016]};
      mid_0[2] = {1'b0,layer_2_0[4031:4024]} - {1'b0, layer_1_0[4031:4024]};
      mid_1[0] = {1'b0,layer_2_1[4015:4008]} - {1'b0, layer_1_1[4015:4008]};
      mid_1[1] = {1'b0,layer_2_1[4023:4016]} - {1'b0, layer_1_1[4023:4016]};
      mid_1[2] = {1'b0,layer_2_1[4031:4024]} - {1'b0, layer_1_1[4031:4024]};
      mid_2[0] = {1'b0,layer_2_2[4015:4008]} - {1'b0, layer_1_2[4015:4008]};
      mid_2[1] = {1'b0,layer_2_2[4023:4016]} - {1'b0, layer_1_2[4023:4016]};
      mid_2[2] = {1'b0,layer_2_2[4031:4024]} - {1'b0, layer_1_2[4031:4024]};
      btm_0[0] = {1'b0,layer_3_0[4015:4008]} - {1'b0, layer_2_0[4015:4008]};
      btm_0[1] = {1'b0,layer_3_0[4023:4016]} - {1'b0, layer_2_0[4023:4016]};
      btm_0[2] = {1'b0,layer_3_0[4031:4024]} - {1'b0, layer_2_0[4031:4024]};
      btm_1[0] = {1'b0,layer_3_1[4015:4008]} - {1'b0, layer_2_1[4015:4008]};
      btm_1[1] = {1'b0,layer_3_1[4023:4016]} - {1'b0, layer_2_1[4023:4016]};
      btm_1[2] = {1'b0,layer_3_1[4031:4024]} - {1'b0, layer_2_1[4031:4024]};
      btm_2[0] = {1'b0,layer_3_2[4015:4008]} - {1'b0, layer_2_2[4015:4008]};
      btm_2[1] = {1'b0,layer_3_2[4023:4016]} - {1'b0, layer_2_2[4023:4016]};
      btm_2[2] = {1'b0,layer_3_2[4031:4024]} - {1'b0, layer_2_2[4031:4024]};
    end
    'd503: begin
      top_0[0] = {1'b0,layer_1_0[4023:4016]} - {1'b0, layer_0_0[4023:4016]};
      top_0[1] = {1'b0,layer_1_0[4031:4024]} - {1'b0, layer_0_0[4031:4024]};
      top_0[2] = {1'b0,layer_1_0[4039:4032]} - {1'b0, layer_0_0[4039:4032]};
      top_1[0] = {1'b0,layer_1_1[4023:4016]} - {1'b0, layer_0_1[4023:4016]};
      top_1[1] = {1'b0,layer_1_1[4031:4024]} - {1'b0, layer_0_1[4031:4024]};
      top_1[2] = {1'b0,layer_1_1[4039:4032]} - {1'b0, layer_0_1[4039:4032]};
      top_2[0] = {1'b0,layer_1_2[4023:4016]} - {1'b0, layer_0_2[4023:4016]};
      top_2[1] = {1'b0,layer_1_2[4031:4024]} - {1'b0, layer_0_2[4031:4024]};
      top_2[2] = {1'b0,layer_1_2[4039:4032]} - {1'b0, layer_0_2[4039:4032]};
      mid_0[0] = {1'b0,layer_2_0[4023:4016]} - {1'b0, layer_1_0[4023:4016]};
      mid_0[1] = {1'b0,layer_2_0[4031:4024]} - {1'b0, layer_1_0[4031:4024]};
      mid_0[2] = {1'b0,layer_2_0[4039:4032]} - {1'b0, layer_1_0[4039:4032]};
      mid_1[0] = {1'b0,layer_2_1[4023:4016]} - {1'b0, layer_1_1[4023:4016]};
      mid_1[1] = {1'b0,layer_2_1[4031:4024]} - {1'b0, layer_1_1[4031:4024]};
      mid_1[2] = {1'b0,layer_2_1[4039:4032]} - {1'b0, layer_1_1[4039:4032]};
      mid_2[0] = {1'b0,layer_2_2[4023:4016]} - {1'b0, layer_1_2[4023:4016]};
      mid_2[1] = {1'b0,layer_2_2[4031:4024]} - {1'b0, layer_1_2[4031:4024]};
      mid_2[2] = {1'b0,layer_2_2[4039:4032]} - {1'b0, layer_1_2[4039:4032]};
      btm_0[0] = {1'b0,layer_3_0[4023:4016]} - {1'b0, layer_2_0[4023:4016]};
      btm_0[1] = {1'b0,layer_3_0[4031:4024]} - {1'b0, layer_2_0[4031:4024]};
      btm_0[2] = {1'b0,layer_3_0[4039:4032]} - {1'b0, layer_2_0[4039:4032]};
      btm_1[0] = {1'b0,layer_3_1[4023:4016]} - {1'b0, layer_2_1[4023:4016]};
      btm_1[1] = {1'b0,layer_3_1[4031:4024]} - {1'b0, layer_2_1[4031:4024]};
      btm_1[2] = {1'b0,layer_3_1[4039:4032]} - {1'b0, layer_2_1[4039:4032]};
      btm_2[0] = {1'b0,layer_3_2[4023:4016]} - {1'b0, layer_2_2[4023:4016]};
      btm_2[1] = {1'b0,layer_3_2[4031:4024]} - {1'b0, layer_2_2[4031:4024]};
      btm_2[2] = {1'b0,layer_3_2[4039:4032]} - {1'b0, layer_2_2[4039:4032]};
    end
    'd504: begin
      top_0[0] = {1'b0,layer_1_0[4031:4024]} - {1'b0, layer_0_0[4031:4024]};
      top_0[1] = {1'b0,layer_1_0[4039:4032]} - {1'b0, layer_0_0[4039:4032]};
      top_0[2] = {1'b0,layer_1_0[4047:4040]} - {1'b0, layer_0_0[4047:4040]};
      top_1[0] = {1'b0,layer_1_1[4031:4024]} - {1'b0, layer_0_1[4031:4024]};
      top_1[1] = {1'b0,layer_1_1[4039:4032]} - {1'b0, layer_0_1[4039:4032]};
      top_1[2] = {1'b0,layer_1_1[4047:4040]} - {1'b0, layer_0_1[4047:4040]};
      top_2[0] = {1'b0,layer_1_2[4031:4024]} - {1'b0, layer_0_2[4031:4024]};
      top_2[1] = {1'b0,layer_1_2[4039:4032]} - {1'b0, layer_0_2[4039:4032]};
      top_2[2] = {1'b0,layer_1_2[4047:4040]} - {1'b0, layer_0_2[4047:4040]};
      mid_0[0] = {1'b0,layer_2_0[4031:4024]} - {1'b0, layer_1_0[4031:4024]};
      mid_0[1] = {1'b0,layer_2_0[4039:4032]} - {1'b0, layer_1_0[4039:4032]};
      mid_0[2] = {1'b0,layer_2_0[4047:4040]} - {1'b0, layer_1_0[4047:4040]};
      mid_1[0] = {1'b0,layer_2_1[4031:4024]} - {1'b0, layer_1_1[4031:4024]};
      mid_1[1] = {1'b0,layer_2_1[4039:4032]} - {1'b0, layer_1_1[4039:4032]};
      mid_1[2] = {1'b0,layer_2_1[4047:4040]} - {1'b0, layer_1_1[4047:4040]};
      mid_2[0] = {1'b0,layer_2_2[4031:4024]} - {1'b0, layer_1_2[4031:4024]};
      mid_2[1] = {1'b0,layer_2_2[4039:4032]} - {1'b0, layer_1_2[4039:4032]};
      mid_2[2] = {1'b0,layer_2_2[4047:4040]} - {1'b0, layer_1_2[4047:4040]};
      btm_0[0] = {1'b0,layer_3_0[4031:4024]} - {1'b0, layer_2_0[4031:4024]};
      btm_0[1] = {1'b0,layer_3_0[4039:4032]} - {1'b0, layer_2_0[4039:4032]};
      btm_0[2] = {1'b0,layer_3_0[4047:4040]} - {1'b0, layer_2_0[4047:4040]};
      btm_1[0] = {1'b0,layer_3_1[4031:4024]} - {1'b0, layer_2_1[4031:4024]};
      btm_1[1] = {1'b0,layer_3_1[4039:4032]} - {1'b0, layer_2_1[4039:4032]};
      btm_1[2] = {1'b0,layer_3_1[4047:4040]} - {1'b0, layer_2_1[4047:4040]};
      btm_2[0] = {1'b0,layer_3_2[4031:4024]} - {1'b0, layer_2_2[4031:4024]};
      btm_2[1] = {1'b0,layer_3_2[4039:4032]} - {1'b0, layer_2_2[4039:4032]};
      btm_2[2] = {1'b0,layer_3_2[4047:4040]} - {1'b0, layer_2_2[4047:4040]};
    end
    'd505: begin
      top_0[0] = {1'b0,layer_1_0[4039:4032]} - {1'b0, layer_0_0[4039:4032]};
      top_0[1] = {1'b0,layer_1_0[4047:4040]} - {1'b0, layer_0_0[4047:4040]};
      top_0[2] = {1'b0,layer_1_0[4055:4048]} - {1'b0, layer_0_0[4055:4048]};
      top_1[0] = {1'b0,layer_1_1[4039:4032]} - {1'b0, layer_0_1[4039:4032]};
      top_1[1] = {1'b0,layer_1_1[4047:4040]} - {1'b0, layer_0_1[4047:4040]};
      top_1[2] = {1'b0,layer_1_1[4055:4048]} - {1'b0, layer_0_1[4055:4048]};
      top_2[0] = {1'b0,layer_1_2[4039:4032]} - {1'b0, layer_0_2[4039:4032]};
      top_2[1] = {1'b0,layer_1_2[4047:4040]} - {1'b0, layer_0_2[4047:4040]};
      top_2[2] = {1'b0,layer_1_2[4055:4048]} - {1'b0, layer_0_2[4055:4048]};
      mid_0[0] = {1'b0,layer_2_0[4039:4032]} - {1'b0, layer_1_0[4039:4032]};
      mid_0[1] = {1'b0,layer_2_0[4047:4040]} - {1'b0, layer_1_0[4047:4040]};
      mid_0[2] = {1'b0,layer_2_0[4055:4048]} - {1'b0, layer_1_0[4055:4048]};
      mid_1[0] = {1'b0,layer_2_1[4039:4032]} - {1'b0, layer_1_1[4039:4032]};
      mid_1[1] = {1'b0,layer_2_1[4047:4040]} - {1'b0, layer_1_1[4047:4040]};
      mid_1[2] = {1'b0,layer_2_1[4055:4048]} - {1'b0, layer_1_1[4055:4048]};
      mid_2[0] = {1'b0,layer_2_2[4039:4032]} - {1'b0, layer_1_2[4039:4032]};
      mid_2[1] = {1'b0,layer_2_2[4047:4040]} - {1'b0, layer_1_2[4047:4040]};
      mid_2[2] = {1'b0,layer_2_2[4055:4048]} - {1'b0, layer_1_2[4055:4048]};
      btm_0[0] = {1'b0,layer_3_0[4039:4032]} - {1'b0, layer_2_0[4039:4032]};
      btm_0[1] = {1'b0,layer_3_0[4047:4040]} - {1'b0, layer_2_0[4047:4040]};
      btm_0[2] = {1'b0,layer_3_0[4055:4048]} - {1'b0, layer_2_0[4055:4048]};
      btm_1[0] = {1'b0,layer_3_1[4039:4032]} - {1'b0, layer_2_1[4039:4032]};
      btm_1[1] = {1'b0,layer_3_1[4047:4040]} - {1'b0, layer_2_1[4047:4040]};
      btm_1[2] = {1'b0,layer_3_1[4055:4048]} - {1'b0, layer_2_1[4055:4048]};
      btm_2[0] = {1'b0,layer_3_2[4039:4032]} - {1'b0, layer_2_2[4039:4032]};
      btm_2[1] = {1'b0,layer_3_2[4047:4040]} - {1'b0, layer_2_2[4047:4040]};
      btm_2[2] = {1'b0,layer_3_2[4055:4048]} - {1'b0, layer_2_2[4055:4048]};
    end
    'd506: begin
      top_0[0] = {1'b0,layer_1_0[4047:4040]} - {1'b0, layer_0_0[4047:4040]};
      top_0[1] = {1'b0,layer_1_0[4055:4048]} - {1'b0, layer_0_0[4055:4048]};
      top_0[2] = {1'b0,layer_1_0[4063:4056]} - {1'b0, layer_0_0[4063:4056]};
      top_1[0] = {1'b0,layer_1_1[4047:4040]} - {1'b0, layer_0_1[4047:4040]};
      top_1[1] = {1'b0,layer_1_1[4055:4048]} - {1'b0, layer_0_1[4055:4048]};
      top_1[2] = {1'b0,layer_1_1[4063:4056]} - {1'b0, layer_0_1[4063:4056]};
      top_2[0] = {1'b0,layer_1_2[4047:4040]} - {1'b0, layer_0_2[4047:4040]};
      top_2[1] = {1'b0,layer_1_2[4055:4048]} - {1'b0, layer_0_2[4055:4048]};
      top_2[2] = {1'b0,layer_1_2[4063:4056]} - {1'b0, layer_0_2[4063:4056]};
      mid_0[0] = {1'b0,layer_2_0[4047:4040]} - {1'b0, layer_1_0[4047:4040]};
      mid_0[1] = {1'b0,layer_2_0[4055:4048]} - {1'b0, layer_1_0[4055:4048]};
      mid_0[2] = {1'b0,layer_2_0[4063:4056]} - {1'b0, layer_1_0[4063:4056]};
      mid_1[0] = {1'b0,layer_2_1[4047:4040]} - {1'b0, layer_1_1[4047:4040]};
      mid_1[1] = {1'b0,layer_2_1[4055:4048]} - {1'b0, layer_1_1[4055:4048]};
      mid_1[2] = {1'b0,layer_2_1[4063:4056]} - {1'b0, layer_1_1[4063:4056]};
      mid_2[0] = {1'b0,layer_2_2[4047:4040]} - {1'b0, layer_1_2[4047:4040]};
      mid_2[1] = {1'b0,layer_2_2[4055:4048]} - {1'b0, layer_1_2[4055:4048]};
      mid_2[2] = {1'b0,layer_2_2[4063:4056]} - {1'b0, layer_1_2[4063:4056]};
      btm_0[0] = {1'b0,layer_3_0[4047:4040]} - {1'b0, layer_2_0[4047:4040]};
      btm_0[1] = {1'b0,layer_3_0[4055:4048]} - {1'b0, layer_2_0[4055:4048]};
      btm_0[2] = {1'b0,layer_3_0[4063:4056]} - {1'b0, layer_2_0[4063:4056]};
      btm_1[0] = {1'b0,layer_3_1[4047:4040]} - {1'b0, layer_2_1[4047:4040]};
      btm_1[1] = {1'b0,layer_3_1[4055:4048]} - {1'b0, layer_2_1[4055:4048]};
      btm_1[2] = {1'b0,layer_3_1[4063:4056]} - {1'b0, layer_2_1[4063:4056]};
      btm_2[0] = {1'b0,layer_3_2[4047:4040]} - {1'b0, layer_2_2[4047:4040]};
      btm_2[1] = {1'b0,layer_3_2[4055:4048]} - {1'b0, layer_2_2[4055:4048]};
      btm_2[2] = {1'b0,layer_3_2[4063:4056]} - {1'b0, layer_2_2[4063:4056]};
    end
    'd507: begin
      top_0[0] = {1'b0,layer_1_0[4055:4048]} - {1'b0, layer_0_0[4055:4048]};
      top_0[1] = {1'b0,layer_1_0[4063:4056]} - {1'b0, layer_0_0[4063:4056]};
      top_0[2] = {1'b0,layer_1_0[4071:4064]} - {1'b0, layer_0_0[4071:4064]};
      top_1[0] = {1'b0,layer_1_1[4055:4048]} - {1'b0, layer_0_1[4055:4048]};
      top_1[1] = {1'b0,layer_1_1[4063:4056]} - {1'b0, layer_0_1[4063:4056]};
      top_1[2] = {1'b0,layer_1_1[4071:4064]} - {1'b0, layer_0_1[4071:4064]};
      top_2[0] = {1'b0,layer_1_2[4055:4048]} - {1'b0, layer_0_2[4055:4048]};
      top_2[1] = {1'b0,layer_1_2[4063:4056]} - {1'b0, layer_0_2[4063:4056]};
      top_2[2] = {1'b0,layer_1_2[4071:4064]} - {1'b0, layer_0_2[4071:4064]};
      mid_0[0] = {1'b0,layer_2_0[4055:4048]} - {1'b0, layer_1_0[4055:4048]};
      mid_0[1] = {1'b0,layer_2_0[4063:4056]} - {1'b0, layer_1_0[4063:4056]};
      mid_0[2] = {1'b0,layer_2_0[4071:4064]} - {1'b0, layer_1_0[4071:4064]};
      mid_1[0] = {1'b0,layer_2_1[4055:4048]} - {1'b0, layer_1_1[4055:4048]};
      mid_1[1] = {1'b0,layer_2_1[4063:4056]} - {1'b0, layer_1_1[4063:4056]};
      mid_1[2] = {1'b0,layer_2_1[4071:4064]} - {1'b0, layer_1_1[4071:4064]};
      mid_2[0] = {1'b0,layer_2_2[4055:4048]} - {1'b0, layer_1_2[4055:4048]};
      mid_2[1] = {1'b0,layer_2_2[4063:4056]} - {1'b0, layer_1_2[4063:4056]};
      mid_2[2] = {1'b0,layer_2_2[4071:4064]} - {1'b0, layer_1_2[4071:4064]};
      btm_0[0] = {1'b0,layer_3_0[4055:4048]} - {1'b0, layer_2_0[4055:4048]};
      btm_0[1] = {1'b0,layer_3_0[4063:4056]} - {1'b0, layer_2_0[4063:4056]};
      btm_0[2] = {1'b0,layer_3_0[4071:4064]} - {1'b0, layer_2_0[4071:4064]};
      btm_1[0] = {1'b0,layer_3_1[4055:4048]} - {1'b0, layer_2_1[4055:4048]};
      btm_1[1] = {1'b0,layer_3_1[4063:4056]} - {1'b0, layer_2_1[4063:4056]};
      btm_1[2] = {1'b0,layer_3_1[4071:4064]} - {1'b0, layer_2_1[4071:4064]};
      btm_2[0] = {1'b0,layer_3_2[4055:4048]} - {1'b0, layer_2_2[4055:4048]};
      btm_2[1] = {1'b0,layer_3_2[4063:4056]} - {1'b0, layer_2_2[4063:4056]};
      btm_2[2] = {1'b0,layer_3_2[4071:4064]} - {1'b0, layer_2_2[4071:4064]};
    end
    'd508: begin
      top_0[0] = {1'b0,layer_1_0[4063:4056]} - {1'b0, layer_0_0[4063:4056]};
      top_0[1] = {1'b0,layer_1_0[4071:4064]} - {1'b0, layer_0_0[4071:4064]};
      top_0[2] = {1'b0,layer_1_0[4079:4072]} - {1'b0, layer_0_0[4079:4072]};
      top_1[0] = {1'b0,layer_1_1[4063:4056]} - {1'b0, layer_0_1[4063:4056]};
      top_1[1] = {1'b0,layer_1_1[4071:4064]} - {1'b0, layer_0_1[4071:4064]};
      top_1[2] = {1'b0,layer_1_1[4079:4072]} - {1'b0, layer_0_1[4079:4072]};
      top_2[0] = {1'b0,layer_1_2[4063:4056]} - {1'b0, layer_0_2[4063:4056]};
      top_2[1] = {1'b0,layer_1_2[4071:4064]} - {1'b0, layer_0_2[4071:4064]};
      top_2[2] = {1'b0,layer_1_2[4079:4072]} - {1'b0, layer_0_2[4079:4072]};
      mid_0[0] = {1'b0,layer_2_0[4063:4056]} - {1'b0, layer_1_0[4063:4056]};
      mid_0[1] = {1'b0,layer_2_0[4071:4064]} - {1'b0, layer_1_0[4071:4064]};
      mid_0[2] = {1'b0,layer_2_0[4079:4072]} - {1'b0, layer_1_0[4079:4072]};
      mid_1[0] = {1'b0,layer_2_1[4063:4056]} - {1'b0, layer_1_1[4063:4056]};
      mid_1[1] = {1'b0,layer_2_1[4071:4064]} - {1'b0, layer_1_1[4071:4064]};
      mid_1[2] = {1'b0,layer_2_1[4079:4072]} - {1'b0, layer_1_1[4079:4072]};
      mid_2[0] = {1'b0,layer_2_2[4063:4056]} - {1'b0, layer_1_2[4063:4056]};
      mid_2[1] = {1'b0,layer_2_2[4071:4064]} - {1'b0, layer_1_2[4071:4064]};
      mid_2[2] = {1'b0,layer_2_2[4079:4072]} - {1'b0, layer_1_2[4079:4072]};
      btm_0[0] = {1'b0,layer_3_0[4063:4056]} - {1'b0, layer_2_0[4063:4056]};
      btm_0[1] = {1'b0,layer_3_0[4071:4064]} - {1'b0, layer_2_0[4071:4064]};
      btm_0[2] = {1'b0,layer_3_0[4079:4072]} - {1'b0, layer_2_0[4079:4072]};
      btm_1[0] = {1'b0,layer_3_1[4063:4056]} - {1'b0, layer_2_1[4063:4056]};
      btm_1[1] = {1'b0,layer_3_1[4071:4064]} - {1'b0, layer_2_1[4071:4064]};
      btm_1[2] = {1'b0,layer_3_1[4079:4072]} - {1'b0, layer_2_1[4079:4072]};
      btm_2[0] = {1'b0,layer_3_2[4063:4056]} - {1'b0, layer_2_2[4063:4056]};
      btm_2[1] = {1'b0,layer_3_2[4071:4064]} - {1'b0, layer_2_2[4071:4064]};
      btm_2[2] = {1'b0,layer_3_2[4079:4072]} - {1'b0, layer_2_2[4079:4072]};
    end
    'd509: begin
      top_0[0] = {1'b0,layer_1_0[4071:4064]} - {1'b0, layer_0_0[4071:4064]};
      top_0[1] = {1'b0,layer_1_0[4079:4072]} - {1'b0, layer_0_0[4079:4072]};
      top_0[2] = {1'b0,layer_1_0[4087:4080]} - {1'b0, layer_0_0[4087:4080]};
      top_1[0] = {1'b0,layer_1_1[4071:4064]} - {1'b0, layer_0_1[4071:4064]};
      top_1[1] = {1'b0,layer_1_1[4079:4072]} - {1'b0, layer_0_1[4079:4072]};
      top_1[2] = {1'b0,layer_1_1[4087:4080]} - {1'b0, layer_0_1[4087:4080]};
      top_2[0] = {1'b0,layer_1_2[4071:4064]} - {1'b0, layer_0_2[4071:4064]};
      top_2[1] = {1'b0,layer_1_2[4079:4072]} - {1'b0, layer_0_2[4079:4072]};
      top_2[2] = {1'b0,layer_1_2[4087:4080]} - {1'b0, layer_0_2[4087:4080]};
      mid_0[0] = {1'b0,layer_2_0[4071:4064]} - {1'b0, layer_1_0[4071:4064]};
      mid_0[1] = {1'b0,layer_2_0[4079:4072]} - {1'b0, layer_1_0[4079:4072]};
      mid_0[2] = {1'b0,layer_2_0[4087:4080]} - {1'b0, layer_1_0[4087:4080]};
      mid_1[0] = {1'b0,layer_2_1[4071:4064]} - {1'b0, layer_1_1[4071:4064]};
      mid_1[1] = {1'b0,layer_2_1[4079:4072]} - {1'b0, layer_1_1[4079:4072]};
      mid_1[2] = {1'b0,layer_2_1[4087:4080]} - {1'b0, layer_1_1[4087:4080]};
      mid_2[0] = {1'b0,layer_2_2[4071:4064]} - {1'b0, layer_1_2[4071:4064]};
      mid_2[1] = {1'b0,layer_2_2[4079:4072]} - {1'b0, layer_1_2[4079:4072]};
      mid_2[2] = {1'b0,layer_2_2[4087:4080]} - {1'b0, layer_1_2[4087:4080]};
      btm_0[0] = {1'b0,layer_3_0[4071:4064]} - {1'b0, layer_2_0[4071:4064]};
      btm_0[1] = {1'b0,layer_3_0[4079:4072]} - {1'b0, layer_2_0[4079:4072]};
      btm_0[2] = {1'b0,layer_3_0[4087:4080]} - {1'b0, layer_2_0[4087:4080]};
      btm_1[0] = {1'b0,layer_3_1[4071:4064]} - {1'b0, layer_2_1[4071:4064]};
      btm_1[1] = {1'b0,layer_3_1[4079:4072]} - {1'b0, layer_2_1[4079:4072]};
      btm_1[2] = {1'b0,layer_3_1[4087:4080]} - {1'b0, layer_2_1[4087:4080]};
      btm_2[0] = {1'b0,layer_3_2[4071:4064]} - {1'b0, layer_2_2[4071:4064]};
      btm_2[1] = {1'b0,layer_3_2[4079:4072]} - {1'b0, layer_2_2[4079:4072]};
      btm_2[2] = {1'b0,layer_3_2[4087:4080]} - {1'b0, layer_2_2[4087:4080]};
    end
    'd510: begin
      top_0[0] = {1'b0,layer_1_0[4079:4072]} - {1'b0, layer_0_0[4079:4072]};
      top_0[1] = {1'b0,layer_1_0[4087:4080]} - {1'b0, layer_0_0[4087:4080]};
      top_0[2] = {1'b0,layer_1_0[4095:4088]} - {1'b0, layer_0_0[4095:4088]};
      top_1[0] = {1'b0,layer_1_1[4079:4072]} - {1'b0, layer_0_1[4079:4072]};
      top_1[1] = {1'b0,layer_1_1[4087:4080]} - {1'b0, layer_0_1[4087:4080]};
      top_1[2] = {1'b0,layer_1_1[4095:4088]} - {1'b0, layer_0_1[4095:4088]};
      top_2[0] = {1'b0,layer_1_2[4079:4072]} - {1'b0, layer_0_2[4079:4072]};
      top_2[1] = {1'b0,layer_1_2[4087:4080]} - {1'b0, layer_0_2[4087:4080]};
      top_2[2] = {1'b0,layer_1_2[4095:4088]} - {1'b0, layer_0_2[4095:4088]};
      mid_0[0] = {1'b0,layer_2_0[4079:4072]} - {1'b0, layer_1_0[4079:4072]};
      mid_0[1] = {1'b0,layer_2_0[4087:4080]} - {1'b0, layer_1_0[4087:4080]};
      mid_0[2] = {1'b0,layer_2_0[4095:4088]} - {1'b0, layer_1_0[4095:4088]};
      mid_1[0] = {1'b0,layer_2_1[4079:4072]} - {1'b0, layer_1_1[4079:4072]};
      mid_1[1] = {1'b0,layer_2_1[4087:4080]} - {1'b0, layer_1_1[4087:4080]};
      mid_1[2] = {1'b0,layer_2_1[4095:4088]} - {1'b0, layer_1_1[4095:4088]};
      mid_2[0] = {1'b0,layer_2_2[4079:4072]} - {1'b0, layer_1_2[4079:4072]};
      mid_2[1] = {1'b0,layer_2_2[4087:4080]} - {1'b0, layer_1_2[4087:4080]};
      mid_2[2] = {1'b0,layer_2_2[4095:4088]} - {1'b0, layer_1_2[4095:4088]};
      btm_0[0] = {1'b0,layer_3_0[4079:4072]} - {1'b0, layer_2_0[4079:4072]};
      btm_0[1] = {1'b0,layer_3_0[4087:4080]} - {1'b0, layer_2_0[4087:4080]};
      btm_0[2] = {1'b0,layer_3_0[4095:4088]} - {1'b0, layer_2_0[4095:4088]};
      btm_1[0] = {1'b0,layer_3_1[4079:4072]} - {1'b0, layer_2_1[4079:4072]};
      btm_1[1] = {1'b0,layer_3_1[4087:4080]} - {1'b0, layer_2_1[4087:4080]};
      btm_1[2] = {1'b0,layer_3_1[4095:4088]} - {1'b0, layer_2_1[4095:4088]};
      btm_2[0] = {1'b0,layer_3_2[4079:4072]} - {1'b0, layer_2_2[4079:4072]};
      btm_2[1] = {1'b0,layer_3_2[4087:4080]} - {1'b0, layer_2_2[4087:4080]};
      btm_2[2] = {1'b0,layer_3_2[4095:4088]} - {1'b0, layer_2_2[4095:4088]};
    end
    'd511: begin
      top_0[0] = {1'b0,layer_1_0[4087:4080]} - {1'b0, layer_0_0[4087:4080]};
      top_0[1] = {1'b0,layer_1_0[4095:4088]} - {1'b0, layer_0_0[4095:4088]};
      top_0[2] = {1'b0,layer_1_0[4103:4096]} - {1'b0, layer_0_0[4103:4096]};
      top_1[0] = {1'b0,layer_1_1[4087:4080]} - {1'b0, layer_0_1[4087:4080]};
      top_1[1] = {1'b0,layer_1_1[4095:4088]} - {1'b0, layer_0_1[4095:4088]};
      top_1[2] = {1'b0,layer_1_1[4103:4096]} - {1'b0, layer_0_1[4103:4096]};
      top_2[0] = {1'b0,layer_1_2[4087:4080]} - {1'b0, layer_0_2[4087:4080]};
      top_2[1] = {1'b0,layer_1_2[4095:4088]} - {1'b0, layer_0_2[4095:4088]};
      top_2[2] = {1'b0,layer_1_2[4103:4096]} - {1'b0, layer_0_2[4103:4096]};
      mid_0[0] = {1'b0,layer_2_0[4087:4080]} - {1'b0, layer_1_0[4087:4080]};
      mid_0[1] = {1'b0,layer_2_0[4095:4088]} - {1'b0, layer_1_0[4095:4088]};
      mid_0[2] = {1'b0,layer_2_0[4103:4096]} - {1'b0, layer_1_0[4103:4096]};
      mid_1[0] = {1'b0,layer_2_1[4087:4080]} - {1'b0, layer_1_1[4087:4080]};
      mid_1[1] = {1'b0,layer_2_1[4095:4088]} - {1'b0, layer_1_1[4095:4088]};
      mid_1[2] = {1'b0,layer_2_1[4103:4096]} - {1'b0, layer_1_1[4103:4096]};
      mid_2[0] = {1'b0,layer_2_2[4087:4080]} - {1'b0, layer_1_2[4087:4080]};
      mid_2[1] = {1'b0,layer_2_2[4095:4088]} - {1'b0, layer_1_2[4095:4088]};
      mid_2[2] = {1'b0,layer_2_2[4103:4096]} - {1'b0, layer_1_2[4103:4096]};
      btm_0[0] = {1'b0,layer_3_0[4087:4080]} - {1'b0, layer_2_0[4087:4080]};
      btm_0[1] = {1'b0,layer_3_0[4095:4088]} - {1'b0, layer_2_0[4095:4088]};
      btm_0[2] = {1'b0,layer_3_0[4103:4096]} - {1'b0, layer_2_0[4103:4096]};
      btm_1[0] = {1'b0,layer_3_1[4087:4080]} - {1'b0, layer_2_1[4087:4080]};
      btm_1[1] = {1'b0,layer_3_1[4095:4088]} - {1'b0, layer_2_1[4095:4088]};
      btm_1[2] = {1'b0,layer_3_1[4103:4096]} - {1'b0, layer_2_1[4103:4096]};
      btm_2[0] = {1'b0,layer_3_2[4087:4080]} - {1'b0, layer_2_2[4087:4080]};
      btm_2[1] = {1'b0,layer_3_2[4095:4088]} - {1'b0, layer_2_2[4095:4088]};
      btm_2[2] = {1'b0,layer_3_2[4103:4096]} - {1'b0, layer_2_2[4103:4096]};
    end
    'd512: begin
      top_0[0] = {1'b0,layer_1_0[4095:4088]} - {1'b0, layer_0_0[4095:4088]};
      top_0[1] = {1'b0,layer_1_0[4103:4096]} - {1'b0, layer_0_0[4103:4096]};
      top_0[2] = {1'b0,layer_1_0[4111:4104]} - {1'b0, layer_0_0[4111:4104]};
      top_1[0] = {1'b0,layer_1_1[4095:4088]} - {1'b0, layer_0_1[4095:4088]};
      top_1[1] = {1'b0,layer_1_1[4103:4096]} - {1'b0, layer_0_1[4103:4096]};
      top_1[2] = {1'b0,layer_1_1[4111:4104]} - {1'b0, layer_0_1[4111:4104]};
      top_2[0] = {1'b0,layer_1_2[4095:4088]} - {1'b0, layer_0_2[4095:4088]};
      top_2[1] = {1'b0,layer_1_2[4103:4096]} - {1'b0, layer_0_2[4103:4096]};
      top_2[2] = {1'b0,layer_1_2[4111:4104]} - {1'b0, layer_0_2[4111:4104]};
      mid_0[0] = {1'b0,layer_2_0[4095:4088]} - {1'b0, layer_1_0[4095:4088]};
      mid_0[1] = {1'b0,layer_2_0[4103:4096]} - {1'b0, layer_1_0[4103:4096]};
      mid_0[2] = {1'b0,layer_2_0[4111:4104]} - {1'b0, layer_1_0[4111:4104]};
      mid_1[0] = {1'b0,layer_2_1[4095:4088]} - {1'b0, layer_1_1[4095:4088]};
      mid_1[1] = {1'b0,layer_2_1[4103:4096]} - {1'b0, layer_1_1[4103:4096]};
      mid_1[2] = {1'b0,layer_2_1[4111:4104]} - {1'b0, layer_1_1[4111:4104]};
      mid_2[0] = {1'b0,layer_2_2[4095:4088]} - {1'b0, layer_1_2[4095:4088]};
      mid_2[1] = {1'b0,layer_2_2[4103:4096]} - {1'b0, layer_1_2[4103:4096]};
      mid_2[2] = {1'b0,layer_2_2[4111:4104]} - {1'b0, layer_1_2[4111:4104]};
      btm_0[0] = {1'b0,layer_3_0[4095:4088]} - {1'b0, layer_2_0[4095:4088]};
      btm_0[1] = {1'b0,layer_3_0[4103:4096]} - {1'b0, layer_2_0[4103:4096]};
      btm_0[2] = {1'b0,layer_3_0[4111:4104]} - {1'b0, layer_2_0[4111:4104]};
      btm_1[0] = {1'b0,layer_3_1[4095:4088]} - {1'b0, layer_2_1[4095:4088]};
      btm_1[1] = {1'b0,layer_3_1[4103:4096]} - {1'b0, layer_2_1[4103:4096]};
      btm_1[2] = {1'b0,layer_3_1[4111:4104]} - {1'b0, layer_2_1[4111:4104]};
      btm_2[0] = {1'b0,layer_3_2[4095:4088]} - {1'b0, layer_2_2[4095:4088]};
      btm_2[1] = {1'b0,layer_3_2[4103:4096]} - {1'b0, layer_2_2[4103:4096]};
      btm_2[2] = {1'b0,layer_3_2[4111:4104]} - {1'b0, layer_2_2[4111:4104]};
    end
    'd513: begin
      top_0[0] = {1'b0,layer_1_0[4103:4096]} - {1'b0, layer_0_0[4103:4096]};
      top_0[1] = {1'b0,layer_1_0[4111:4104]} - {1'b0, layer_0_0[4111:4104]};
      top_0[2] = {1'b0,layer_1_0[4119:4112]} - {1'b0, layer_0_0[4119:4112]};
      top_1[0] = {1'b0,layer_1_1[4103:4096]} - {1'b0, layer_0_1[4103:4096]};
      top_1[1] = {1'b0,layer_1_1[4111:4104]} - {1'b0, layer_0_1[4111:4104]};
      top_1[2] = {1'b0,layer_1_1[4119:4112]} - {1'b0, layer_0_1[4119:4112]};
      top_2[0] = {1'b0,layer_1_2[4103:4096]} - {1'b0, layer_0_2[4103:4096]};
      top_2[1] = {1'b0,layer_1_2[4111:4104]} - {1'b0, layer_0_2[4111:4104]};
      top_2[2] = {1'b0,layer_1_2[4119:4112]} - {1'b0, layer_0_2[4119:4112]};
      mid_0[0] = {1'b0,layer_2_0[4103:4096]} - {1'b0, layer_1_0[4103:4096]};
      mid_0[1] = {1'b0,layer_2_0[4111:4104]} - {1'b0, layer_1_0[4111:4104]};
      mid_0[2] = {1'b0,layer_2_0[4119:4112]} - {1'b0, layer_1_0[4119:4112]};
      mid_1[0] = {1'b0,layer_2_1[4103:4096]} - {1'b0, layer_1_1[4103:4096]};
      mid_1[1] = {1'b0,layer_2_1[4111:4104]} - {1'b0, layer_1_1[4111:4104]};
      mid_1[2] = {1'b0,layer_2_1[4119:4112]} - {1'b0, layer_1_1[4119:4112]};
      mid_2[0] = {1'b0,layer_2_2[4103:4096]} - {1'b0, layer_1_2[4103:4096]};
      mid_2[1] = {1'b0,layer_2_2[4111:4104]} - {1'b0, layer_1_2[4111:4104]};
      mid_2[2] = {1'b0,layer_2_2[4119:4112]} - {1'b0, layer_1_2[4119:4112]};
      btm_0[0] = {1'b0,layer_3_0[4103:4096]} - {1'b0, layer_2_0[4103:4096]};
      btm_0[1] = {1'b0,layer_3_0[4111:4104]} - {1'b0, layer_2_0[4111:4104]};
      btm_0[2] = {1'b0,layer_3_0[4119:4112]} - {1'b0, layer_2_0[4119:4112]};
      btm_1[0] = {1'b0,layer_3_1[4103:4096]} - {1'b0, layer_2_1[4103:4096]};
      btm_1[1] = {1'b0,layer_3_1[4111:4104]} - {1'b0, layer_2_1[4111:4104]};
      btm_1[2] = {1'b0,layer_3_1[4119:4112]} - {1'b0, layer_2_1[4119:4112]};
      btm_2[0] = {1'b0,layer_3_2[4103:4096]} - {1'b0, layer_2_2[4103:4096]};
      btm_2[1] = {1'b0,layer_3_2[4111:4104]} - {1'b0, layer_2_2[4111:4104]};
      btm_2[2] = {1'b0,layer_3_2[4119:4112]} - {1'b0, layer_2_2[4119:4112]};
    end
    'd514: begin
      top_0[0] = {1'b0,layer_1_0[4111:4104]} - {1'b0, layer_0_0[4111:4104]};
      top_0[1] = {1'b0,layer_1_0[4119:4112]} - {1'b0, layer_0_0[4119:4112]};
      top_0[2] = {1'b0,layer_1_0[4127:4120]} - {1'b0, layer_0_0[4127:4120]};
      top_1[0] = {1'b0,layer_1_1[4111:4104]} - {1'b0, layer_0_1[4111:4104]};
      top_1[1] = {1'b0,layer_1_1[4119:4112]} - {1'b0, layer_0_1[4119:4112]};
      top_1[2] = {1'b0,layer_1_1[4127:4120]} - {1'b0, layer_0_1[4127:4120]};
      top_2[0] = {1'b0,layer_1_2[4111:4104]} - {1'b0, layer_0_2[4111:4104]};
      top_2[1] = {1'b0,layer_1_2[4119:4112]} - {1'b0, layer_0_2[4119:4112]};
      top_2[2] = {1'b0,layer_1_2[4127:4120]} - {1'b0, layer_0_2[4127:4120]};
      mid_0[0] = {1'b0,layer_2_0[4111:4104]} - {1'b0, layer_1_0[4111:4104]};
      mid_0[1] = {1'b0,layer_2_0[4119:4112]} - {1'b0, layer_1_0[4119:4112]};
      mid_0[2] = {1'b0,layer_2_0[4127:4120]} - {1'b0, layer_1_0[4127:4120]};
      mid_1[0] = {1'b0,layer_2_1[4111:4104]} - {1'b0, layer_1_1[4111:4104]};
      mid_1[1] = {1'b0,layer_2_1[4119:4112]} - {1'b0, layer_1_1[4119:4112]};
      mid_1[2] = {1'b0,layer_2_1[4127:4120]} - {1'b0, layer_1_1[4127:4120]};
      mid_2[0] = {1'b0,layer_2_2[4111:4104]} - {1'b0, layer_1_2[4111:4104]};
      mid_2[1] = {1'b0,layer_2_2[4119:4112]} - {1'b0, layer_1_2[4119:4112]};
      mid_2[2] = {1'b0,layer_2_2[4127:4120]} - {1'b0, layer_1_2[4127:4120]};
      btm_0[0] = {1'b0,layer_3_0[4111:4104]} - {1'b0, layer_2_0[4111:4104]};
      btm_0[1] = {1'b0,layer_3_0[4119:4112]} - {1'b0, layer_2_0[4119:4112]};
      btm_0[2] = {1'b0,layer_3_0[4127:4120]} - {1'b0, layer_2_0[4127:4120]};
      btm_1[0] = {1'b0,layer_3_1[4111:4104]} - {1'b0, layer_2_1[4111:4104]};
      btm_1[1] = {1'b0,layer_3_1[4119:4112]} - {1'b0, layer_2_1[4119:4112]};
      btm_1[2] = {1'b0,layer_3_1[4127:4120]} - {1'b0, layer_2_1[4127:4120]};
      btm_2[0] = {1'b0,layer_3_2[4111:4104]} - {1'b0, layer_2_2[4111:4104]};
      btm_2[1] = {1'b0,layer_3_2[4119:4112]} - {1'b0, layer_2_2[4119:4112]};
      btm_2[2] = {1'b0,layer_3_2[4127:4120]} - {1'b0, layer_2_2[4127:4120]};
    end
    'd515: begin
      top_0[0] = {1'b0,layer_1_0[4119:4112]} - {1'b0, layer_0_0[4119:4112]};
      top_0[1] = {1'b0,layer_1_0[4127:4120]} - {1'b0, layer_0_0[4127:4120]};
      top_0[2] = {1'b0,layer_1_0[4135:4128]} - {1'b0, layer_0_0[4135:4128]};
      top_1[0] = {1'b0,layer_1_1[4119:4112]} - {1'b0, layer_0_1[4119:4112]};
      top_1[1] = {1'b0,layer_1_1[4127:4120]} - {1'b0, layer_0_1[4127:4120]};
      top_1[2] = {1'b0,layer_1_1[4135:4128]} - {1'b0, layer_0_1[4135:4128]};
      top_2[0] = {1'b0,layer_1_2[4119:4112]} - {1'b0, layer_0_2[4119:4112]};
      top_2[1] = {1'b0,layer_1_2[4127:4120]} - {1'b0, layer_0_2[4127:4120]};
      top_2[2] = {1'b0,layer_1_2[4135:4128]} - {1'b0, layer_0_2[4135:4128]};
      mid_0[0] = {1'b0,layer_2_0[4119:4112]} - {1'b0, layer_1_0[4119:4112]};
      mid_0[1] = {1'b0,layer_2_0[4127:4120]} - {1'b0, layer_1_0[4127:4120]};
      mid_0[2] = {1'b0,layer_2_0[4135:4128]} - {1'b0, layer_1_0[4135:4128]};
      mid_1[0] = {1'b0,layer_2_1[4119:4112]} - {1'b0, layer_1_1[4119:4112]};
      mid_1[1] = {1'b0,layer_2_1[4127:4120]} - {1'b0, layer_1_1[4127:4120]};
      mid_1[2] = {1'b0,layer_2_1[4135:4128]} - {1'b0, layer_1_1[4135:4128]};
      mid_2[0] = {1'b0,layer_2_2[4119:4112]} - {1'b0, layer_1_2[4119:4112]};
      mid_2[1] = {1'b0,layer_2_2[4127:4120]} - {1'b0, layer_1_2[4127:4120]};
      mid_2[2] = {1'b0,layer_2_2[4135:4128]} - {1'b0, layer_1_2[4135:4128]};
      btm_0[0] = {1'b0,layer_3_0[4119:4112]} - {1'b0, layer_2_0[4119:4112]};
      btm_0[1] = {1'b0,layer_3_0[4127:4120]} - {1'b0, layer_2_0[4127:4120]};
      btm_0[2] = {1'b0,layer_3_0[4135:4128]} - {1'b0, layer_2_0[4135:4128]};
      btm_1[0] = {1'b0,layer_3_1[4119:4112]} - {1'b0, layer_2_1[4119:4112]};
      btm_1[1] = {1'b0,layer_3_1[4127:4120]} - {1'b0, layer_2_1[4127:4120]};
      btm_1[2] = {1'b0,layer_3_1[4135:4128]} - {1'b0, layer_2_1[4135:4128]};
      btm_2[0] = {1'b0,layer_3_2[4119:4112]} - {1'b0, layer_2_2[4119:4112]};
      btm_2[1] = {1'b0,layer_3_2[4127:4120]} - {1'b0, layer_2_2[4127:4120]};
      btm_2[2] = {1'b0,layer_3_2[4135:4128]} - {1'b0, layer_2_2[4135:4128]};
    end
    'd516: begin
      top_0[0] = {1'b0,layer_1_0[4127:4120]} - {1'b0, layer_0_0[4127:4120]};
      top_0[1] = {1'b0,layer_1_0[4135:4128]} - {1'b0, layer_0_0[4135:4128]};
      top_0[2] = {1'b0,layer_1_0[4143:4136]} - {1'b0, layer_0_0[4143:4136]};
      top_1[0] = {1'b0,layer_1_1[4127:4120]} - {1'b0, layer_0_1[4127:4120]};
      top_1[1] = {1'b0,layer_1_1[4135:4128]} - {1'b0, layer_0_1[4135:4128]};
      top_1[2] = {1'b0,layer_1_1[4143:4136]} - {1'b0, layer_0_1[4143:4136]};
      top_2[0] = {1'b0,layer_1_2[4127:4120]} - {1'b0, layer_0_2[4127:4120]};
      top_2[1] = {1'b0,layer_1_2[4135:4128]} - {1'b0, layer_0_2[4135:4128]};
      top_2[2] = {1'b0,layer_1_2[4143:4136]} - {1'b0, layer_0_2[4143:4136]};
      mid_0[0] = {1'b0,layer_2_0[4127:4120]} - {1'b0, layer_1_0[4127:4120]};
      mid_0[1] = {1'b0,layer_2_0[4135:4128]} - {1'b0, layer_1_0[4135:4128]};
      mid_0[2] = {1'b0,layer_2_0[4143:4136]} - {1'b0, layer_1_0[4143:4136]};
      mid_1[0] = {1'b0,layer_2_1[4127:4120]} - {1'b0, layer_1_1[4127:4120]};
      mid_1[1] = {1'b0,layer_2_1[4135:4128]} - {1'b0, layer_1_1[4135:4128]};
      mid_1[2] = {1'b0,layer_2_1[4143:4136]} - {1'b0, layer_1_1[4143:4136]};
      mid_2[0] = {1'b0,layer_2_2[4127:4120]} - {1'b0, layer_1_2[4127:4120]};
      mid_2[1] = {1'b0,layer_2_2[4135:4128]} - {1'b0, layer_1_2[4135:4128]};
      mid_2[2] = {1'b0,layer_2_2[4143:4136]} - {1'b0, layer_1_2[4143:4136]};
      btm_0[0] = {1'b0,layer_3_0[4127:4120]} - {1'b0, layer_2_0[4127:4120]};
      btm_0[1] = {1'b0,layer_3_0[4135:4128]} - {1'b0, layer_2_0[4135:4128]};
      btm_0[2] = {1'b0,layer_3_0[4143:4136]} - {1'b0, layer_2_0[4143:4136]};
      btm_1[0] = {1'b0,layer_3_1[4127:4120]} - {1'b0, layer_2_1[4127:4120]};
      btm_1[1] = {1'b0,layer_3_1[4135:4128]} - {1'b0, layer_2_1[4135:4128]};
      btm_1[2] = {1'b0,layer_3_1[4143:4136]} - {1'b0, layer_2_1[4143:4136]};
      btm_2[0] = {1'b0,layer_3_2[4127:4120]} - {1'b0, layer_2_2[4127:4120]};
      btm_2[1] = {1'b0,layer_3_2[4135:4128]} - {1'b0, layer_2_2[4135:4128]};
      btm_2[2] = {1'b0,layer_3_2[4143:4136]} - {1'b0, layer_2_2[4143:4136]};
    end
    'd517: begin
      top_0[0] = {1'b0,layer_1_0[4135:4128]} - {1'b0, layer_0_0[4135:4128]};
      top_0[1] = {1'b0,layer_1_0[4143:4136]} - {1'b0, layer_0_0[4143:4136]};
      top_0[2] = {1'b0,layer_1_0[4151:4144]} - {1'b0, layer_0_0[4151:4144]};
      top_1[0] = {1'b0,layer_1_1[4135:4128]} - {1'b0, layer_0_1[4135:4128]};
      top_1[1] = {1'b0,layer_1_1[4143:4136]} - {1'b0, layer_0_1[4143:4136]};
      top_1[2] = {1'b0,layer_1_1[4151:4144]} - {1'b0, layer_0_1[4151:4144]};
      top_2[0] = {1'b0,layer_1_2[4135:4128]} - {1'b0, layer_0_2[4135:4128]};
      top_2[1] = {1'b0,layer_1_2[4143:4136]} - {1'b0, layer_0_2[4143:4136]};
      top_2[2] = {1'b0,layer_1_2[4151:4144]} - {1'b0, layer_0_2[4151:4144]};
      mid_0[0] = {1'b0,layer_2_0[4135:4128]} - {1'b0, layer_1_0[4135:4128]};
      mid_0[1] = {1'b0,layer_2_0[4143:4136]} - {1'b0, layer_1_0[4143:4136]};
      mid_0[2] = {1'b0,layer_2_0[4151:4144]} - {1'b0, layer_1_0[4151:4144]};
      mid_1[0] = {1'b0,layer_2_1[4135:4128]} - {1'b0, layer_1_1[4135:4128]};
      mid_1[1] = {1'b0,layer_2_1[4143:4136]} - {1'b0, layer_1_1[4143:4136]};
      mid_1[2] = {1'b0,layer_2_1[4151:4144]} - {1'b0, layer_1_1[4151:4144]};
      mid_2[0] = {1'b0,layer_2_2[4135:4128]} - {1'b0, layer_1_2[4135:4128]};
      mid_2[1] = {1'b0,layer_2_2[4143:4136]} - {1'b0, layer_1_2[4143:4136]};
      mid_2[2] = {1'b0,layer_2_2[4151:4144]} - {1'b0, layer_1_2[4151:4144]};
      btm_0[0] = {1'b0,layer_3_0[4135:4128]} - {1'b0, layer_2_0[4135:4128]};
      btm_0[1] = {1'b0,layer_3_0[4143:4136]} - {1'b0, layer_2_0[4143:4136]};
      btm_0[2] = {1'b0,layer_3_0[4151:4144]} - {1'b0, layer_2_0[4151:4144]};
      btm_1[0] = {1'b0,layer_3_1[4135:4128]} - {1'b0, layer_2_1[4135:4128]};
      btm_1[1] = {1'b0,layer_3_1[4143:4136]} - {1'b0, layer_2_1[4143:4136]};
      btm_1[2] = {1'b0,layer_3_1[4151:4144]} - {1'b0, layer_2_1[4151:4144]};
      btm_2[0] = {1'b0,layer_3_2[4135:4128]} - {1'b0, layer_2_2[4135:4128]};
      btm_2[1] = {1'b0,layer_3_2[4143:4136]} - {1'b0, layer_2_2[4143:4136]};
      btm_2[2] = {1'b0,layer_3_2[4151:4144]} - {1'b0, layer_2_2[4151:4144]};
    end
    'd518: begin
      top_0[0] = {1'b0,layer_1_0[4143:4136]} - {1'b0, layer_0_0[4143:4136]};
      top_0[1] = {1'b0,layer_1_0[4151:4144]} - {1'b0, layer_0_0[4151:4144]};
      top_0[2] = {1'b0,layer_1_0[4159:4152]} - {1'b0, layer_0_0[4159:4152]};
      top_1[0] = {1'b0,layer_1_1[4143:4136]} - {1'b0, layer_0_1[4143:4136]};
      top_1[1] = {1'b0,layer_1_1[4151:4144]} - {1'b0, layer_0_1[4151:4144]};
      top_1[2] = {1'b0,layer_1_1[4159:4152]} - {1'b0, layer_0_1[4159:4152]};
      top_2[0] = {1'b0,layer_1_2[4143:4136]} - {1'b0, layer_0_2[4143:4136]};
      top_2[1] = {1'b0,layer_1_2[4151:4144]} - {1'b0, layer_0_2[4151:4144]};
      top_2[2] = {1'b0,layer_1_2[4159:4152]} - {1'b0, layer_0_2[4159:4152]};
      mid_0[0] = {1'b0,layer_2_0[4143:4136]} - {1'b0, layer_1_0[4143:4136]};
      mid_0[1] = {1'b0,layer_2_0[4151:4144]} - {1'b0, layer_1_0[4151:4144]};
      mid_0[2] = {1'b0,layer_2_0[4159:4152]} - {1'b0, layer_1_0[4159:4152]};
      mid_1[0] = {1'b0,layer_2_1[4143:4136]} - {1'b0, layer_1_1[4143:4136]};
      mid_1[1] = {1'b0,layer_2_1[4151:4144]} - {1'b0, layer_1_1[4151:4144]};
      mid_1[2] = {1'b0,layer_2_1[4159:4152]} - {1'b0, layer_1_1[4159:4152]};
      mid_2[0] = {1'b0,layer_2_2[4143:4136]} - {1'b0, layer_1_2[4143:4136]};
      mid_2[1] = {1'b0,layer_2_2[4151:4144]} - {1'b0, layer_1_2[4151:4144]};
      mid_2[2] = {1'b0,layer_2_2[4159:4152]} - {1'b0, layer_1_2[4159:4152]};
      btm_0[0] = {1'b0,layer_3_0[4143:4136]} - {1'b0, layer_2_0[4143:4136]};
      btm_0[1] = {1'b0,layer_3_0[4151:4144]} - {1'b0, layer_2_0[4151:4144]};
      btm_0[2] = {1'b0,layer_3_0[4159:4152]} - {1'b0, layer_2_0[4159:4152]};
      btm_1[0] = {1'b0,layer_3_1[4143:4136]} - {1'b0, layer_2_1[4143:4136]};
      btm_1[1] = {1'b0,layer_3_1[4151:4144]} - {1'b0, layer_2_1[4151:4144]};
      btm_1[2] = {1'b0,layer_3_1[4159:4152]} - {1'b0, layer_2_1[4159:4152]};
      btm_2[0] = {1'b0,layer_3_2[4143:4136]} - {1'b0, layer_2_2[4143:4136]};
      btm_2[1] = {1'b0,layer_3_2[4151:4144]} - {1'b0, layer_2_2[4151:4144]};
      btm_2[2] = {1'b0,layer_3_2[4159:4152]} - {1'b0, layer_2_2[4159:4152]};
    end
    'd519: begin
      top_0[0] = {1'b0,layer_1_0[4151:4144]} - {1'b0, layer_0_0[4151:4144]};
      top_0[1] = {1'b0,layer_1_0[4159:4152]} - {1'b0, layer_0_0[4159:4152]};
      top_0[2] = {1'b0,layer_1_0[4167:4160]} - {1'b0, layer_0_0[4167:4160]};
      top_1[0] = {1'b0,layer_1_1[4151:4144]} - {1'b0, layer_0_1[4151:4144]};
      top_1[1] = {1'b0,layer_1_1[4159:4152]} - {1'b0, layer_0_1[4159:4152]};
      top_1[2] = {1'b0,layer_1_1[4167:4160]} - {1'b0, layer_0_1[4167:4160]};
      top_2[0] = {1'b0,layer_1_2[4151:4144]} - {1'b0, layer_0_2[4151:4144]};
      top_2[1] = {1'b0,layer_1_2[4159:4152]} - {1'b0, layer_0_2[4159:4152]};
      top_2[2] = {1'b0,layer_1_2[4167:4160]} - {1'b0, layer_0_2[4167:4160]};
      mid_0[0] = {1'b0,layer_2_0[4151:4144]} - {1'b0, layer_1_0[4151:4144]};
      mid_0[1] = {1'b0,layer_2_0[4159:4152]} - {1'b0, layer_1_0[4159:4152]};
      mid_0[2] = {1'b0,layer_2_0[4167:4160]} - {1'b0, layer_1_0[4167:4160]};
      mid_1[0] = {1'b0,layer_2_1[4151:4144]} - {1'b0, layer_1_1[4151:4144]};
      mid_1[1] = {1'b0,layer_2_1[4159:4152]} - {1'b0, layer_1_1[4159:4152]};
      mid_1[2] = {1'b0,layer_2_1[4167:4160]} - {1'b0, layer_1_1[4167:4160]};
      mid_2[0] = {1'b0,layer_2_2[4151:4144]} - {1'b0, layer_1_2[4151:4144]};
      mid_2[1] = {1'b0,layer_2_2[4159:4152]} - {1'b0, layer_1_2[4159:4152]};
      mid_2[2] = {1'b0,layer_2_2[4167:4160]} - {1'b0, layer_1_2[4167:4160]};
      btm_0[0] = {1'b0,layer_3_0[4151:4144]} - {1'b0, layer_2_0[4151:4144]};
      btm_0[1] = {1'b0,layer_3_0[4159:4152]} - {1'b0, layer_2_0[4159:4152]};
      btm_0[2] = {1'b0,layer_3_0[4167:4160]} - {1'b0, layer_2_0[4167:4160]};
      btm_1[0] = {1'b0,layer_3_1[4151:4144]} - {1'b0, layer_2_1[4151:4144]};
      btm_1[1] = {1'b0,layer_3_1[4159:4152]} - {1'b0, layer_2_1[4159:4152]};
      btm_1[2] = {1'b0,layer_3_1[4167:4160]} - {1'b0, layer_2_1[4167:4160]};
      btm_2[0] = {1'b0,layer_3_2[4151:4144]} - {1'b0, layer_2_2[4151:4144]};
      btm_2[1] = {1'b0,layer_3_2[4159:4152]} - {1'b0, layer_2_2[4159:4152]};
      btm_2[2] = {1'b0,layer_3_2[4167:4160]} - {1'b0, layer_2_2[4167:4160]};
    end
    'd520: begin
      top_0[0] = {1'b0,layer_1_0[4159:4152]} - {1'b0, layer_0_0[4159:4152]};
      top_0[1] = {1'b0,layer_1_0[4167:4160]} - {1'b0, layer_0_0[4167:4160]};
      top_0[2] = {1'b0,layer_1_0[4175:4168]} - {1'b0, layer_0_0[4175:4168]};
      top_1[0] = {1'b0,layer_1_1[4159:4152]} - {1'b0, layer_0_1[4159:4152]};
      top_1[1] = {1'b0,layer_1_1[4167:4160]} - {1'b0, layer_0_1[4167:4160]};
      top_1[2] = {1'b0,layer_1_1[4175:4168]} - {1'b0, layer_0_1[4175:4168]};
      top_2[0] = {1'b0,layer_1_2[4159:4152]} - {1'b0, layer_0_2[4159:4152]};
      top_2[1] = {1'b0,layer_1_2[4167:4160]} - {1'b0, layer_0_2[4167:4160]};
      top_2[2] = {1'b0,layer_1_2[4175:4168]} - {1'b0, layer_0_2[4175:4168]};
      mid_0[0] = {1'b0,layer_2_0[4159:4152]} - {1'b0, layer_1_0[4159:4152]};
      mid_0[1] = {1'b0,layer_2_0[4167:4160]} - {1'b0, layer_1_0[4167:4160]};
      mid_0[2] = {1'b0,layer_2_0[4175:4168]} - {1'b0, layer_1_0[4175:4168]};
      mid_1[0] = {1'b0,layer_2_1[4159:4152]} - {1'b0, layer_1_1[4159:4152]};
      mid_1[1] = {1'b0,layer_2_1[4167:4160]} - {1'b0, layer_1_1[4167:4160]};
      mid_1[2] = {1'b0,layer_2_1[4175:4168]} - {1'b0, layer_1_1[4175:4168]};
      mid_2[0] = {1'b0,layer_2_2[4159:4152]} - {1'b0, layer_1_2[4159:4152]};
      mid_2[1] = {1'b0,layer_2_2[4167:4160]} - {1'b0, layer_1_2[4167:4160]};
      mid_2[2] = {1'b0,layer_2_2[4175:4168]} - {1'b0, layer_1_2[4175:4168]};
      btm_0[0] = {1'b0,layer_3_0[4159:4152]} - {1'b0, layer_2_0[4159:4152]};
      btm_0[1] = {1'b0,layer_3_0[4167:4160]} - {1'b0, layer_2_0[4167:4160]};
      btm_0[2] = {1'b0,layer_3_0[4175:4168]} - {1'b0, layer_2_0[4175:4168]};
      btm_1[0] = {1'b0,layer_3_1[4159:4152]} - {1'b0, layer_2_1[4159:4152]};
      btm_1[1] = {1'b0,layer_3_1[4167:4160]} - {1'b0, layer_2_1[4167:4160]};
      btm_1[2] = {1'b0,layer_3_1[4175:4168]} - {1'b0, layer_2_1[4175:4168]};
      btm_2[0] = {1'b0,layer_3_2[4159:4152]} - {1'b0, layer_2_2[4159:4152]};
      btm_2[1] = {1'b0,layer_3_2[4167:4160]} - {1'b0, layer_2_2[4167:4160]};
      btm_2[2] = {1'b0,layer_3_2[4175:4168]} - {1'b0, layer_2_2[4175:4168]};
    end
    'd521: begin
      top_0[0] = {1'b0,layer_1_0[4167:4160]} - {1'b0, layer_0_0[4167:4160]};
      top_0[1] = {1'b0,layer_1_0[4175:4168]} - {1'b0, layer_0_0[4175:4168]};
      top_0[2] = {1'b0,layer_1_0[4183:4176]} - {1'b0, layer_0_0[4183:4176]};
      top_1[0] = {1'b0,layer_1_1[4167:4160]} - {1'b0, layer_0_1[4167:4160]};
      top_1[1] = {1'b0,layer_1_1[4175:4168]} - {1'b0, layer_0_1[4175:4168]};
      top_1[2] = {1'b0,layer_1_1[4183:4176]} - {1'b0, layer_0_1[4183:4176]};
      top_2[0] = {1'b0,layer_1_2[4167:4160]} - {1'b0, layer_0_2[4167:4160]};
      top_2[1] = {1'b0,layer_1_2[4175:4168]} - {1'b0, layer_0_2[4175:4168]};
      top_2[2] = {1'b0,layer_1_2[4183:4176]} - {1'b0, layer_0_2[4183:4176]};
      mid_0[0] = {1'b0,layer_2_0[4167:4160]} - {1'b0, layer_1_0[4167:4160]};
      mid_0[1] = {1'b0,layer_2_0[4175:4168]} - {1'b0, layer_1_0[4175:4168]};
      mid_0[2] = {1'b0,layer_2_0[4183:4176]} - {1'b0, layer_1_0[4183:4176]};
      mid_1[0] = {1'b0,layer_2_1[4167:4160]} - {1'b0, layer_1_1[4167:4160]};
      mid_1[1] = {1'b0,layer_2_1[4175:4168]} - {1'b0, layer_1_1[4175:4168]};
      mid_1[2] = {1'b0,layer_2_1[4183:4176]} - {1'b0, layer_1_1[4183:4176]};
      mid_2[0] = {1'b0,layer_2_2[4167:4160]} - {1'b0, layer_1_2[4167:4160]};
      mid_2[1] = {1'b0,layer_2_2[4175:4168]} - {1'b0, layer_1_2[4175:4168]};
      mid_2[2] = {1'b0,layer_2_2[4183:4176]} - {1'b0, layer_1_2[4183:4176]};
      btm_0[0] = {1'b0,layer_3_0[4167:4160]} - {1'b0, layer_2_0[4167:4160]};
      btm_0[1] = {1'b0,layer_3_0[4175:4168]} - {1'b0, layer_2_0[4175:4168]};
      btm_0[2] = {1'b0,layer_3_0[4183:4176]} - {1'b0, layer_2_0[4183:4176]};
      btm_1[0] = {1'b0,layer_3_1[4167:4160]} - {1'b0, layer_2_1[4167:4160]};
      btm_1[1] = {1'b0,layer_3_1[4175:4168]} - {1'b0, layer_2_1[4175:4168]};
      btm_1[2] = {1'b0,layer_3_1[4183:4176]} - {1'b0, layer_2_1[4183:4176]};
      btm_2[0] = {1'b0,layer_3_2[4167:4160]} - {1'b0, layer_2_2[4167:4160]};
      btm_2[1] = {1'b0,layer_3_2[4175:4168]} - {1'b0, layer_2_2[4175:4168]};
      btm_2[2] = {1'b0,layer_3_2[4183:4176]} - {1'b0, layer_2_2[4183:4176]};
    end
    'd522: begin
      top_0[0] = {1'b0,layer_1_0[4175:4168]} - {1'b0, layer_0_0[4175:4168]};
      top_0[1] = {1'b0,layer_1_0[4183:4176]} - {1'b0, layer_0_0[4183:4176]};
      top_0[2] = {1'b0,layer_1_0[4191:4184]} - {1'b0, layer_0_0[4191:4184]};
      top_1[0] = {1'b0,layer_1_1[4175:4168]} - {1'b0, layer_0_1[4175:4168]};
      top_1[1] = {1'b0,layer_1_1[4183:4176]} - {1'b0, layer_0_1[4183:4176]};
      top_1[2] = {1'b0,layer_1_1[4191:4184]} - {1'b0, layer_0_1[4191:4184]};
      top_2[0] = {1'b0,layer_1_2[4175:4168]} - {1'b0, layer_0_2[4175:4168]};
      top_2[1] = {1'b0,layer_1_2[4183:4176]} - {1'b0, layer_0_2[4183:4176]};
      top_2[2] = {1'b0,layer_1_2[4191:4184]} - {1'b0, layer_0_2[4191:4184]};
      mid_0[0] = {1'b0,layer_2_0[4175:4168]} - {1'b0, layer_1_0[4175:4168]};
      mid_0[1] = {1'b0,layer_2_0[4183:4176]} - {1'b0, layer_1_0[4183:4176]};
      mid_0[2] = {1'b0,layer_2_0[4191:4184]} - {1'b0, layer_1_0[4191:4184]};
      mid_1[0] = {1'b0,layer_2_1[4175:4168]} - {1'b0, layer_1_1[4175:4168]};
      mid_1[1] = {1'b0,layer_2_1[4183:4176]} - {1'b0, layer_1_1[4183:4176]};
      mid_1[2] = {1'b0,layer_2_1[4191:4184]} - {1'b0, layer_1_1[4191:4184]};
      mid_2[0] = {1'b0,layer_2_2[4175:4168]} - {1'b0, layer_1_2[4175:4168]};
      mid_2[1] = {1'b0,layer_2_2[4183:4176]} - {1'b0, layer_1_2[4183:4176]};
      mid_2[2] = {1'b0,layer_2_2[4191:4184]} - {1'b0, layer_1_2[4191:4184]};
      btm_0[0] = {1'b0,layer_3_0[4175:4168]} - {1'b0, layer_2_0[4175:4168]};
      btm_0[1] = {1'b0,layer_3_0[4183:4176]} - {1'b0, layer_2_0[4183:4176]};
      btm_0[2] = {1'b0,layer_3_0[4191:4184]} - {1'b0, layer_2_0[4191:4184]};
      btm_1[0] = {1'b0,layer_3_1[4175:4168]} - {1'b0, layer_2_1[4175:4168]};
      btm_1[1] = {1'b0,layer_3_1[4183:4176]} - {1'b0, layer_2_1[4183:4176]};
      btm_1[2] = {1'b0,layer_3_1[4191:4184]} - {1'b0, layer_2_1[4191:4184]};
      btm_2[0] = {1'b0,layer_3_2[4175:4168]} - {1'b0, layer_2_2[4175:4168]};
      btm_2[1] = {1'b0,layer_3_2[4183:4176]} - {1'b0, layer_2_2[4183:4176]};
      btm_2[2] = {1'b0,layer_3_2[4191:4184]} - {1'b0, layer_2_2[4191:4184]};
    end
    'd523: begin
      top_0[0] = {1'b0,layer_1_0[4183:4176]} - {1'b0, layer_0_0[4183:4176]};
      top_0[1] = {1'b0,layer_1_0[4191:4184]} - {1'b0, layer_0_0[4191:4184]};
      top_0[2] = {1'b0,layer_1_0[4199:4192]} - {1'b0, layer_0_0[4199:4192]};
      top_1[0] = {1'b0,layer_1_1[4183:4176]} - {1'b0, layer_0_1[4183:4176]};
      top_1[1] = {1'b0,layer_1_1[4191:4184]} - {1'b0, layer_0_1[4191:4184]};
      top_1[2] = {1'b0,layer_1_1[4199:4192]} - {1'b0, layer_0_1[4199:4192]};
      top_2[0] = {1'b0,layer_1_2[4183:4176]} - {1'b0, layer_0_2[4183:4176]};
      top_2[1] = {1'b0,layer_1_2[4191:4184]} - {1'b0, layer_0_2[4191:4184]};
      top_2[2] = {1'b0,layer_1_2[4199:4192]} - {1'b0, layer_0_2[4199:4192]};
      mid_0[0] = {1'b0,layer_2_0[4183:4176]} - {1'b0, layer_1_0[4183:4176]};
      mid_0[1] = {1'b0,layer_2_0[4191:4184]} - {1'b0, layer_1_0[4191:4184]};
      mid_0[2] = {1'b0,layer_2_0[4199:4192]} - {1'b0, layer_1_0[4199:4192]};
      mid_1[0] = {1'b0,layer_2_1[4183:4176]} - {1'b0, layer_1_1[4183:4176]};
      mid_1[1] = {1'b0,layer_2_1[4191:4184]} - {1'b0, layer_1_1[4191:4184]};
      mid_1[2] = {1'b0,layer_2_1[4199:4192]} - {1'b0, layer_1_1[4199:4192]};
      mid_2[0] = {1'b0,layer_2_2[4183:4176]} - {1'b0, layer_1_2[4183:4176]};
      mid_2[1] = {1'b0,layer_2_2[4191:4184]} - {1'b0, layer_1_2[4191:4184]};
      mid_2[2] = {1'b0,layer_2_2[4199:4192]} - {1'b0, layer_1_2[4199:4192]};
      btm_0[0] = {1'b0,layer_3_0[4183:4176]} - {1'b0, layer_2_0[4183:4176]};
      btm_0[1] = {1'b0,layer_3_0[4191:4184]} - {1'b0, layer_2_0[4191:4184]};
      btm_0[2] = {1'b0,layer_3_0[4199:4192]} - {1'b0, layer_2_0[4199:4192]};
      btm_1[0] = {1'b0,layer_3_1[4183:4176]} - {1'b0, layer_2_1[4183:4176]};
      btm_1[1] = {1'b0,layer_3_1[4191:4184]} - {1'b0, layer_2_1[4191:4184]};
      btm_1[2] = {1'b0,layer_3_1[4199:4192]} - {1'b0, layer_2_1[4199:4192]};
      btm_2[0] = {1'b0,layer_3_2[4183:4176]} - {1'b0, layer_2_2[4183:4176]};
      btm_2[1] = {1'b0,layer_3_2[4191:4184]} - {1'b0, layer_2_2[4191:4184]};
      btm_2[2] = {1'b0,layer_3_2[4199:4192]} - {1'b0, layer_2_2[4199:4192]};
    end
    'd524: begin
      top_0[0] = {1'b0,layer_1_0[4191:4184]} - {1'b0, layer_0_0[4191:4184]};
      top_0[1] = {1'b0,layer_1_0[4199:4192]} - {1'b0, layer_0_0[4199:4192]};
      top_0[2] = {1'b0,layer_1_0[4207:4200]} - {1'b0, layer_0_0[4207:4200]};
      top_1[0] = {1'b0,layer_1_1[4191:4184]} - {1'b0, layer_0_1[4191:4184]};
      top_1[1] = {1'b0,layer_1_1[4199:4192]} - {1'b0, layer_0_1[4199:4192]};
      top_1[2] = {1'b0,layer_1_1[4207:4200]} - {1'b0, layer_0_1[4207:4200]};
      top_2[0] = {1'b0,layer_1_2[4191:4184]} - {1'b0, layer_0_2[4191:4184]};
      top_2[1] = {1'b0,layer_1_2[4199:4192]} - {1'b0, layer_0_2[4199:4192]};
      top_2[2] = {1'b0,layer_1_2[4207:4200]} - {1'b0, layer_0_2[4207:4200]};
      mid_0[0] = {1'b0,layer_2_0[4191:4184]} - {1'b0, layer_1_0[4191:4184]};
      mid_0[1] = {1'b0,layer_2_0[4199:4192]} - {1'b0, layer_1_0[4199:4192]};
      mid_0[2] = {1'b0,layer_2_0[4207:4200]} - {1'b0, layer_1_0[4207:4200]};
      mid_1[0] = {1'b0,layer_2_1[4191:4184]} - {1'b0, layer_1_1[4191:4184]};
      mid_1[1] = {1'b0,layer_2_1[4199:4192]} - {1'b0, layer_1_1[4199:4192]};
      mid_1[2] = {1'b0,layer_2_1[4207:4200]} - {1'b0, layer_1_1[4207:4200]};
      mid_2[0] = {1'b0,layer_2_2[4191:4184]} - {1'b0, layer_1_2[4191:4184]};
      mid_2[1] = {1'b0,layer_2_2[4199:4192]} - {1'b0, layer_1_2[4199:4192]};
      mid_2[2] = {1'b0,layer_2_2[4207:4200]} - {1'b0, layer_1_2[4207:4200]};
      btm_0[0] = {1'b0,layer_3_0[4191:4184]} - {1'b0, layer_2_0[4191:4184]};
      btm_0[1] = {1'b0,layer_3_0[4199:4192]} - {1'b0, layer_2_0[4199:4192]};
      btm_0[2] = {1'b0,layer_3_0[4207:4200]} - {1'b0, layer_2_0[4207:4200]};
      btm_1[0] = {1'b0,layer_3_1[4191:4184]} - {1'b0, layer_2_1[4191:4184]};
      btm_1[1] = {1'b0,layer_3_1[4199:4192]} - {1'b0, layer_2_1[4199:4192]};
      btm_1[2] = {1'b0,layer_3_1[4207:4200]} - {1'b0, layer_2_1[4207:4200]};
      btm_2[0] = {1'b0,layer_3_2[4191:4184]} - {1'b0, layer_2_2[4191:4184]};
      btm_2[1] = {1'b0,layer_3_2[4199:4192]} - {1'b0, layer_2_2[4199:4192]};
      btm_2[2] = {1'b0,layer_3_2[4207:4200]} - {1'b0, layer_2_2[4207:4200]};
    end
    'd525: begin
      top_0[0] = {1'b0,layer_1_0[4199:4192]} - {1'b0, layer_0_0[4199:4192]};
      top_0[1] = {1'b0,layer_1_0[4207:4200]} - {1'b0, layer_0_0[4207:4200]};
      top_0[2] = {1'b0,layer_1_0[4215:4208]} - {1'b0, layer_0_0[4215:4208]};
      top_1[0] = {1'b0,layer_1_1[4199:4192]} - {1'b0, layer_0_1[4199:4192]};
      top_1[1] = {1'b0,layer_1_1[4207:4200]} - {1'b0, layer_0_1[4207:4200]};
      top_1[2] = {1'b0,layer_1_1[4215:4208]} - {1'b0, layer_0_1[4215:4208]};
      top_2[0] = {1'b0,layer_1_2[4199:4192]} - {1'b0, layer_0_2[4199:4192]};
      top_2[1] = {1'b0,layer_1_2[4207:4200]} - {1'b0, layer_0_2[4207:4200]};
      top_2[2] = {1'b0,layer_1_2[4215:4208]} - {1'b0, layer_0_2[4215:4208]};
      mid_0[0] = {1'b0,layer_2_0[4199:4192]} - {1'b0, layer_1_0[4199:4192]};
      mid_0[1] = {1'b0,layer_2_0[4207:4200]} - {1'b0, layer_1_0[4207:4200]};
      mid_0[2] = {1'b0,layer_2_0[4215:4208]} - {1'b0, layer_1_0[4215:4208]};
      mid_1[0] = {1'b0,layer_2_1[4199:4192]} - {1'b0, layer_1_1[4199:4192]};
      mid_1[1] = {1'b0,layer_2_1[4207:4200]} - {1'b0, layer_1_1[4207:4200]};
      mid_1[2] = {1'b0,layer_2_1[4215:4208]} - {1'b0, layer_1_1[4215:4208]};
      mid_2[0] = {1'b0,layer_2_2[4199:4192]} - {1'b0, layer_1_2[4199:4192]};
      mid_2[1] = {1'b0,layer_2_2[4207:4200]} - {1'b0, layer_1_2[4207:4200]};
      mid_2[2] = {1'b0,layer_2_2[4215:4208]} - {1'b0, layer_1_2[4215:4208]};
      btm_0[0] = {1'b0,layer_3_0[4199:4192]} - {1'b0, layer_2_0[4199:4192]};
      btm_0[1] = {1'b0,layer_3_0[4207:4200]} - {1'b0, layer_2_0[4207:4200]};
      btm_0[2] = {1'b0,layer_3_0[4215:4208]} - {1'b0, layer_2_0[4215:4208]};
      btm_1[0] = {1'b0,layer_3_1[4199:4192]} - {1'b0, layer_2_1[4199:4192]};
      btm_1[1] = {1'b0,layer_3_1[4207:4200]} - {1'b0, layer_2_1[4207:4200]};
      btm_1[2] = {1'b0,layer_3_1[4215:4208]} - {1'b0, layer_2_1[4215:4208]};
      btm_2[0] = {1'b0,layer_3_2[4199:4192]} - {1'b0, layer_2_2[4199:4192]};
      btm_2[1] = {1'b0,layer_3_2[4207:4200]} - {1'b0, layer_2_2[4207:4200]};
      btm_2[2] = {1'b0,layer_3_2[4215:4208]} - {1'b0, layer_2_2[4215:4208]};
    end
    'd526: begin
      top_0[0] = {1'b0,layer_1_0[4207:4200]} - {1'b0, layer_0_0[4207:4200]};
      top_0[1] = {1'b0,layer_1_0[4215:4208]} - {1'b0, layer_0_0[4215:4208]};
      top_0[2] = {1'b0,layer_1_0[4223:4216]} - {1'b0, layer_0_0[4223:4216]};
      top_1[0] = {1'b0,layer_1_1[4207:4200]} - {1'b0, layer_0_1[4207:4200]};
      top_1[1] = {1'b0,layer_1_1[4215:4208]} - {1'b0, layer_0_1[4215:4208]};
      top_1[2] = {1'b0,layer_1_1[4223:4216]} - {1'b0, layer_0_1[4223:4216]};
      top_2[0] = {1'b0,layer_1_2[4207:4200]} - {1'b0, layer_0_2[4207:4200]};
      top_2[1] = {1'b0,layer_1_2[4215:4208]} - {1'b0, layer_0_2[4215:4208]};
      top_2[2] = {1'b0,layer_1_2[4223:4216]} - {1'b0, layer_0_2[4223:4216]};
      mid_0[0] = {1'b0,layer_2_0[4207:4200]} - {1'b0, layer_1_0[4207:4200]};
      mid_0[1] = {1'b0,layer_2_0[4215:4208]} - {1'b0, layer_1_0[4215:4208]};
      mid_0[2] = {1'b0,layer_2_0[4223:4216]} - {1'b0, layer_1_0[4223:4216]};
      mid_1[0] = {1'b0,layer_2_1[4207:4200]} - {1'b0, layer_1_1[4207:4200]};
      mid_1[1] = {1'b0,layer_2_1[4215:4208]} - {1'b0, layer_1_1[4215:4208]};
      mid_1[2] = {1'b0,layer_2_1[4223:4216]} - {1'b0, layer_1_1[4223:4216]};
      mid_2[0] = {1'b0,layer_2_2[4207:4200]} - {1'b0, layer_1_2[4207:4200]};
      mid_2[1] = {1'b0,layer_2_2[4215:4208]} - {1'b0, layer_1_2[4215:4208]};
      mid_2[2] = {1'b0,layer_2_2[4223:4216]} - {1'b0, layer_1_2[4223:4216]};
      btm_0[0] = {1'b0,layer_3_0[4207:4200]} - {1'b0, layer_2_0[4207:4200]};
      btm_0[1] = {1'b0,layer_3_0[4215:4208]} - {1'b0, layer_2_0[4215:4208]};
      btm_0[2] = {1'b0,layer_3_0[4223:4216]} - {1'b0, layer_2_0[4223:4216]};
      btm_1[0] = {1'b0,layer_3_1[4207:4200]} - {1'b0, layer_2_1[4207:4200]};
      btm_1[1] = {1'b0,layer_3_1[4215:4208]} - {1'b0, layer_2_1[4215:4208]};
      btm_1[2] = {1'b0,layer_3_1[4223:4216]} - {1'b0, layer_2_1[4223:4216]};
      btm_2[0] = {1'b0,layer_3_2[4207:4200]} - {1'b0, layer_2_2[4207:4200]};
      btm_2[1] = {1'b0,layer_3_2[4215:4208]} - {1'b0, layer_2_2[4215:4208]};
      btm_2[2] = {1'b0,layer_3_2[4223:4216]} - {1'b0, layer_2_2[4223:4216]};
    end
    'd527: begin
      top_0[0] = {1'b0,layer_1_0[4215:4208]} - {1'b0, layer_0_0[4215:4208]};
      top_0[1] = {1'b0,layer_1_0[4223:4216]} - {1'b0, layer_0_0[4223:4216]};
      top_0[2] = {1'b0,layer_1_0[4231:4224]} - {1'b0, layer_0_0[4231:4224]};
      top_1[0] = {1'b0,layer_1_1[4215:4208]} - {1'b0, layer_0_1[4215:4208]};
      top_1[1] = {1'b0,layer_1_1[4223:4216]} - {1'b0, layer_0_1[4223:4216]};
      top_1[2] = {1'b0,layer_1_1[4231:4224]} - {1'b0, layer_0_1[4231:4224]};
      top_2[0] = {1'b0,layer_1_2[4215:4208]} - {1'b0, layer_0_2[4215:4208]};
      top_2[1] = {1'b0,layer_1_2[4223:4216]} - {1'b0, layer_0_2[4223:4216]};
      top_2[2] = {1'b0,layer_1_2[4231:4224]} - {1'b0, layer_0_2[4231:4224]};
      mid_0[0] = {1'b0,layer_2_0[4215:4208]} - {1'b0, layer_1_0[4215:4208]};
      mid_0[1] = {1'b0,layer_2_0[4223:4216]} - {1'b0, layer_1_0[4223:4216]};
      mid_0[2] = {1'b0,layer_2_0[4231:4224]} - {1'b0, layer_1_0[4231:4224]};
      mid_1[0] = {1'b0,layer_2_1[4215:4208]} - {1'b0, layer_1_1[4215:4208]};
      mid_1[1] = {1'b0,layer_2_1[4223:4216]} - {1'b0, layer_1_1[4223:4216]};
      mid_1[2] = {1'b0,layer_2_1[4231:4224]} - {1'b0, layer_1_1[4231:4224]};
      mid_2[0] = {1'b0,layer_2_2[4215:4208]} - {1'b0, layer_1_2[4215:4208]};
      mid_2[1] = {1'b0,layer_2_2[4223:4216]} - {1'b0, layer_1_2[4223:4216]};
      mid_2[2] = {1'b0,layer_2_2[4231:4224]} - {1'b0, layer_1_2[4231:4224]};
      btm_0[0] = {1'b0,layer_3_0[4215:4208]} - {1'b0, layer_2_0[4215:4208]};
      btm_0[1] = {1'b0,layer_3_0[4223:4216]} - {1'b0, layer_2_0[4223:4216]};
      btm_0[2] = {1'b0,layer_3_0[4231:4224]} - {1'b0, layer_2_0[4231:4224]};
      btm_1[0] = {1'b0,layer_3_1[4215:4208]} - {1'b0, layer_2_1[4215:4208]};
      btm_1[1] = {1'b0,layer_3_1[4223:4216]} - {1'b0, layer_2_1[4223:4216]};
      btm_1[2] = {1'b0,layer_3_1[4231:4224]} - {1'b0, layer_2_1[4231:4224]};
      btm_2[0] = {1'b0,layer_3_2[4215:4208]} - {1'b0, layer_2_2[4215:4208]};
      btm_2[1] = {1'b0,layer_3_2[4223:4216]} - {1'b0, layer_2_2[4223:4216]};
      btm_2[2] = {1'b0,layer_3_2[4231:4224]} - {1'b0, layer_2_2[4231:4224]};
    end
    'd528: begin
      top_0[0] = {1'b0,layer_1_0[4223:4216]} - {1'b0, layer_0_0[4223:4216]};
      top_0[1] = {1'b0,layer_1_0[4231:4224]} - {1'b0, layer_0_0[4231:4224]};
      top_0[2] = {1'b0,layer_1_0[4239:4232]} - {1'b0, layer_0_0[4239:4232]};
      top_1[0] = {1'b0,layer_1_1[4223:4216]} - {1'b0, layer_0_1[4223:4216]};
      top_1[1] = {1'b0,layer_1_1[4231:4224]} - {1'b0, layer_0_1[4231:4224]};
      top_1[2] = {1'b0,layer_1_1[4239:4232]} - {1'b0, layer_0_1[4239:4232]};
      top_2[0] = {1'b0,layer_1_2[4223:4216]} - {1'b0, layer_0_2[4223:4216]};
      top_2[1] = {1'b0,layer_1_2[4231:4224]} - {1'b0, layer_0_2[4231:4224]};
      top_2[2] = {1'b0,layer_1_2[4239:4232]} - {1'b0, layer_0_2[4239:4232]};
      mid_0[0] = {1'b0,layer_2_0[4223:4216]} - {1'b0, layer_1_0[4223:4216]};
      mid_0[1] = {1'b0,layer_2_0[4231:4224]} - {1'b0, layer_1_0[4231:4224]};
      mid_0[2] = {1'b0,layer_2_0[4239:4232]} - {1'b0, layer_1_0[4239:4232]};
      mid_1[0] = {1'b0,layer_2_1[4223:4216]} - {1'b0, layer_1_1[4223:4216]};
      mid_1[1] = {1'b0,layer_2_1[4231:4224]} - {1'b0, layer_1_1[4231:4224]};
      mid_1[2] = {1'b0,layer_2_1[4239:4232]} - {1'b0, layer_1_1[4239:4232]};
      mid_2[0] = {1'b0,layer_2_2[4223:4216]} - {1'b0, layer_1_2[4223:4216]};
      mid_2[1] = {1'b0,layer_2_2[4231:4224]} - {1'b0, layer_1_2[4231:4224]};
      mid_2[2] = {1'b0,layer_2_2[4239:4232]} - {1'b0, layer_1_2[4239:4232]};
      btm_0[0] = {1'b0,layer_3_0[4223:4216]} - {1'b0, layer_2_0[4223:4216]};
      btm_0[1] = {1'b0,layer_3_0[4231:4224]} - {1'b0, layer_2_0[4231:4224]};
      btm_0[2] = {1'b0,layer_3_0[4239:4232]} - {1'b0, layer_2_0[4239:4232]};
      btm_1[0] = {1'b0,layer_3_1[4223:4216]} - {1'b0, layer_2_1[4223:4216]};
      btm_1[1] = {1'b0,layer_3_1[4231:4224]} - {1'b0, layer_2_1[4231:4224]};
      btm_1[2] = {1'b0,layer_3_1[4239:4232]} - {1'b0, layer_2_1[4239:4232]};
      btm_2[0] = {1'b0,layer_3_2[4223:4216]} - {1'b0, layer_2_2[4223:4216]};
      btm_2[1] = {1'b0,layer_3_2[4231:4224]} - {1'b0, layer_2_2[4231:4224]};
      btm_2[2] = {1'b0,layer_3_2[4239:4232]} - {1'b0, layer_2_2[4239:4232]};
    end
    'd529: begin
      top_0[0] = {1'b0,layer_1_0[4231:4224]} - {1'b0, layer_0_0[4231:4224]};
      top_0[1] = {1'b0,layer_1_0[4239:4232]} - {1'b0, layer_0_0[4239:4232]};
      top_0[2] = {1'b0,layer_1_0[4247:4240]} - {1'b0, layer_0_0[4247:4240]};
      top_1[0] = {1'b0,layer_1_1[4231:4224]} - {1'b0, layer_0_1[4231:4224]};
      top_1[1] = {1'b0,layer_1_1[4239:4232]} - {1'b0, layer_0_1[4239:4232]};
      top_1[2] = {1'b0,layer_1_1[4247:4240]} - {1'b0, layer_0_1[4247:4240]};
      top_2[0] = {1'b0,layer_1_2[4231:4224]} - {1'b0, layer_0_2[4231:4224]};
      top_2[1] = {1'b0,layer_1_2[4239:4232]} - {1'b0, layer_0_2[4239:4232]};
      top_2[2] = {1'b0,layer_1_2[4247:4240]} - {1'b0, layer_0_2[4247:4240]};
      mid_0[0] = {1'b0,layer_2_0[4231:4224]} - {1'b0, layer_1_0[4231:4224]};
      mid_0[1] = {1'b0,layer_2_0[4239:4232]} - {1'b0, layer_1_0[4239:4232]};
      mid_0[2] = {1'b0,layer_2_0[4247:4240]} - {1'b0, layer_1_0[4247:4240]};
      mid_1[0] = {1'b0,layer_2_1[4231:4224]} - {1'b0, layer_1_1[4231:4224]};
      mid_1[1] = {1'b0,layer_2_1[4239:4232]} - {1'b0, layer_1_1[4239:4232]};
      mid_1[2] = {1'b0,layer_2_1[4247:4240]} - {1'b0, layer_1_1[4247:4240]};
      mid_2[0] = {1'b0,layer_2_2[4231:4224]} - {1'b0, layer_1_2[4231:4224]};
      mid_2[1] = {1'b0,layer_2_2[4239:4232]} - {1'b0, layer_1_2[4239:4232]};
      mid_2[2] = {1'b0,layer_2_2[4247:4240]} - {1'b0, layer_1_2[4247:4240]};
      btm_0[0] = {1'b0,layer_3_0[4231:4224]} - {1'b0, layer_2_0[4231:4224]};
      btm_0[1] = {1'b0,layer_3_0[4239:4232]} - {1'b0, layer_2_0[4239:4232]};
      btm_0[2] = {1'b0,layer_3_0[4247:4240]} - {1'b0, layer_2_0[4247:4240]};
      btm_1[0] = {1'b0,layer_3_1[4231:4224]} - {1'b0, layer_2_1[4231:4224]};
      btm_1[1] = {1'b0,layer_3_1[4239:4232]} - {1'b0, layer_2_1[4239:4232]};
      btm_1[2] = {1'b0,layer_3_1[4247:4240]} - {1'b0, layer_2_1[4247:4240]};
      btm_2[0] = {1'b0,layer_3_2[4231:4224]} - {1'b0, layer_2_2[4231:4224]};
      btm_2[1] = {1'b0,layer_3_2[4239:4232]} - {1'b0, layer_2_2[4239:4232]};
      btm_2[2] = {1'b0,layer_3_2[4247:4240]} - {1'b0, layer_2_2[4247:4240]};
    end
    'd530: begin
      top_0[0] = {1'b0,layer_1_0[4239:4232]} - {1'b0, layer_0_0[4239:4232]};
      top_0[1] = {1'b0,layer_1_0[4247:4240]} - {1'b0, layer_0_0[4247:4240]};
      top_0[2] = {1'b0,layer_1_0[4255:4248]} - {1'b0, layer_0_0[4255:4248]};
      top_1[0] = {1'b0,layer_1_1[4239:4232]} - {1'b0, layer_0_1[4239:4232]};
      top_1[1] = {1'b0,layer_1_1[4247:4240]} - {1'b0, layer_0_1[4247:4240]};
      top_1[2] = {1'b0,layer_1_1[4255:4248]} - {1'b0, layer_0_1[4255:4248]};
      top_2[0] = {1'b0,layer_1_2[4239:4232]} - {1'b0, layer_0_2[4239:4232]};
      top_2[1] = {1'b0,layer_1_2[4247:4240]} - {1'b0, layer_0_2[4247:4240]};
      top_2[2] = {1'b0,layer_1_2[4255:4248]} - {1'b0, layer_0_2[4255:4248]};
      mid_0[0] = {1'b0,layer_2_0[4239:4232]} - {1'b0, layer_1_0[4239:4232]};
      mid_0[1] = {1'b0,layer_2_0[4247:4240]} - {1'b0, layer_1_0[4247:4240]};
      mid_0[2] = {1'b0,layer_2_0[4255:4248]} - {1'b0, layer_1_0[4255:4248]};
      mid_1[0] = {1'b0,layer_2_1[4239:4232]} - {1'b0, layer_1_1[4239:4232]};
      mid_1[1] = {1'b0,layer_2_1[4247:4240]} - {1'b0, layer_1_1[4247:4240]};
      mid_1[2] = {1'b0,layer_2_1[4255:4248]} - {1'b0, layer_1_1[4255:4248]};
      mid_2[0] = {1'b0,layer_2_2[4239:4232]} - {1'b0, layer_1_2[4239:4232]};
      mid_2[1] = {1'b0,layer_2_2[4247:4240]} - {1'b0, layer_1_2[4247:4240]};
      mid_2[2] = {1'b0,layer_2_2[4255:4248]} - {1'b0, layer_1_2[4255:4248]};
      btm_0[0] = {1'b0,layer_3_0[4239:4232]} - {1'b0, layer_2_0[4239:4232]};
      btm_0[1] = {1'b0,layer_3_0[4247:4240]} - {1'b0, layer_2_0[4247:4240]};
      btm_0[2] = {1'b0,layer_3_0[4255:4248]} - {1'b0, layer_2_0[4255:4248]};
      btm_1[0] = {1'b0,layer_3_1[4239:4232]} - {1'b0, layer_2_1[4239:4232]};
      btm_1[1] = {1'b0,layer_3_1[4247:4240]} - {1'b0, layer_2_1[4247:4240]};
      btm_1[2] = {1'b0,layer_3_1[4255:4248]} - {1'b0, layer_2_1[4255:4248]};
      btm_2[0] = {1'b0,layer_3_2[4239:4232]} - {1'b0, layer_2_2[4239:4232]};
      btm_2[1] = {1'b0,layer_3_2[4247:4240]} - {1'b0, layer_2_2[4247:4240]};
      btm_2[2] = {1'b0,layer_3_2[4255:4248]} - {1'b0, layer_2_2[4255:4248]};
    end
    'd531: begin
      top_0[0] = {1'b0,layer_1_0[4247:4240]} - {1'b0, layer_0_0[4247:4240]};
      top_0[1] = {1'b0,layer_1_0[4255:4248]} - {1'b0, layer_0_0[4255:4248]};
      top_0[2] = {1'b0,layer_1_0[4263:4256]} - {1'b0, layer_0_0[4263:4256]};
      top_1[0] = {1'b0,layer_1_1[4247:4240]} - {1'b0, layer_0_1[4247:4240]};
      top_1[1] = {1'b0,layer_1_1[4255:4248]} - {1'b0, layer_0_1[4255:4248]};
      top_1[2] = {1'b0,layer_1_1[4263:4256]} - {1'b0, layer_0_1[4263:4256]};
      top_2[0] = {1'b0,layer_1_2[4247:4240]} - {1'b0, layer_0_2[4247:4240]};
      top_2[1] = {1'b0,layer_1_2[4255:4248]} - {1'b0, layer_0_2[4255:4248]};
      top_2[2] = {1'b0,layer_1_2[4263:4256]} - {1'b0, layer_0_2[4263:4256]};
      mid_0[0] = {1'b0,layer_2_0[4247:4240]} - {1'b0, layer_1_0[4247:4240]};
      mid_0[1] = {1'b0,layer_2_0[4255:4248]} - {1'b0, layer_1_0[4255:4248]};
      mid_0[2] = {1'b0,layer_2_0[4263:4256]} - {1'b0, layer_1_0[4263:4256]};
      mid_1[0] = {1'b0,layer_2_1[4247:4240]} - {1'b0, layer_1_1[4247:4240]};
      mid_1[1] = {1'b0,layer_2_1[4255:4248]} - {1'b0, layer_1_1[4255:4248]};
      mid_1[2] = {1'b0,layer_2_1[4263:4256]} - {1'b0, layer_1_1[4263:4256]};
      mid_2[0] = {1'b0,layer_2_2[4247:4240]} - {1'b0, layer_1_2[4247:4240]};
      mid_2[1] = {1'b0,layer_2_2[4255:4248]} - {1'b0, layer_1_2[4255:4248]};
      mid_2[2] = {1'b0,layer_2_2[4263:4256]} - {1'b0, layer_1_2[4263:4256]};
      btm_0[0] = {1'b0,layer_3_0[4247:4240]} - {1'b0, layer_2_0[4247:4240]};
      btm_0[1] = {1'b0,layer_3_0[4255:4248]} - {1'b0, layer_2_0[4255:4248]};
      btm_0[2] = {1'b0,layer_3_0[4263:4256]} - {1'b0, layer_2_0[4263:4256]};
      btm_1[0] = {1'b0,layer_3_1[4247:4240]} - {1'b0, layer_2_1[4247:4240]};
      btm_1[1] = {1'b0,layer_3_1[4255:4248]} - {1'b0, layer_2_1[4255:4248]};
      btm_1[2] = {1'b0,layer_3_1[4263:4256]} - {1'b0, layer_2_1[4263:4256]};
      btm_2[0] = {1'b0,layer_3_2[4247:4240]} - {1'b0, layer_2_2[4247:4240]};
      btm_2[1] = {1'b0,layer_3_2[4255:4248]} - {1'b0, layer_2_2[4255:4248]};
      btm_2[2] = {1'b0,layer_3_2[4263:4256]} - {1'b0, layer_2_2[4263:4256]};
    end
    'd532: begin
      top_0[0] = {1'b0,layer_1_0[4255:4248]} - {1'b0, layer_0_0[4255:4248]};
      top_0[1] = {1'b0,layer_1_0[4263:4256]} - {1'b0, layer_0_0[4263:4256]};
      top_0[2] = {1'b0,layer_1_0[4271:4264]} - {1'b0, layer_0_0[4271:4264]};
      top_1[0] = {1'b0,layer_1_1[4255:4248]} - {1'b0, layer_0_1[4255:4248]};
      top_1[1] = {1'b0,layer_1_1[4263:4256]} - {1'b0, layer_0_1[4263:4256]};
      top_1[2] = {1'b0,layer_1_1[4271:4264]} - {1'b0, layer_0_1[4271:4264]};
      top_2[0] = {1'b0,layer_1_2[4255:4248]} - {1'b0, layer_0_2[4255:4248]};
      top_2[1] = {1'b0,layer_1_2[4263:4256]} - {1'b0, layer_0_2[4263:4256]};
      top_2[2] = {1'b0,layer_1_2[4271:4264]} - {1'b0, layer_0_2[4271:4264]};
      mid_0[0] = {1'b0,layer_2_0[4255:4248]} - {1'b0, layer_1_0[4255:4248]};
      mid_0[1] = {1'b0,layer_2_0[4263:4256]} - {1'b0, layer_1_0[4263:4256]};
      mid_0[2] = {1'b0,layer_2_0[4271:4264]} - {1'b0, layer_1_0[4271:4264]};
      mid_1[0] = {1'b0,layer_2_1[4255:4248]} - {1'b0, layer_1_1[4255:4248]};
      mid_1[1] = {1'b0,layer_2_1[4263:4256]} - {1'b0, layer_1_1[4263:4256]};
      mid_1[2] = {1'b0,layer_2_1[4271:4264]} - {1'b0, layer_1_1[4271:4264]};
      mid_2[0] = {1'b0,layer_2_2[4255:4248]} - {1'b0, layer_1_2[4255:4248]};
      mid_2[1] = {1'b0,layer_2_2[4263:4256]} - {1'b0, layer_1_2[4263:4256]};
      mid_2[2] = {1'b0,layer_2_2[4271:4264]} - {1'b0, layer_1_2[4271:4264]};
      btm_0[0] = {1'b0,layer_3_0[4255:4248]} - {1'b0, layer_2_0[4255:4248]};
      btm_0[1] = {1'b0,layer_3_0[4263:4256]} - {1'b0, layer_2_0[4263:4256]};
      btm_0[2] = {1'b0,layer_3_0[4271:4264]} - {1'b0, layer_2_0[4271:4264]};
      btm_1[0] = {1'b0,layer_3_1[4255:4248]} - {1'b0, layer_2_1[4255:4248]};
      btm_1[1] = {1'b0,layer_3_1[4263:4256]} - {1'b0, layer_2_1[4263:4256]};
      btm_1[2] = {1'b0,layer_3_1[4271:4264]} - {1'b0, layer_2_1[4271:4264]};
      btm_2[0] = {1'b0,layer_3_2[4255:4248]} - {1'b0, layer_2_2[4255:4248]};
      btm_2[1] = {1'b0,layer_3_2[4263:4256]} - {1'b0, layer_2_2[4263:4256]};
      btm_2[2] = {1'b0,layer_3_2[4271:4264]} - {1'b0, layer_2_2[4271:4264]};
    end
    'd533: begin
      top_0[0] = {1'b0,layer_1_0[4263:4256]} - {1'b0, layer_0_0[4263:4256]};
      top_0[1] = {1'b0,layer_1_0[4271:4264]} - {1'b0, layer_0_0[4271:4264]};
      top_0[2] = {1'b0,layer_1_0[4279:4272]} - {1'b0, layer_0_0[4279:4272]};
      top_1[0] = {1'b0,layer_1_1[4263:4256]} - {1'b0, layer_0_1[4263:4256]};
      top_1[1] = {1'b0,layer_1_1[4271:4264]} - {1'b0, layer_0_1[4271:4264]};
      top_1[2] = {1'b0,layer_1_1[4279:4272]} - {1'b0, layer_0_1[4279:4272]};
      top_2[0] = {1'b0,layer_1_2[4263:4256]} - {1'b0, layer_0_2[4263:4256]};
      top_2[1] = {1'b0,layer_1_2[4271:4264]} - {1'b0, layer_0_2[4271:4264]};
      top_2[2] = {1'b0,layer_1_2[4279:4272]} - {1'b0, layer_0_2[4279:4272]};
      mid_0[0] = {1'b0,layer_2_0[4263:4256]} - {1'b0, layer_1_0[4263:4256]};
      mid_0[1] = {1'b0,layer_2_0[4271:4264]} - {1'b0, layer_1_0[4271:4264]};
      mid_0[2] = {1'b0,layer_2_0[4279:4272]} - {1'b0, layer_1_0[4279:4272]};
      mid_1[0] = {1'b0,layer_2_1[4263:4256]} - {1'b0, layer_1_1[4263:4256]};
      mid_1[1] = {1'b0,layer_2_1[4271:4264]} - {1'b0, layer_1_1[4271:4264]};
      mid_1[2] = {1'b0,layer_2_1[4279:4272]} - {1'b0, layer_1_1[4279:4272]};
      mid_2[0] = {1'b0,layer_2_2[4263:4256]} - {1'b0, layer_1_2[4263:4256]};
      mid_2[1] = {1'b0,layer_2_2[4271:4264]} - {1'b0, layer_1_2[4271:4264]};
      mid_2[2] = {1'b0,layer_2_2[4279:4272]} - {1'b0, layer_1_2[4279:4272]};
      btm_0[0] = {1'b0,layer_3_0[4263:4256]} - {1'b0, layer_2_0[4263:4256]};
      btm_0[1] = {1'b0,layer_3_0[4271:4264]} - {1'b0, layer_2_0[4271:4264]};
      btm_0[2] = {1'b0,layer_3_0[4279:4272]} - {1'b0, layer_2_0[4279:4272]};
      btm_1[0] = {1'b0,layer_3_1[4263:4256]} - {1'b0, layer_2_1[4263:4256]};
      btm_1[1] = {1'b0,layer_3_1[4271:4264]} - {1'b0, layer_2_1[4271:4264]};
      btm_1[2] = {1'b0,layer_3_1[4279:4272]} - {1'b0, layer_2_1[4279:4272]};
      btm_2[0] = {1'b0,layer_3_2[4263:4256]} - {1'b0, layer_2_2[4263:4256]};
      btm_2[1] = {1'b0,layer_3_2[4271:4264]} - {1'b0, layer_2_2[4271:4264]};
      btm_2[2] = {1'b0,layer_3_2[4279:4272]} - {1'b0, layer_2_2[4279:4272]};
    end
    'd534: begin
      top_0[0] = {1'b0,layer_1_0[4271:4264]} - {1'b0, layer_0_0[4271:4264]};
      top_0[1] = {1'b0,layer_1_0[4279:4272]} - {1'b0, layer_0_0[4279:4272]};
      top_0[2] = {1'b0,layer_1_0[4287:4280]} - {1'b0, layer_0_0[4287:4280]};
      top_1[0] = {1'b0,layer_1_1[4271:4264]} - {1'b0, layer_0_1[4271:4264]};
      top_1[1] = {1'b0,layer_1_1[4279:4272]} - {1'b0, layer_0_1[4279:4272]};
      top_1[2] = {1'b0,layer_1_1[4287:4280]} - {1'b0, layer_0_1[4287:4280]};
      top_2[0] = {1'b0,layer_1_2[4271:4264]} - {1'b0, layer_0_2[4271:4264]};
      top_2[1] = {1'b0,layer_1_2[4279:4272]} - {1'b0, layer_0_2[4279:4272]};
      top_2[2] = {1'b0,layer_1_2[4287:4280]} - {1'b0, layer_0_2[4287:4280]};
      mid_0[0] = {1'b0,layer_2_0[4271:4264]} - {1'b0, layer_1_0[4271:4264]};
      mid_0[1] = {1'b0,layer_2_0[4279:4272]} - {1'b0, layer_1_0[4279:4272]};
      mid_0[2] = {1'b0,layer_2_0[4287:4280]} - {1'b0, layer_1_0[4287:4280]};
      mid_1[0] = {1'b0,layer_2_1[4271:4264]} - {1'b0, layer_1_1[4271:4264]};
      mid_1[1] = {1'b0,layer_2_1[4279:4272]} - {1'b0, layer_1_1[4279:4272]};
      mid_1[2] = {1'b0,layer_2_1[4287:4280]} - {1'b0, layer_1_1[4287:4280]};
      mid_2[0] = {1'b0,layer_2_2[4271:4264]} - {1'b0, layer_1_2[4271:4264]};
      mid_2[1] = {1'b0,layer_2_2[4279:4272]} - {1'b0, layer_1_2[4279:4272]};
      mid_2[2] = {1'b0,layer_2_2[4287:4280]} - {1'b0, layer_1_2[4287:4280]};
      btm_0[0] = {1'b0,layer_3_0[4271:4264]} - {1'b0, layer_2_0[4271:4264]};
      btm_0[1] = {1'b0,layer_3_0[4279:4272]} - {1'b0, layer_2_0[4279:4272]};
      btm_0[2] = {1'b0,layer_3_0[4287:4280]} - {1'b0, layer_2_0[4287:4280]};
      btm_1[0] = {1'b0,layer_3_1[4271:4264]} - {1'b0, layer_2_1[4271:4264]};
      btm_1[1] = {1'b0,layer_3_1[4279:4272]} - {1'b0, layer_2_1[4279:4272]};
      btm_1[2] = {1'b0,layer_3_1[4287:4280]} - {1'b0, layer_2_1[4287:4280]};
      btm_2[0] = {1'b0,layer_3_2[4271:4264]} - {1'b0, layer_2_2[4271:4264]};
      btm_2[1] = {1'b0,layer_3_2[4279:4272]} - {1'b0, layer_2_2[4279:4272]};
      btm_2[2] = {1'b0,layer_3_2[4287:4280]} - {1'b0, layer_2_2[4287:4280]};
    end
    'd535: begin
      top_0[0] = {1'b0,layer_1_0[4279:4272]} - {1'b0, layer_0_0[4279:4272]};
      top_0[1] = {1'b0,layer_1_0[4287:4280]} - {1'b0, layer_0_0[4287:4280]};
      top_0[2] = {1'b0,layer_1_0[4295:4288]} - {1'b0, layer_0_0[4295:4288]};
      top_1[0] = {1'b0,layer_1_1[4279:4272]} - {1'b0, layer_0_1[4279:4272]};
      top_1[1] = {1'b0,layer_1_1[4287:4280]} - {1'b0, layer_0_1[4287:4280]};
      top_1[2] = {1'b0,layer_1_1[4295:4288]} - {1'b0, layer_0_1[4295:4288]};
      top_2[0] = {1'b0,layer_1_2[4279:4272]} - {1'b0, layer_0_2[4279:4272]};
      top_2[1] = {1'b0,layer_1_2[4287:4280]} - {1'b0, layer_0_2[4287:4280]};
      top_2[2] = {1'b0,layer_1_2[4295:4288]} - {1'b0, layer_0_2[4295:4288]};
      mid_0[0] = {1'b0,layer_2_0[4279:4272]} - {1'b0, layer_1_0[4279:4272]};
      mid_0[1] = {1'b0,layer_2_0[4287:4280]} - {1'b0, layer_1_0[4287:4280]};
      mid_0[2] = {1'b0,layer_2_0[4295:4288]} - {1'b0, layer_1_0[4295:4288]};
      mid_1[0] = {1'b0,layer_2_1[4279:4272]} - {1'b0, layer_1_1[4279:4272]};
      mid_1[1] = {1'b0,layer_2_1[4287:4280]} - {1'b0, layer_1_1[4287:4280]};
      mid_1[2] = {1'b0,layer_2_1[4295:4288]} - {1'b0, layer_1_1[4295:4288]};
      mid_2[0] = {1'b0,layer_2_2[4279:4272]} - {1'b0, layer_1_2[4279:4272]};
      mid_2[1] = {1'b0,layer_2_2[4287:4280]} - {1'b0, layer_1_2[4287:4280]};
      mid_2[2] = {1'b0,layer_2_2[4295:4288]} - {1'b0, layer_1_2[4295:4288]};
      btm_0[0] = {1'b0,layer_3_0[4279:4272]} - {1'b0, layer_2_0[4279:4272]};
      btm_0[1] = {1'b0,layer_3_0[4287:4280]} - {1'b0, layer_2_0[4287:4280]};
      btm_0[2] = {1'b0,layer_3_0[4295:4288]} - {1'b0, layer_2_0[4295:4288]};
      btm_1[0] = {1'b0,layer_3_1[4279:4272]} - {1'b0, layer_2_1[4279:4272]};
      btm_1[1] = {1'b0,layer_3_1[4287:4280]} - {1'b0, layer_2_1[4287:4280]};
      btm_1[2] = {1'b0,layer_3_1[4295:4288]} - {1'b0, layer_2_1[4295:4288]};
      btm_2[0] = {1'b0,layer_3_2[4279:4272]} - {1'b0, layer_2_2[4279:4272]};
      btm_2[1] = {1'b0,layer_3_2[4287:4280]} - {1'b0, layer_2_2[4287:4280]};
      btm_2[2] = {1'b0,layer_3_2[4295:4288]} - {1'b0, layer_2_2[4295:4288]};
    end
    'd536: begin
      top_0[0] = {1'b0,layer_1_0[4287:4280]} - {1'b0, layer_0_0[4287:4280]};
      top_0[1] = {1'b0,layer_1_0[4295:4288]} - {1'b0, layer_0_0[4295:4288]};
      top_0[2] = {1'b0,layer_1_0[4303:4296]} - {1'b0, layer_0_0[4303:4296]};
      top_1[0] = {1'b0,layer_1_1[4287:4280]} - {1'b0, layer_0_1[4287:4280]};
      top_1[1] = {1'b0,layer_1_1[4295:4288]} - {1'b0, layer_0_1[4295:4288]};
      top_1[2] = {1'b0,layer_1_1[4303:4296]} - {1'b0, layer_0_1[4303:4296]};
      top_2[0] = {1'b0,layer_1_2[4287:4280]} - {1'b0, layer_0_2[4287:4280]};
      top_2[1] = {1'b0,layer_1_2[4295:4288]} - {1'b0, layer_0_2[4295:4288]};
      top_2[2] = {1'b0,layer_1_2[4303:4296]} - {1'b0, layer_0_2[4303:4296]};
      mid_0[0] = {1'b0,layer_2_0[4287:4280]} - {1'b0, layer_1_0[4287:4280]};
      mid_0[1] = {1'b0,layer_2_0[4295:4288]} - {1'b0, layer_1_0[4295:4288]};
      mid_0[2] = {1'b0,layer_2_0[4303:4296]} - {1'b0, layer_1_0[4303:4296]};
      mid_1[0] = {1'b0,layer_2_1[4287:4280]} - {1'b0, layer_1_1[4287:4280]};
      mid_1[1] = {1'b0,layer_2_1[4295:4288]} - {1'b0, layer_1_1[4295:4288]};
      mid_1[2] = {1'b0,layer_2_1[4303:4296]} - {1'b0, layer_1_1[4303:4296]};
      mid_2[0] = {1'b0,layer_2_2[4287:4280]} - {1'b0, layer_1_2[4287:4280]};
      mid_2[1] = {1'b0,layer_2_2[4295:4288]} - {1'b0, layer_1_2[4295:4288]};
      mid_2[2] = {1'b0,layer_2_2[4303:4296]} - {1'b0, layer_1_2[4303:4296]};
      btm_0[0] = {1'b0,layer_3_0[4287:4280]} - {1'b0, layer_2_0[4287:4280]};
      btm_0[1] = {1'b0,layer_3_0[4295:4288]} - {1'b0, layer_2_0[4295:4288]};
      btm_0[2] = {1'b0,layer_3_0[4303:4296]} - {1'b0, layer_2_0[4303:4296]};
      btm_1[0] = {1'b0,layer_3_1[4287:4280]} - {1'b0, layer_2_1[4287:4280]};
      btm_1[1] = {1'b0,layer_3_1[4295:4288]} - {1'b0, layer_2_1[4295:4288]};
      btm_1[2] = {1'b0,layer_3_1[4303:4296]} - {1'b0, layer_2_1[4303:4296]};
      btm_2[0] = {1'b0,layer_3_2[4287:4280]} - {1'b0, layer_2_2[4287:4280]};
      btm_2[1] = {1'b0,layer_3_2[4295:4288]} - {1'b0, layer_2_2[4295:4288]};
      btm_2[2] = {1'b0,layer_3_2[4303:4296]} - {1'b0, layer_2_2[4303:4296]};
    end
    'd537: begin
      top_0[0] = {1'b0,layer_1_0[4295:4288]} - {1'b0, layer_0_0[4295:4288]};
      top_0[1] = {1'b0,layer_1_0[4303:4296]} - {1'b0, layer_0_0[4303:4296]};
      top_0[2] = {1'b0,layer_1_0[4311:4304]} - {1'b0, layer_0_0[4311:4304]};
      top_1[0] = {1'b0,layer_1_1[4295:4288]} - {1'b0, layer_0_1[4295:4288]};
      top_1[1] = {1'b0,layer_1_1[4303:4296]} - {1'b0, layer_0_1[4303:4296]};
      top_1[2] = {1'b0,layer_1_1[4311:4304]} - {1'b0, layer_0_1[4311:4304]};
      top_2[0] = {1'b0,layer_1_2[4295:4288]} - {1'b0, layer_0_2[4295:4288]};
      top_2[1] = {1'b0,layer_1_2[4303:4296]} - {1'b0, layer_0_2[4303:4296]};
      top_2[2] = {1'b0,layer_1_2[4311:4304]} - {1'b0, layer_0_2[4311:4304]};
      mid_0[0] = {1'b0,layer_2_0[4295:4288]} - {1'b0, layer_1_0[4295:4288]};
      mid_0[1] = {1'b0,layer_2_0[4303:4296]} - {1'b0, layer_1_0[4303:4296]};
      mid_0[2] = {1'b0,layer_2_0[4311:4304]} - {1'b0, layer_1_0[4311:4304]};
      mid_1[0] = {1'b0,layer_2_1[4295:4288]} - {1'b0, layer_1_1[4295:4288]};
      mid_1[1] = {1'b0,layer_2_1[4303:4296]} - {1'b0, layer_1_1[4303:4296]};
      mid_1[2] = {1'b0,layer_2_1[4311:4304]} - {1'b0, layer_1_1[4311:4304]};
      mid_2[0] = {1'b0,layer_2_2[4295:4288]} - {1'b0, layer_1_2[4295:4288]};
      mid_2[1] = {1'b0,layer_2_2[4303:4296]} - {1'b0, layer_1_2[4303:4296]};
      mid_2[2] = {1'b0,layer_2_2[4311:4304]} - {1'b0, layer_1_2[4311:4304]};
      btm_0[0] = {1'b0,layer_3_0[4295:4288]} - {1'b0, layer_2_0[4295:4288]};
      btm_0[1] = {1'b0,layer_3_0[4303:4296]} - {1'b0, layer_2_0[4303:4296]};
      btm_0[2] = {1'b0,layer_3_0[4311:4304]} - {1'b0, layer_2_0[4311:4304]};
      btm_1[0] = {1'b0,layer_3_1[4295:4288]} - {1'b0, layer_2_1[4295:4288]};
      btm_1[1] = {1'b0,layer_3_1[4303:4296]} - {1'b0, layer_2_1[4303:4296]};
      btm_1[2] = {1'b0,layer_3_1[4311:4304]} - {1'b0, layer_2_1[4311:4304]};
      btm_2[0] = {1'b0,layer_3_2[4295:4288]} - {1'b0, layer_2_2[4295:4288]};
      btm_2[1] = {1'b0,layer_3_2[4303:4296]} - {1'b0, layer_2_2[4303:4296]};
      btm_2[2] = {1'b0,layer_3_2[4311:4304]} - {1'b0, layer_2_2[4311:4304]};
    end
    'd538: begin
      top_0[0] = {1'b0,layer_1_0[4303:4296]} - {1'b0, layer_0_0[4303:4296]};
      top_0[1] = {1'b0,layer_1_0[4311:4304]} - {1'b0, layer_0_0[4311:4304]};
      top_0[2] = {1'b0,layer_1_0[4319:4312]} - {1'b0, layer_0_0[4319:4312]};
      top_1[0] = {1'b0,layer_1_1[4303:4296]} - {1'b0, layer_0_1[4303:4296]};
      top_1[1] = {1'b0,layer_1_1[4311:4304]} - {1'b0, layer_0_1[4311:4304]};
      top_1[2] = {1'b0,layer_1_1[4319:4312]} - {1'b0, layer_0_1[4319:4312]};
      top_2[0] = {1'b0,layer_1_2[4303:4296]} - {1'b0, layer_0_2[4303:4296]};
      top_2[1] = {1'b0,layer_1_2[4311:4304]} - {1'b0, layer_0_2[4311:4304]};
      top_2[2] = {1'b0,layer_1_2[4319:4312]} - {1'b0, layer_0_2[4319:4312]};
      mid_0[0] = {1'b0,layer_2_0[4303:4296]} - {1'b0, layer_1_0[4303:4296]};
      mid_0[1] = {1'b0,layer_2_0[4311:4304]} - {1'b0, layer_1_0[4311:4304]};
      mid_0[2] = {1'b0,layer_2_0[4319:4312]} - {1'b0, layer_1_0[4319:4312]};
      mid_1[0] = {1'b0,layer_2_1[4303:4296]} - {1'b0, layer_1_1[4303:4296]};
      mid_1[1] = {1'b0,layer_2_1[4311:4304]} - {1'b0, layer_1_1[4311:4304]};
      mid_1[2] = {1'b0,layer_2_1[4319:4312]} - {1'b0, layer_1_1[4319:4312]};
      mid_2[0] = {1'b0,layer_2_2[4303:4296]} - {1'b0, layer_1_2[4303:4296]};
      mid_2[1] = {1'b0,layer_2_2[4311:4304]} - {1'b0, layer_1_2[4311:4304]};
      mid_2[2] = {1'b0,layer_2_2[4319:4312]} - {1'b0, layer_1_2[4319:4312]};
      btm_0[0] = {1'b0,layer_3_0[4303:4296]} - {1'b0, layer_2_0[4303:4296]};
      btm_0[1] = {1'b0,layer_3_0[4311:4304]} - {1'b0, layer_2_0[4311:4304]};
      btm_0[2] = {1'b0,layer_3_0[4319:4312]} - {1'b0, layer_2_0[4319:4312]};
      btm_1[0] = {1'b0,layer_3_1[4303:4296]} - {1'b0, layer_2_1[4303:4296]};
      btm_1[1] = {1'b0,layer_3_1[4311:4304]} - {1'b0, layer_2_1[4311:4304]};
      btm_1[2] = {1'b0,layer_3_1[4319:4312]} - {1'b0, layer_2_1[4319:4312]};
      btm_2[0] = {1'b0,layer_3_2[4303:4296]} - {1'b0, layer_2_2[4303:4296]};
      btm_2[1] = {1'b0,layer_3_2[4311:4304]} - {1'b0, layer_2_2[4311:4304]};
      btm_2[2] = {1'b0,layer_3_2[4319:4312]} - {1'b0, layer_2_2[4319:4312]};
    end
    'd539: begin
      top_0[0] = {1'b0,layer_1_0[4311:4304]} - {1'b0, layer_0_0[4311:4304]};
      top_0[1] = {1'b0,layer_1_0[4319:4312]} - {1'b0, layer_0_0[4319:4312]};
      top_0[2] = {1'b0,layer_1_0[4327:4320]} - {1'b0, layer_0_0[4327:4320]};
      top_1[0] = {1'b0,layer_1_1[4311:4304]} - {1'b0, layer_0_1[4311:4304]};
      top_1[1] = {1'b0,layer_1_1[4319:4312]} - {1'b0, layer_0_1[4319:4312]};
      top_1[2] = {1'b0,layer_1_1[4327:4320]} - {1'b0, layer_0_1[4327:4320]};
      top_2[0] = {1'b0,layer_1_2[4311:4304]} - {1'b0, layer_0_2[4311:4304]};
      top_2[1] = {1'b0,layer_1_2[4319:4312]} - {1'b0, layer_0_2[4319:4312]};
      top_2[2] = {1'b0,layer_1_2[4327:4320]} - {1'b0, layer_0_2[4327:4320]};
      mid_0[0] = {1'b0,layer_2_0[4311:4304]} - {1'b0, layer_1_0[4311:4304]};
      mid_0[1] = {1'b0,layer_2_0[4319:4312]} - {1'b0, layer_1_0[4319:4312]};
      mid_0[2] = {1'b0,layer_2_0[4327:4320]} - {1'b0, layer_1_0[4327:4320]};
      mid_1[0] = {1'b0,layer_2_1[4311:4304]} - {1'b0, layer_1_1[4311:4304]};
      mid_1[1] = {1'b0,layer_2_1[4319:4312]} - {1'b0, layer_1_1[4319:4312]};
      mid_1[2] = {1'b0,layer_2_1[4327:4320]} - {1'b0, layer_1_1[4327:4320]};
      mid_2[0] = {1'b0,layer_2_2[4311:4304]} - {1'b0, layer_1_2[4311:4304]};
      mid_2[1] = {1'b0,layer_2_2[4319:4312]} - {1'b0, layer_1_2[4319:4312]};
      mid_2[2] = {1'b0,layer_2_2[4327:4320]} - {1'b0, layer_1_2[4327:4320]};
      btm_0[0] = {1'b0,layer_3_0[4311:4304]} - {1'b0, layer_2_0[4311:4304]};
      btm_0[1] = {1'b0,layer_3_0[4319:4312]} - {1'b0, layer_2_0[4319:4312]};
      btm_0[2] = {1'b0,layer_3_0[4327:4320]} - {1'b0, layer_2_0[4327:4320]};
      btm_1[0] = {1'b0,layer_3_1[4311:4304]} - {1'b0, layer_2_1[4311:4304]};
      btm_1[1] = {1'b0,layer_3_1[4319:4312]} - {1'b0, layer_2_1[4319:4312]};
      btm_1[2] = {1'b0,layer_3_1[4327:4320]} - {1'b0, layer_2_1[4327:4320]};
      btm_2[0] = {1'b0,layer_3_2[4311:4304]} - {1'b0, layer_2_2[4311:4304]};
      btm_2[1] = {1'b0,layer_3_2[4319:4312]} - {1'b0, layer_2_2[4319:4312]};
      btm_2[2] = {1'b0,layer_3_2[4327:4320]} - {1'b0, layer_2_2[4327:4320]};
    end
    'd540: begin
      top_0[0] = {1'b0,layer_1_0[4319:4312]} - {1'b0, layer_0_0[4319:4312]};
      top_0[1] = {1'b0,layer_1_0[4327:4320]} - {1'b0, layer_0_0[4327:4320]};
      top_0[2] = {1'b0,layer_1_0[4335:4328]} - {1'b0, layer_0_0[4335:4328]};
      top_1[0] = {1'b0,layer_1_1[4319:4312]} - {1'b0, layer_0_1[4319:4312]};
      top_1[1] = {1'b0,layer_1_1[4327:4320]} - {1'b0, layer_0_1[4327:4320]};
      top_1[2] = {1'b0,layer_1_1[4335:4328]} - {1'b0, layer_0_1[4335:4328]};
      top_2[0] = {1'b0,layer_1_2[4319:4312]} - {1'b0, layer_0_2[4319:4312]};
      top_2[1] = {1'b0,layer_1_2[4327:4320]} - {1'b0, layer_0_2[4327:4320]};
      top_2[2] = {1'b0,layer_1_2[4335:4328]} - {1'b0, layer_0_2[4335:4328]};
      mid_0[0] = {1'b0,layer_2_0[4319:4312]} - {1'b0, layer_1_0[4319:4312]};
      mid_0[1] = {1'b0,layer_2_0[4327:4320]} - {1'b0, layer_1_0[4327:4320]};
      mid_0[2] = {1'b0,layer_2_0[4335:4328]} - {1'b0, layer_1_0[4335:4328]};
      mid_1[0] = {1'b0,layer_2_1[4319:4312]} - {1'b0, layer_1_1[4319:4312]};
      mid_1[1] = {1'b0,layer_2_1[4327:4320]} - {1'b0, layer_1_1[4327:4320]};
      mid_1[2] = {1'b0,layer_2_1[4335:4328]} - {1'b0, layer_1_1[4335:4328]};
      mid_2[0] = {1'b0,layer_2_2[4319:4312]} - {1'b0, layer_1_2[4319:4312]};
      mid_2[1] = {1'b0,layer_2_2[4327:4320]} - {1'b0, layer_1_2[4327:4320]};
      mid_2[2] = {1'b0,layer_2_2[4335:4328]} - {1'b0, layer_1_2[4335:4328]};
      btm_0[0] = {1'b0,layer_3_0[4319:4312]} - {1'b0, layer_2_0[4319:4312]};
      btm_0[1] = {1'b0,layer_3_0[4327:4320]} - {1'b0, layer_2_0[4327:4320]};
      btm_0[2] = {1'b0,layer_3_0[4335:4328]} - {1'b0, layer_2_0[4335:4328]};
      btm_1[0] = {1'b0,layer_3_1[4319:4312]} - {1'b0, layer_2_1[4319:4312]};
      btm_1[1] = {1'b0,layer_3_1[4327:4320]} - {1'b0, layer_2_1[4327:4320]};
      btm_1[2] = {1'b0,layer_3_1[4335:4328]} - {1'b0, layer_2_1[4335:4328]};
      btm_2[0] = {1'b0,layer_3_2[4319:4312]} - {1'b0, layer_2_2[4319:4312]};
      btm_2[1] = {1'b0,layer_3_2[4327:4320]} - {1'b0, layer_2_2[4327:4320]};
      btm_2[2] = {1'b0,layer_3_2[4335:4328]} - {1'b0, layer_2_2[4335:4328]};
    end
    'd541: begin
      top_0[0] = {1'b0,layer_1_0[4327:4320]} - {1'b0, layer_0_0[4327:4320]};
      top_0[1] = {1'b0,layer_1_0[4335:4328]} - {1'b0, layer_0_0[4335:4328]};
      top_0[2] = {1'b0,layer_1_0[4343:4336]} - {1'b0, layer_0_0[4343:4336]};
      top_1[0] = {1'b0,layer_1_1[4327:4320]} - {1'b0, layer_0_1[4327:4320]};
      top_1[1] = {1'b0,layer_1_1[4335:4328]} - {1'b0, layer_0_1[4335:4328]};
      top_1[2] = {1'b0,layer_1_1[4343:4336]} - {1'b0, layer_0_1[4343:4336]};
      top_2[0] = {1'b0,layer_1_2[4327:4320]} - {1'b0, layer_0_2[4327:4320]};
      top_2[1] = {1'b0,layer_1_2[4335:4328]} - {1'b0, layer_0_2[4335:4328]};
      top_2[2] = {1'b0,layer_1_2[4343:4336]} - {1'b0, layer_0_2[4343:4336]};
      mid_0[0] = {1'b0,layer_2_0[4327:4320]} - {1'b0, layer_1_0[4327:4320]};
      mid_0[1] = {1'b0,layer_2_0[4335:4328]} - {1'b0, layer_1_0[4335:4328]};
      mid_0[2] = {1'b0,layer_2_0[4343:4336]} - {1'b0, layer_1_0[4343:4336]};
      mid_1[0] = {1'b0,layer_2_1[4327:4320]} - {1'b0, layer_1_1[4327:4320]};
      mid_1[1] = {1'b0,layer_2_1[4335:4328]} - {1'b0, layer_1_1[4335:4328]};
      mid_1[2] = {1'b0,layer_2_1[4343:4336]} - {1'b0, layer_1_1[4343:4336]};
      mid_2[0] = {1'b0,layer_2_2[4327:4320]} - {1'b0, layer_1_2[4327:4320]};
      mid_2[1] = {1'b0,layer_2_2[4335:4328]} - {1'b0, layer_1_2[4335:4328]};
      mid_2[2] = {1'b0,layer_2_2[4343:4336]} - {1'b0, layer_1_2[4343:4336]};
      btm_0[0] = {1'b0,layer_3_0[4327:4320]} - {1'b0, layer_2_0[4327:4320]};
      btm_0[1] = {1'b0,layer_3_0[4335:4328]} - {1'b0, layer_2_0[4335:4328]};
      btm_0[2] = {1'b0,layer_3_0[4343:4336]} - {1'b0, layer_2_0[4343:4336]};
      btm_1[0] = {1'b0,layer_3_1[4327:4320]} - {1'b0, layer_2_1[4327:4320]};
      btm_1[1] = {1'b0,layer_3_1[4335:4328]} - {1'b0, layer_2_1[4335:4328]};
      btm_1[2] = {1'b0,layer_3_1[4343:4336]} - {1'b0, layer_2_1[4343:4336]};
      btm_2[0] = {1'b0,layer_3_2[4327:4320]} - {1'b0, layer_2_2[4327:4320]};
      btm_2[1] = {1'b0,layer_3_2[4335:4328]} - {1'b0, layer_2_2[4335:4328]};
      btm_2[2] = {1'b0,layer_3_2[4343:4336]} - {1'b0, layer_2_2[4343:4336]};
    end
    'd542: begin
      top_0[0] = {1'b0,layer_1_0[4335:4328]} - {1'b0, layer_0_0[4335:4328]};
      top_0[1] = {1'b0,layer_1_0[4343:4336]} - {1'b0, layer_0_0[4343:4336]};
      top_0[2] = {1'b0,layer_1_0[4351:4344]} - {1'b0, layer_0_0[4351:4344]};
      top_1[0] = {1'b0,layer_1_1[4335:4328]} - {1'b0, layer_0_1[4335:4328]};
      top_1[1] = {1'b0,layer_1_1[4343:4336]} - {1'b0, layer_0_1[4343:4336]};
      top_1[2] = {1'b0,layer_1_1[4351:4344]} - {1'b0, layer_0_1[4351:4344]};
      top_2[0] = {1'b0,layer_1_2[4335:4328]} - {1'b0, layer_0_2[4335:4328]};
      top_2[1] = {1'b0,layer_1_2[4343:4336]} - {1'b0, layer_0_2[4343:4336]};
      top_2[2] = {1'b0,layer_1_2[4351:4344]} - {1'b0, layer_0_2[4351:4344]};
      mid_0[0] = {1'b0,layer_2_0[4335:4328]} - {1'b0, layer_1_0[4335:4328]};
      mid_0[1] = {1'b0,layer_2_0[4343:4336]} - {1'b0, layer_1_0[4343:4336]};
      mid_0[2] = {1'b0,layer_2_0[4351:4344]} - {1'b0, layer_1_0[4351:4344]};
      mid_1[0] = {1'b0,layer_2_1[4335:4328]} - {1'b0, layer_1_1[4335:4328]};
      mid_1[1] = {1'b0,layer_2_1[4343:4336]} - {1'b0, layer_1_1[4343:4336]};
      mid_1[2] = {1'b0,layer_2_1[4351:4344]} - {1'b0, layer_1_1[4351:4344]};
      mid_2[0] = {1'b0,layer_2_2[4335:4328]} - {1'b0, layer_1_2[4335:4328]};
      mid_2[1] = {1'b0,layer_2_2[4343:4336]} - {1'b0, layer_1_2[4343:4336]};
      mid_2[2] = {1'b0,layer_2_2[4351:4344]} - {1'b0, layer_1_2[4351:4344]};
      btm_0[0] = {1'b0,layer_3_0[4335:4328]} - {1'b0, layer_2_0[4335:4328]};
      btm_0[1] = {1'b0,layer_3_0[4343:4336]} - {1'b0, layer_2_0[4343:4336]};
      btm_0[2] = {1'b0,layer_3_0[4351:4344]} - {1'b0, layer_2_0[4351:4344]};
      btm_1[0] = {1'b0,layer_3_1[4335:4328]} - {1'b0, layer_2_1[4335:4328]};
      btm_1[1] = {1'b0,layer_3_1[4343:4336]} - {1'b0, layer_2_1[4343:4336]};
      btm_1[2] = {1'b0,layer_3_1[4351:4344]} - {1'b0, layer_2_1[4351:4344]};
      btm_2[0] = {1'b0,layer_3_2[4335:4328]} - {1'b0, layer_2_2[4335:4328]};
      btm_2[1] = {1'b0,layer_3_2[4343:4336]} - {1'b0, layer_2_2[4343:4336]};
      btm_2[2] = {1'b0,layer_3_2[4351:4344]} - {1'b0, layer_2_2[4351:4344]};
    end
    'd543: begin
      top_0[0] = {1'b0,layer_1_0[4343:4336]} - {1'b0, layer_0_0[4343:4336]};
      top_0[1] = {1'b0,layer_1_0[4351:4344]} - {1'b0, layer_0_0[4351:4344]};
      top_0[2] = {1'b0,layer_1_0[4359:4352]} - {1'b0, layer_0_0[4359:4352]};
      top_1[0] = {1'b0,layer_1_1[4343:4336]} - {1'b0, layer_0_1[4343:4336]};
      top_1[1] = {1'b0,layer_1_1[4351:4344]} - {1'b0, layer_0_1[4351:4344]};
      top_1[2] = {1'b0,layer_1_1[4359:4352]} - {1'b0, layer_0_1[4359:4352]};
      top_2[0] = {1'b0,layer_1_2[4343:4336]} - {1'b0, layer_0_2[4343:4336]};
      top_2[1] = {1'b0,layer_1_2[4351:4344]} - {1'b0, layer_0_2[4351:4344]};
      top_2[2] = {1'b0,layer_1_2[4359:4352]} - {1'b0, layer_0_2[4359:4352]};
      mid_0[0] = {1'b0,layer_2_0[4343:4336]} - {1'b0, layer_1_0[4343:4336]};
      mid_0[1] = {1'b0,layer_2_0[4351:4344]} - {1'b0, layer_1_0[4351:4344]};
      mid_0[2] = {1'b0,layer_2_0[4359:4352]} - {1'b0, layer_1_0[4359:4352]};
      mid_1[0] = {1'b0,layer_2_1[4343:4336]} - {1'b0, layer_1_1[4343:4336]};
      mid_1[1] = {1'b0,layer_2_1[4351:4344]} - {1'b0, layer_1_1[4351:4344]};
      mid_1[2] = {1'b0,layer_2_1[4359:4352]} - {1'b0, layer_1_1[4359:4352]};
      mid_2[0] = {1'b0,layer_2_2[4343:4336]} - {1'b0, layer_1_2[4343:4336]};
      mid_2[1] = {1'b0,layer_2_2[4351:4344]} - {1'b0, layer_1_2[4351:4344]};
      mid_2[2] = {1'b0,layer_2_2[4359:4352]} - {1'b0, layer_1_2[4359:4352]};
      btm_0[0] = {1'b0,layer_3_0[4343:4336]} - {1'b0, layer_2_0[4343:4336]};
      btm_0[1] = {1'b0,layer_3_0[4351:4344]} - {1'b0, layer_2_0[4351:4344]};
      btm_0[2] = {1'b0,layer_3_0[4359:4352]} - {1'b0, layer_2_0[4359:4352]};
      btm_1[0] = {1'b0,layer_3_1[4343:4336]} - {1'b0, layer_2_1[4343:4336]};
      btm_1[1] = {1'b0,layer_3_1[4351:4344]} - {1'b0, layer_2_1[4351:4344]};
      btm_1[2] = {1'b0,layer_3_1[4359:4352]} - {1'b0, layer_2_1[4359:4352]};
      btm_2[0] = {1'b0,layer_3_2[4343:4336]} - {1'b0, layer_2_2[4343:4336]};
      btm_2[1] = {1'b0,layer_3_2[4351:4344]} - {1'b0, layer_2_2[4351:4344]};
      btm_2[2] = {1'b0,layer_3_2[4359:4352]} - {1'b0, layer_2_2[4359:4352]};
    end
    'd544: begin
      top_0[0] = {1'b0,layer_1_0[4351:4344]} - {1'b0, layer_0_0[4351:4344]};
      top_0[1] = {1'b0,layer_1_0[4359:4352]} - {1'b0, layer_0_0[4359:4352]};
      top_0[2] = {1'b0,layer_1_0[4367:4360]} - {1'b0, layer_0_0[4367:4360]};
      top_1[0] = {1'b0,layer_1_1[4351:4344]} - {1'b0, layer_0_1[4351:4344]};
      top_1[1] = {1'b0,layer_1_1[4359:4352]} - {1'b0, layer_0_1[4359:4352]};
      top_1[2] = {1'b0,layer_1_1[4367:4360]} - {1'b0, layer_0_1[4367:4360]};
      top_2[0] = {1'b0,layer_1_2[4351:4344]} - {1'b0, layer_0_2[4351:4344]};
      top_2[1] = {1'b0,layer_1_2[4359:4352]} - {1'b0, layer_0_2[4359:4352]};
      top_2[2] = {1'b0,layer_1_2[4367:4360]} - {1'b0, layer_0_2[4367:4360]};
      mid_0[0] = {1'b0,layer_2_0[4351:4344]} - {1'b0, layer_1_0[4351:4344]};
      mid_0[1] = {1'b0,layer_2_0[4359:4352]} - {1'b0, layer_1_0[4359:4352]};
      mid_0[2] = {1'b0,layer_2_0[4367:4360]} - {1'b0, layer_1_0[4367:4360]};
      mid_1[0] = {1'b0,layer_2_1[4351:4344]} - {1'b0, layer_1_1[4351:4344]};
      mid_1[1] = {1'b0,layer_2_1[4359:4352]} - {1'b0, layer_1_1[4359:4352]};
      mid_1[2] = {1'b0,layer_2_1[4367:4360]} - {1'b0, layer_1_1[4367:4360]};
      mid_2[0] = {1'b0,layer_2_2[4351:4344]} - {1'b0, layer_1_2[4351:4344]};
      mid_2[1] = {1'b0,layer_2_2[4359:4352]} - {1'b0, layer_1_2[4359:4352]};
      mid_2[2] = {1'b0,layer_2_2[4367:4360]} - {1'b0, layer_1_2[4367:4360]};
      btm_0[0] = {1'b0,layer_3_0[4351:4344]} - {1'b0, layer_2_0[4351:4344]};
      btm_0[1] = {1'b0,layer_3_0[4359:4352]} - {1'b0, layer_2_0[4359:4352]};
      btm_0[2] = {1'b0,layer_3_0[4367:4360]} - {1'b0, layer_2_0[4367:4360]};
      btm_1[0] = {1'b0,layer_3_1[4351:4344]} - {1'b0, layer_2_1[4351:4344]};
      btm_1[1] = {1'b0,layer_3_1[4359:4352]} - {1'b0, layer_2_1[4359:4352]};
      btm_1[2] = {1'b0,layer_3_1[4367:4360]} - {1'b0, layer_2_1[4367:4360]};
      btm_2[0] = {1'b0,layer_3_2[4351:4344]} - {1'b0, layer_2_2[4351:4344]};
      btm_2[1] = {1'b0,layer_3_2[4359:4352]} - {1'b0, layer_2_2[4359:4352]};
      btm_2[2] = {1'b0,layer_3_2[4367:4360]} - {1'b0, layer_2_2[4367:4360]};
    end
    'd545: begin
      top_0[0] = {1'b0,layer_1_0[4359:4352]} - {1'b0, layer_0_0[4359:4352]};
      top_0[1] = {1'b0,layer_1_0[4367:4360]} - {1'b0, layer_0_0[4367:4360]};
      top_0[2] = {1'b0,layer_1_0[4375:4368]} - {1'b0, layer_0_0[4375:4368]};
      top_1[0] = {1'b0,layer_1_1[4359:4352]} - {1'b0, layer_0_1[4359:4352]};
      top_1[1] = {1'b0,layer_1_1[4367:4360]} - {1'b0, layer_0_1[4367:4360]};
      top_1[2] = {1'b0,layer_1_1[4375:4368]} - {1'b0, layer_0_1[4375:4368]};
      top_2[0] = {1'b0,layer_1_2[4359:4352]} - {1'b0, layer_0_2[4359:4352]};
      top_2[1] = {1'b0,layer_1_2[4367:4360]} - {1'b0, layer_0_2[4367:4360]};
      top_2[2] = {1'b0,layer_1_2[4375:4368]} - {1'b0, layer_0_2[4375:4368]};
      mid_0[0] = {1'b0,layer_2_0[4359:4352]} - {1'b0, layer_1_0[4359:4352]};
      mid_0[1] = {1'b0,layer_2_0[4367:4360]} - {1'b0, layer_1_0[4367:4360]};
      mid_0[2] = {1'b0,layer_2_0[4375:4368]} - {1'b0, layer_1_0[4375:4368]};
      mid_1[0] = {1'b0,layer_2_1[4359:4352]} - {1'b0, layer_1_1[4359:4352]};
      mid_1[1] = {1'b0,layer_2_1[4367:4360]} - {1'b0, layer_1_1[4367:4360]};
      mid_1[2] = {1'b0,layer_2_1[4375:4368]} - {1'b0, layer_1_1[4375:4368]};
      mid_2[0] = {1'b0,layer_2_2[4359:4352]} - {1'b0, layer_1_2[4359:4352]};
      mid_2[1] = {1'b0,layer_2_2[4367:4360]} - {1'b0, layer_1_2[4367:4360]};
      mid_2[2] = {1'b0,layer_2_2[4375:4368]} - {1'b0, layer_1_2[4375:4368]};
      btm_0[0] = {1'b0,layer_3_0[4359:4352]} - {1'b0, layer_2_0[4359:4352]};
      btm_0[1] = {1'b0,layer_3_0[4367:4360]} - {1'b0, layer_2_0[4367:4360]};
      btm_0[2] = {1'b0,layer_3_0[4375:4368]} - {1'b0, layer_2_0[4375:4368]};
      btm_1[0] = {1'b0,layer_3_1[4359:4352]} - {1'b0, layer_2_1[4359:4352]};
      btm_1[1] = {1'b0,layer_3_1[4367:4360]} - {1'b0, layer_2_1[4367:4360]};
      btm_1[2] = {1'b0,layer_3_1[4375:4368]} - {1'b0, layer_2_1[4375:4368]};
      btm_2[0] = {1'b0,layer_3_2[4359:4352]} - {1'b0, layer_2_2[4359:4352]};
      btm_2[1] = {1'b0,layer_3_2[4367:4360]} - {1'b0, layer_2_2[4367:4360]};
      btm_2[2] = {1'b0,layer_3_2[4375:4368]} - {1'b0, layer_2_2[4375:4368]};
    end
    'd546: begin
      top_0[0] = {1'b0,layer_1_0[4367:4360]} - {1'b0, layer_0_0[4367:4360]};
      top_0[1] = {1'b0,layer_1_0[4375:4368]} - {1'b0, layer_0_0[4375:4368]};
      top_0[2] = {1'b0,layer_1_0[4383:4376]} - {1'b0, layer_0_0[4383:4376]};
      top_1[0] = {1'b0,layer_1_1[4367:4360]} - {1'b0, layer_0_1[4367:4360]};
      top_1[1] = {1'b0,layer_1_1[4375:4368]} - {1'b0, layer_0_1[4375:4368]};
      top_1[2] = {1'b0,layer_1_1[4383:4376]} - {1'b0, layer_0_1[4383:4376]};
      top_2[0] = {1'b0,layer_1_2[4367:4360]} - {1'b0, layer_0_2[4367:4360]};
      top_2[1] = {1'b0,layer_1_2[4375:4368]} - {1'b0, layer_0_2[4375:4368]};
      top_2[2] = {1'b0,layer_1_2[4383:4376]} - {1'b0, layer_0_2[4383:4376]};
      mid_0[0] = {1'b0,layer_2_0[4367:4360]} - {1'b0, layer_1_0[4367:4360]};
      mid_0[1] = {1'b0,layer_2_0[4375:4368]} - {1'b0, layer_1_0[4375:4368]};
      mid_0[2] = {1'b0,layer_2_0[4383:4376]} - {1'b0, layer_1_0[4383:4376]};
      mid_1[0] = {1'b0,layer_2_1[4367:4360]} - {1'b0, layer_1_1[4367:4360]};
      mid_1[1] = {1'b0,layer_2_1[4375:4368]} - {1'b0, layer_1_1[4375:4368]};
      mid_1[2] = {1'b0,layer_2_1[4383:4376]} - {1'b0, layer_1_1[4383:4376]};
      mid_2[0] = {1'b0,layer_2_2[4367:4360]} - {1'b0, layer_1_2[4367:4360]};
      mid_2[1] = {1'b0,layer_2_2[4375:4368]} - {1'b0, layer_1_2[4375:4368]};
      mid_2[2] = {1'b0,layer_2_2[4383:4376]} - {1'b0, layer_1_2[4383:4376]};
      btm_0[0] = {1'b0,layer_3_0[4367:4360]} - {1'b0, layer_2_0[4367:4360]};
      btm_0[1] = {1'b0,layer_3_0[4375:4368]} - {1'b0, layer_2_0[4375:4368]};
      btm_0[2] = {1'b0,layer_3_0[4383:4376]} - {1'b0, layer_2_0[4383:4376]};
      btm_1[0] = {1'b0,layer_3_1[4367:4360]} - {1'b0, layer_2_1[4367:4360]};
      btm_1[1] = {1'b0,layer_3_1[4375:4368]} - {1'b0, layer_2_1[4375:4368]};
      btm_1[2] = {1'b0,layer_3_1[4383:4376]} - {1'b0, layer_2_1[4383:4376]};
      btm_2[0] = {1'b0,layer_3_2[4367:4360]} - {1'b0, layer_2_2[4367:4360]};
      btm_2[1] = {1'b0,layer_3_2[4375:4368]} - {1'b0, layer_2_2[4375:4368]};
      btm_2[2] = {1'b0,layer_3_2[4383:4376]} - {1'b0, layer_2_2[4383:4376]};
    end
    'd547: begin
      top_0[0] = {1'b0,layer_1_0[4375:4368]} - {1'b0, layer_0_0[4375:4368]};
      top_0[1] = {1'b0,layer_1_0[4383:4376]} - {1'b0, layer_0_0[4383:4376]};
      top_0[2] = {1'b0,layer_1_0[4391:4384]} - {1'b0, layer_0_0[4391:4384]};
      top_1[0] = {1'b0,layer_1_1[4375:4368]} - {1'b0, layer_0_1[4375:4368]};
      top_1[1] = {1'b0,layer_1_1[4383:4376]} - {1'b0, layer_0_1[4383:4376]};
      top_1[2] = {1'b0,layer_1_1[4391:4384]} - {1'b0, layer_0_1[4391:4384]};
      top_2[0] = {1'b0,layer_1_2[4375:4368]} - {1'b0, layer_0_2[4375:4368]};
      top_2[1] = {1'b0,layer_1_2[4383:4376]} - {1'b0, layer_0_2[4383:4376]};
      top_2[2] = {1'b0,layer_1_2[4391:4384]} - {1'b0, layer_0_2[4391:4384]};
      mid_0[0] = {1'b0,layer_2_0[4375:4368]} - {1'b0, layer_1_0[4375:4368]};
      mid_0[1] = {1'b0,layer_2_0[4383:4376]} - {1'b0, layer_1_0[4383:4376]};
      mid_0[2] = {1'b0,layer_2_0[4391:4384]} - {1'b0, layer_1_0[4391:4384]};
      mid_1[0] = {1'b0,layer_2_1[4375:4368]} - {1'b0, layer_1_1[4375:4368]};
      mid_1[1] = {1'b0,layer_2_1[4383:4376]} - {1'b0, layer_1_1[4383:4376]};
      mid_1[2] = {1'b0,layer_2_1[4391:4384]} - {1'b0, layer_1_1[4391:4384]};
      mid_2[0] = {1'b0,layer_2_2[4375:4368]} - {1'b0, layer_1_2[4375:4368]};
      mid_2[1] = {1'b0,layer_2_2[4383:4376]} - {1'b0, layer_1_2[4383:4376]};
      mid_2[2] = {1'b0,layer_2_2[4391:4384]} - {1'b0, layer_1_2[4391:4384]};
      btm_0[0] = {1'b0,layer_3_0[4375:4368]} - {1'b0, layer_2_0[4375:4368]};
      btm_0[1] = {1'b0,layer_3_0[4383:4376]} - {1'b0, layer_2_0[4383:4376]};
      btm_0[2] = {1'b0,layer_3_0[4391:4384]} - {1'b0, layer_2_0[4391:4384]};
      btm_1[0] = {1'b0,layer_3_1[4375:4368]} - {1'b0, layer_2_1[4375:4368]};
      btm_1[1] = {1'b0,layer_3_1[4383:4376]} - {1'b0, layer_2_1[4383:4376]};
      btm_1[2] = {1'b0,layer_3_1[4391:4384]} - {1'b0, layer_2_1[4391:4384]};
      btm_2[0] = {1'b0,layer_3_2[4375:4368]} - {1'b0, layer_2_2[4375:4368]};
      btm_2[1] = {1'b0,layer_3_2[4383:4376]} - {1'b0, layer_2_2[4383:4376]};
      btm_2[2] = {1'b0,layer_3_2[4391:4384]} - {1'b0, layer_2_2[4391:4384]};
    end
    'd548: begin
      top_0[0] = {1'b0,layer_1_0[4383:4376]} - {1'b0, layer_0_0[4383:4376]};
      top_0[1] = {1'b0,layer_1_0[4391:4384]} - {1'b0, layer_0_0[4391:4384]};
      top_0[2] = {1'b0,layer_1_0[4399:4392]} - {1'b0, layer_0_0[4399:4392]};
      top_1[0] = {1'b0,layer_1_1[4383:4376]} - {1'b0, layer_0_1[4383:4376]};
      top_1[1] = {1'b0,layer_1_1[4391:4384]} - {1'b0, layer_0_1[4391:4384]};
      top_1[2] = {1'b0,layer_1_1[4399:4392]} - {1'b0, layer_0_1[4399:4392]};
      top_2[0] = {1'b0,layer_1_2[4383:4376]} - {1'b0, layer_0_2[4383:4376]};
      top_2[1] = {1'b0,layer_1_2[4391:4384]} - {1'b0, layer_0_2[4391:4384]};
      top_2[2] = {1'b0,layer_1_2[4399:4392]} - {1'b0, layer_0_2[4399:4392]};
      mid_0[0] = {1'b0,layer_2_0[4383:4376]} - {1'b0, layer_1_0[4383:4376]};
      mid_0[1] = {1'b0,layer_2_0[4391:4384]} - {1'b0, layer_1_0[4391:4384]};
      mid_0[2] = {1'b0,layer_2_0[4399:4392]} - {1'b0, layer_1_0[4399:4392]};
      mid_1[0] = {1'b0,layer_2_1[4383:4376]} - {1'b0, layer_1_1[4383:4376]};
      mid_1[1] = {1'b0,layer_2_1[4391:4384]} - {1'b0, layer_1_1[4391:4384]};
      mid_1[2] = {1'b0,layer_2_1[4399:4392]} - {1'b0, layer_1_1[4399:4392]};
      mid_2[0] = {1'b0,layer_2_2[4383:4376]} - {1'b0, layer_1_2[4383:4376]};
      mid_2[1] = {1'b0,layer_2_2[4391:4384]} - {1'b0, layer_1_2[4391:4384]};
      mid_2[2] = {1'b0,layer_2_2[4399:4392]} - {1'b0, layer_1_2[4399:4392]};
      btm_0[0] = {1'b0,layer_3_0[4383:4376]} - {1'b0, layer_2_0[4383:4376]};
      btm_0[1] = {1'b0,layer_3_0[4391:4384]} - {1'b0, layer_2_0[4391:4384]};
      btm_0[2] = {1'b0,layer_3_0[4399:4392]} - {1'b0, layer_2_0[4399:4392]};
      btm_1[0] = {1'b0,layer_3_1[4383:4376]} - {1'b0, layer_2_1[4383:4376]};
      btm_1[1] = {1'b0,layer_3_1[4391:4384]} - {1'b0, layer_2_1[4391:4384]};
      btm_1[2] = {1'b0,layer_3_1[4399:4392]} - {1'b0, layer_2_1[4399:4392]};
      btm_2[0] = {1'b0,layer_3_2[4383:4376]} - {1'b0, layer_2_2[4383:4376]};
      btm_2[1] = {1'b0,layer_3_2[4391:4384]} - {1'b0, layer_2_2[4391:4384]};
      btm_2[2] = {1'b0,layer_3_2[4399:4392]} - {1'b0, layer_2_2[4399:4392]};
    end
    'd549: begin
      top_0[0] = {1'b0,layer_1_0[4391:4384]} - {1'b0, layer_0_0[4391:4384]};
      top_0[1] = {1'b0,layer_1_0[4399:4392]} - {1'b0, layer_0_0[4399:4392]};
      top_0[2] = {1'b0,layer_1_0[4407:4400]} - {1'b0, layer_0_0[4407:4400]};
      top_1[0] = {1'b0,layer_1_1[4391:4384]} - {1'b0, layer_0_1[4391:4384]};
      top_1[1] = {1'b0,layer_1_1[4399:4392]} - {1'b0, layer_0_1[4399:4392]};
      top_1[2] = {1'b0,layer_1_1[4407:4400]} - {1'b0, layer_0_1[4407:4400]};
      top_2[0] = {1'b0,layer_1_2[4391:4384]} - {1'b0, layer_0_2[4391:4384]};
      top_2[1] = {1'b0,layer_1_2[4399:4392]} - {1'b0, layer_0_2[4399:4392]};
      top_2[2] = {1'b0,layer_1_2[4407:4400]} - {1'b0, layer_0_2[4407:4400]};
      mid_0[0] = {1'b0,layer_2_0[4391:4384]} - {1'b0, layer_1_0[4391:4384]};
      mid_0[1] = {1'b0,layer_2_0[4399:4392]} - {1'b0, layer_1_0[4399:4392]};
      mid_0[2] = {1'b0,layer_2_0[4407:4400]} - {1'b0, layer_1_0[4407:4400]};
      mid_1[0] = {1'b0,layer_2_1[4391:4384]} - {1'b0, layer_1_1[4391:4384]};
      mid_1[1] = {1'b0,layer_2_1[4399:4392]} - {1'b0, layer_1_1[4399:4392]};
      mid_1[2] = {1'b0,layer_2_1[4407:4400]} - {1'b0, layer_1_1[4407:4400]};
      mid_2[0] = {1'b0,layer_2_2[4391:4384]} - {1'b0, layer_1_2[4391:4384]};
      mid_2[1] = {1'b0,layer_2_2[4399:4392]} - {1'b0, layer_1_2[4399:4392]};
      mid_2[2] = {1'b0,layer_2_2[4407:4400]} - {1'b0, layer_1_2[4407:4400]};
      btm_0[0] = {1'b0,layer_3_0[4391:4384]} - {1'b0, layer_2_0[4391:4384]};
      btm_0[1] = {1'b0,layer_3_0[4399:4392]} - {1'b0, layer_2_0[4399:4392]};
      btm_0[2] = {1'b0,layer_3_0[4407:4400]} - {1'b0, layer_2_0[4407:4400]};
      btm_1[0] = {1'b0,layer_3_1[4391:4384]} - {1'b0, layer_2_1[4391:4384]};
      btm_1[1] = {1'b0,layer_3_1[4399:4392]} - {1'b0, layer_2_1[4399:4392]};
      btm_1[2] = {1'b0,layer_3_1[4407:4400]} - {1'b0, layer_2_1[4407:4400]};
      btm_2[0] = {1'b0,layer_3_2[4391:4384]} - {1'b0, layer_2_2[4391:4384]};
      btm_2[1] = {1'b0,layer_3_2[4399:4392]} - {1'b0, layer_2_2[4399:4392]};
      btm_2[2] = {1'b0,layer_3_2[4407:4400]} - {1'b0, layer_2_2[4407:4400]};
    end
    'd550: begin
      top_0[0] = {1'b0,layer_1_0[4399:4392]} - {1'b0, layer_0_0[4399:4392]};
      top_0[1] = {1'b0,layer_1_0[4407:4400]} - {1'b0, layer_0_0[4407:4400]};
      top_0[2] = {1'b0,layer_1_0[4415:4408]} - {1'b0, layer_0_0[4415:4408]};
      top_1[0] = {1'b0,layer_1_1[4399:4392]} - {1'b0, layer_0_1[4399:4392]};
      top_1[1] = {1'b0,layer_1_1[4407:4400]} - {1'b0, layer_0_1[4407:4400]};
      top_1[2] = {1'b0,layer_1_1[4415:4408]} - {1'b0, layer_0_1[4415:4408]};
      top_2[0] = {1'b0,layer_1_2[4399:4392]} - {1'b0, layer_0_2[4399:4392]};
      top_2[1] = {1'b0,layer_1_2[4407:4400]} - {1'b0, layer_0_2[4407:4400]};
      top_2[2] = {1'b0,layer_1_2[4415:4408]} - {1'b0, layer_0_2[4415:4408]};
      mid_0[0] = {1'b0,layer_2_0[4399:4392]} - {1'b0, layer_1_0[4399:4392]};
      mid_0[1] = {1'b0,layer_2_0[4407:4400]} - {1'b0, layer_1_0[4407:4400]};
      mid_0[2] = {1'b0,layer_2_0[4415:4408]} - {1'b0, layer_1_0[4415:4408]};
      mid_1[0] = {1'b0,layer_2_1[4399:4392]} - {1'b0, layer_1_1[4399:4392]};
      mid_1[1] = {1'b0,layer_2_1[4407:4400]} - {1'b0, layer_1_1[4407:4400]};
      mid_1[2] = {1'b0,layer_2_1[4415:4408]} - {1'b0, layer_1_1[4415:4408]};
      mid_2[0] = {1'b0,layer_2_2[4399:4392]} - {1'b0, layer_1_2[4399:4392]};
      mid_2[1] = {1'b0,layer_2_2[4407:4400]} - {1'b0, layer_1_2[4407:4400]};
      mid_2[2] = {1'b0,layer_2_2[4415:4408]} - {1'b0, layer_1_2[4415:4408]};
      btm_0[0] = {1'b0,layer_3_0[4399:4392]} - {1'b0, layer_2_0[4399:4392]};
      btm_0[1] = {1'b0,layer_3_0[4407:4400]} - {1'b0, layer_2_0[4407:4400]};
      btm_0[2] = {1'b0,layer_3_0[4415:4408]} - {1'b0, layer_2_0[4415:4408]};
      btm_1[0] = {1'b0,layer_3_1[4399:4392]} - {1'b0, layer_2_1[4399:4392]};
      btm_1[1] = {1'b0,layer_3_1[4407:4400]} - {1'b0, layer_2_1[4407:4400]};
      btm_1[2] = {1'b0,layer_3_1[4415:4408]} - {1'b0, layer_2_1[4415:4408]};
      btm_2[0] = {1'b0,layer_3_2[4399:4392]} - {1'b0, layer_2_2[4399:4392]};
      btm_2[1] = {1'b0,layer_3_2[4407:4400]} - {1'b0, layer_2_2[4407:4400]};
      btm_2[2] = {1'b0,layer_3_2[4415:4408]} - {1'b0, layer_2_2[4415:4408]};
    end
    'd551: begin
      top_0[0] = {1'b0,layer_1_0[4407:4400]} - {1'b0, layer_0_0[4407:4400]};
      top_0[1] = {1'b0,layer_1_0[4415:4408]} - {1'b0, layer_0_0[4415:4408]};
      top_0[2] = {1'b0,layer_1_0[4423:4416]} - {1'b0, layer_0_0[4423:4416]};
      top_1[0] = {1'b0,layer_1_1[4407:4400]} - {1'b0, layer_0_1[4407:4400]};
      top_1[1] = {1'b0,layer_1_1[4415:4408]} - {1'b0, layer_0_1[4415:4408]};
      top_1[2] = {1'b0,layer_1_1[4423:4416]} - {1'b0, layer_0_1[4423:4416]};
      top_2[0] = {1'b0,layer_1_2[4407:4400]} - {1'b0, layer_0_2[4407:4400]};
      top_2[1] = {1'b0,layer_1_2[4415:4408]} - {1'b0, layer_0_2[4415:4408]};
      top_2[2] = {1'b0,layer_1_2[4423:4416]} - {1'b0, layer_0_2[4423:4416]};
      mid_0[0] = {1'b0,layer_2_0[4407:4400]} - {1'b0, layer_1_0[4407:4400]};
      mid_0[1] = {1'b0,layer_2_0[4415:4408]} - {1'b0, layer_1_0[4415:4408]};
      mid_0[2] = {1'b0,layer_2_0[4423:4416]} - {1'b0, layer_1_0[4423:4416]};
      mid_1[0] = {1'b0,layer_2_1[4407:4400]} - {1'b0, layer_1_1[4407:4400]};
      mid_1[1] = {1'b0,layer_2_1[4415:4408]} - {1'b0, layer_1_1[4415:4408]};
      mid_1[2] = {1'b0,layer_2_1[4423:4416]} - {1'b0, layer_1_1[4423:4416]};
      mid_2[0] = {1'b0,layer_2_2[4407:4400]} - {1'b0, layer_1_2[4407:4400]};
      mid_2[1] = {1'b0,layer_2_2[4415:4408]} - {1'b0, layer_1_2[4415:4408]};
      mid_2[2] = {1'b0,layer_2_2[4423:4416]} - {1'b0, layer_1_2[4423:4416]};
      btm_0[0] = {1'b0,layer_3_0[4407:4400]} - {1'b0, layer_2_0[4407:4400]};
      btm_0[1] = {1'b0,layer_3_0[4415:4408]} - {1'b0, layer_2_0[4415:4408]};
      btm_0[2] = {1'b0,layer_3_0[4423:4416]} - {1'b0, layer_2_0[4423:4416]};
      btm_1[0] = {1'b0,layer_3_1[4407:4400]} - {1'b0, layer_2_1[4407:4400]};
      btm_1[1] = {1'b0,layer_3_1[4415:4408]} - {1'b0, layer_2_1[4415:4408]};
      btm_1[2] = {1'b0,layer_3_1[4423:4416]} - {1'b0, layer_2_1[4423:4416]};
      btm_2[0] = {1'b0,layer_3_2[4407:4400]} - {1'b0, layer_2_2[4407:4400]};
      btm_2[1] = {1'b0,layer_3_2[4415:4408]} - {1'b0, layer_2_2[4415:4408]};
      btm_2[2] = {1'b0,layer_3_2[4423:4416]} - {1'b0, layer_2_2[4423:4416]};
    end
    'd552: begin
      top_0[0] = {1'b0,layer_1_0[4415:4408]} - {1'b0, layer_0_0[4415:4408]};
      top_0[1] = {1'b0,layer_1_0[4423:4416]} - {1'b0, layer_0_0[4423:4416]};
      top_0[2] = {1'b0,layer_1_0[4431:4424]} - {1'b0, layer_0_0[4431:4424]};
      top_1[0] = {1'b0,layer_1_1[4415:4408]} - {1'b0, layer_0_1[4415:4408]};
      top_1[1] = {1'b0,layer_1_1[4423:4416]} - {1'b0, layer_0_1[4423:4416]};
      top_1[2] = {1'b0,layer_1_1[4431:4424]} - {1'b0, layer_0_1[4431:4424]};
      top_2[0] = {1'b0,layer_1_2[4415:4408]} - {1'b0, layer_0_2[4415:4408]};
      top_2[1] = {1'b0,layer_1_2[4423:4416]} - {1'b0, layer_0_2[4423:4416]};
      top_2[2] = {1'b0,layer_1_2[4431:4424]} - {1'b0, layer_0_2[4431:4424]};
      mid_0[0] = {1'b0,layer_2_0[4415:4408]} - {1'b0, layer_1_0[4415:4408]};
      mid_0[1] = {1'b0,layer_2_0[4423:4416]} - {1'b0, layer_1_0[4423:4416]};
      mid_0[2] = {1'b0,layer_2_0[4431:4424]} - {1'b0, layer_1_0[4431:4424]};
      mid_1[0] = {1'b0,layer_2_1[4415:4408]} - {1'b0, layer_1_1[4415:4408]};
      mid_1[1] = {1'b0,layer_2_1[4423:4416]} - {1'b0, layer_1_1[4423:4416]};
      mid_1[2] = {1'b0,layer_2_1[4431:4424]} - {1'b0, layer_1_1[4431:4424]};
      mid_2[0] = {1'b0,layer_2_2[4415:4408]} - {1'b0, layer_1_2[4415:4408]};
      mid_2[1] = {1'b0,layer_2_2[4423:4416]} - {1'b0, layer_1_2[4423:4416]};
      mid_2[2] = {1'b0,layer_2_2[4431:4424]} - {1'b0, layer_1_2[4431:4424]};
      btm_0[0] = {1'b0,layer_3_0[4415:4408]} - {1'b0, layer_2_0[4415:4408]};
      btm_0[1] = {1'b0,layer_3_0[4423:4416]} - {1'b0, layer_2_0[4423:4416]};
      btm_0[2] = {1'b0,layer_3_0[4431:4424]} - {1'b0, layer_2_0[4431:4424]};
      btm_1[0] = {1'b0,layer_3_1[4415:4408]} - {1'b0, layer_2_1[4415:4408]};
      btm_1[1] = {1'b0,layer_3_1[4423:4416]} - {1'b0, layer_2_1[4423:4416]};
      btm_1[2] = {1'b0,layer_3_1[4431:4424]} - {1'b0, layer_2_1[4431:4424]};
      btm_2[0] = {1'b0,layer_3_2[4415:4408]} - {1'b0, layer_2_2[4415:4408]};
      btm_2[1] = {1'b0,layer_3_2[4423:4416]} - {1'b0, layer_2_2[4423:4416]};
      btm_2[2] = {1'b0,layer_3_2[4431:4424]} - {1'b0, layer_2_2[4431:4424]};
    end
    'd553: begin
      top_0[0] = {1'b0,layer_1_0[4423:4416]} - {1'b0, layer_0_0[4423:4416]};
      top_0[1] = {1'b0,layer_1_0[4431:4424]} - {1'b0, layer_0_0[4431:4424]};
      top_0[2] = {1'b0,layer_1_0[4439:4432]} - {1'b0, layer_0_0[4439:4432]};
      top_1[0] = {1'b0,layer_1_1[4423:4416]} - {1'b0, layer_0_1[4423:4416]};
      top_1[1] = {1'b0,layer_1_1[4431:4424]} - {1'b0, layer_0_1[4431:4424]};
      top_1[2] = {1'b0,layer_1_1[4439:4432]} - {1'b0, layer_0_1[4439:4432]};
      top_2[0] = {1'b0,layer_1_2[4423:4416]} - {1'b0, layer_0_2[4423:4416]};
      top_2[1] = {1'b0,layer_1_2[4431:4424]} - {1'b0, layer_0_2[4431:4424]};
      top_2[2] = {1'b0,layer_1_2[4439:4432]} - {1'b0, layer_0_2[4439:4432]};
      mid_0[0] = {1'b0,layer_2_0[4423:4416]} - {1'b0, layer_1_0[4423:4416]};
      mid_0[1] = {1'b0,layer_2_0[4431:4424]} - {1'b0, layer_1_0[4431:4424]};
      mid_0[2] = {1'b0,layer_2_0[4439:4432]} - {1'b0, layer_1_0[4439:4432]};
      mid_1[0] = {1'b0,layer_2_1[4423:4416]} - {1'b0, layer_1_1[4423:4416]};
      mid_1[1] = {1'b0,layer_2_1[4431:4424]} - {1'b0, layer_1_1[4431:4424]};
      mid_1[2] = {1'b0,layer_2_1[4439:4432]} - {1'b0, layer_1_1[4439:4432]};
      mid_2[0] = {1'b0,layer_2_2[4423:4416]} - {1'b0, layer_1_2[4423:4416]};
      mid_2[1] = {1'b0,layer_2_2[4431:4424]} - {1'b0, layer_1_2[4431:4424]};
      mid_2[2] = {1'b0,layer_2_2[4439:4432]} - {1'b0, layer_1_2[4439:4432]};
      btm_0[0] = {1'b0,layer_3_0[4423:4416]} - {1'b0, layer_2_0[4423:4416]};
      btm_0[1] = {1'b0,layer_3_0[4431:4424]} - {1'b0, layer_2_0[4431:4424]};
      btm_0[2] = {1'b0,layer_3_0[4439:4432]} - {1'b0, layer_2_0[4439:4432]};
      btm_1[0] = {1'b0,layer_3_1[4423:4416]} - {1'b0, layer_2_1[4423:4416]};
      btm_1[1] = {1'b0,layer_3_1[4431:4424]} - {1'b0, layer_2_1[4431:4424]};
      btm_1[2] = {1'b0,layer_3_1[4439:4432]} - {1'b0, layer_2_1[4439:4432]};
      btm_2[0] = {1'b0,layer_3_2[4423:4416]} - {1'b0, layer_2_2[4423:4416]};
      btm_2[1] = {1'b0,layer_3_2[4431:4424]} - {1'b0, layer_2_2[4431:4424]};
      btm_2[2] = {1'b0,layer_3_2[4439:4432]} - {1'b0, layer_2_2[4439:4432]};
    end
    'd554: begin
      top_0[0] = {1'b0,layer_1_0[4431:4424]} - {1'b0, layer_0_0[4431:4424]};
      top_0[1] = {1'b0,layer_1_0[4439:4432]} - {1'b0, layer_0_0[4439:4432]};
      top_0[2] = {1'b0,layer_1_0[4447:4440]} - {1'b0, layer_0_0[4447:4440]};
      top_1[0] = {1'b0,layer_1_1[4431:4424]} - {1'b0, layer_0_1[4431:4424]};
      top_1[1] = {1'b0,layer_1_1[4439:4432]} - {1'b0, layer_0_1[4439:4432]};
      top_1[2] = {1'b0,layer_1_1[4447:4440]} - {1'b0, layer_0_1[4447:4440]};
      top_2[0] = {1'b0,layer_1_2[4431:4424]} - {1'b0, layer_0_2[4431:4424]};
      top_2[1] = {1'b0,layer_1_2[4439:4432]} - {1'b0, layer_0_2[4439:4432]};
      top_2[2] = {1'b0,layer_1_2[4447:4440]} - {1'b0, layer_0_2[4447:4440]};
      mid_0[0] = {1'b0,layer_2_0[4431:4424]} - {1'b0, layer_1_0[4431:4424]};
      mid_0[1] = {1'b0,layer_2_0[4439:4432]} - {1'b0, layer_1_0[4439:4432]};
      mid_0[2] = {1'b0,layer_2_0[4447:4440]} - {1'b0, layer_1_0[4447:4440]};
      mid_1[0] = {1'b0,layer_2_1[4431:4424]} - {1'b0, layer_1_1[4431:4424]};
      mid_1[1] = {1'b0,layer_2_1[4439:4432]} - {1'b0, layer_1_1[4439:4432]};
      mid_1[2] = {1'b0,layer_2_1[4447:4440]} - {1'b0, layer_1_1[4447:4440]};
      mid_2[0] = {1'b0,layer_2_2[4431:4424]} - {1'b0, layer_1_2[4431:4424]};
      mid_2[1] = {1'b0,layer_2_2[4439:4432]} - {1'b0, layer_1_2[4439:4432]};
      mid_2[2] = {1'b0,layer_2_2[4447:4440]} - {1'b0, layer_1_2[4447:4440]};
      btm_0[0] = {1'b0,layer_3_0[4431:4424]} - {1'b0, layer_2_0[4431:4424]};
      btm_0[1] = {1'b0,layer_3_0[4439:4432]} - {1'b0, layer_2_0[4439:4432]};
      btm_0[2] = {1'b0,layer_3_0[4447:4440]} - {1'b0, layer_2_0[4447:4440]};
      btm_1[0] = {1'b0,layer_3_1[4431:4424]} - {1'b0, layer_2_1[4431:4424]};
      btm_1[1] = {1'b0,layer_3_1[4439:4432]} - {1'b0, layer_2_1[4439:4432]};
      btm_1[2] = {1'b0,layer_3_1[4447:4440]} - {1'b0, layer_2_1[4447:4440]};
      btm_2[0] = {1'b0,layer_3_2[4431:4424]} - {1'b0, layer_2_2[4431:4424]};
      btm_2[1] = {1'b0,layer_3_2[4439:4432]} - {1'b0, layer_2_2[4439:4432]};
      btm_2[2] = {1'b0,layer_3_2[4447:4440]} - {1'b0, layer_2_2[4447:4440]};
    end
    'd555: begin
      top_0[0] = {1'b0,layer_1_0[4439:4432]} - {1'b0, layer_0_0[4439:4432]};
      top_0[1] = {1'b0,layer_1_0[4447:4440]} - {1'b0, layer_0_0[4447:4440]};
      top_0[2] = {1'b0,layer_1_0[4455:4448]} - {1'b0, layer_0_0[4455:4448]};
      top_1[0] = {1'b0,layer_1_1[4439:4432]} - {1'b0, layer_0_1[4439:4432]};
      top_1[1] = {1'b0,layer_1_1[4447:4440]} - {1'b0, layer_0_1[4447:4440]};
      top_1[2] = {1'b0,layer_1_1[4455:4448]} - {1'b0, layer_0_1[4455:4448]};
      top_2[0] = {1'b0,layer_1_2[4439:4432]} - {1'b0, layer_0_2[4439:4432]};
      top_2[1] = {1'b0,layer_1_2[4447:4440]} - {1'b0, layer_0_2[4447:4440]};
      top_2[2] = {1'b0,layer_1_2[4455:4448]} - {1'b0, layer_0_2[4455:4448]};
      mid_0[0] = {1'b0,layer_2_0[4439:4432]} - {1'b0, layer_1_0[4439:4432]};
      mid_0[1] = {1'b0,layer_2_0[4447:4440]} - {1'b0, layer_1_0[4447:4440]};
      mid_0[2] = {1'b0,layer_2_0[4455:4448]} - {1'b0, layer_1_0[4455:4448]};
      mid_1[0] = {1'b0,layer_2_1[4439:4432]} - {1'b0, layer_1_1[4439:4432]};
      mid_1[1] = {1'b0,layer_2_1[4447:4440]} - {1'b0, layer_1_1[4447:4440]};
      mid_1[2] = {1'b0,layer_2_1[4455:4448]} - {1'b0, layer_1_1[4455:4448]};
      mid_2[0] = {1'b0,layer_2_2[4439:4432]} - {1'b0, layer_1_2[4439:4432]};
      mid_2[1] = {1'b0,layer_2_2[4447:4440]} - {1'b0, layer_1_2[4447:4440]};
      mid_2[2] = {1'b0,layer_2_2[4455:4448]} - {1'b0, layer_1_2[4455:4448]};
      btm_0[0] = {1'b0,layer_3_0[4439:4432]} - {1'b0, layer_2_0[4439:4432]};
      btm_0[1] = {1'b0,layer_3_0[4447:4440]} - {1'b0, layer_2_0[4447:4440]};
      btm_0[2] = {1'b0,layer_3_0[4455:4448]} - {1'b0, layer_2_0[4455:4448]};
      btm_1[0] = {1'b0,layer_3_1[4439:4432]} - {1'b0, layer_2_1[4439:4432]};
      btm_1[1] = {1'b0,layer_3_1[4447:4440]} - {1'b0, layer_2_1[4447:4440]};
      btm_1[2] = {1'b0,layer_3_1[4455:4448]} - {1'b0, layer_2_1[4455:4448]};
      btm_2[0] = {1'b0,layer_3_2[4439:4432]} - {1'b0, layer_2_2[4439:4432]};
      btm_2[1] = {1'b0,layer_3_2[4447:4440]} - {1'b0, layer_2_2[4447:4440]};
      btm_2[2] = {1'b0,layer_3_2[4455:4448]} - {1'b0, layer_2_2[4455:4448]};
    end
    'd556: begin
      top_0[0] = {1'b0,layer_1_0[4447:4440]} - {1'b0, layer_0_0[4447:4440]};
      top_0[1] = {1'b0,layer_1_0[4455:4448]} - {1'b0, layer_0_0[4455:4448]};
      top_0[2] = {1'b0,layer_1_0[4463:4456]} - {1'b0, layer_0_0[4463:4456]};
      top_1[0] = {1'b0,layer_1_1[4447:4440]} - {1'b0, layer_0_1[4447:4440]};
      top_1[1] = {1'b0,layer_1_1[4455:4448]} - {1'b0, layer_0_1[4455:4448]};
      top_1[2] = {1'b0,layer_1_1[4463:4456]} - {1'b0, layer_0_1[4463:4456]};
      top_2[0] = {1'b0,layer_1_2[4447:4440]} - {1'b0, layer_0_2[4447:4440]};
      top_2[1] = {1'b0,layer_1_2[4455:4448]} - {1'b0, layer_0_2[4455:4448]};
      top_2[2] = {1'b0,layer_1_2[4463:4456]} - {1'b0, layer_0_2[4463:4456]};
      mid_0[0] = {1'b0,layer_2_0[4447:4440]} - {1'b0, layer_1_0[4447:4440]};
      mid_0[1] = {1'b0,layer_2_0[4455:4448]} - {1'b0, layer_1_0[4455:4448]};
      mid_0[2] = {1'b0,layer_2_0[4463:4456]} - {1'b0, layer_1_0[4463:4456]};
      mid_1[0] = {1'b0,layer_2_1[4447:4440]} - {1'b0, layer_1_1[4447:4440]};
      mid_1[1] = {1'b0,layer_2_1[4455:4448]} - {1'b0, layer_1_1[4455:4448]};
      mid_1[2] = {1'b0,layer_2_1[4463:4456]} - {1'b0, layer_1_1[4463:4456]};
      mid_2[0] = {1'b0,layer_2_2[4447:4440]} - {1'b0, layer_1_2[4447:4440]};
      mid_2[1] = {1'b0,layer_2_2[4455:4448]} - {1'b0, layer_1_2[4455:4448]};
      mid_2[2] = {1'b0,layer_2_2[4463:4456]} - {1'b0, layer_1_2[4463:4456]};
      btm_0[0] = {1'b0,layer_3_0[4447:4440]} - {1'b0, layer_2_0[4447:4440]};
      btm_0[1] = {1'b0,layer_3_0[4455:4448]} - {1'b0, layer_2_0[4455:4448]};
      btm_0[2] = {1'b0,layer_3_0[4463:4456]} - {1'b0, layer_2_0[4463:4456]};
      btm_1[0] = {1'b0,layer_3_1[4447:4440]} - {1'b0, layer_2_1[4447:4440]};
      btm_1[1] = {1'b0,layer_3_1[4455:4448]} - {1'b0, layer_2_1[4455:4448]};
      btm_1[2] = {1'b0,layer_3_1[4463:4456]} - {1'b0, layer_2_1[4463:4456]};
      btm_2[0] = {1'b0,layer_3_2[4447:4440]} - {1'b0, layer_2_2[4447:4440]};
      btm_2[1] = {1'b0,layer_3_2[4455:4448]} - {1'b0, layer_2_2[4455:4448]};
      btm_2[2] = {1'b0,layer_3_2[4463:4456]} - {1'b0, layer_2_2[4463:4456]};
    end
    'd557: begin
      top_0[0] = {1'b0,layer_1_0[4455:4448]} - {1'b0, layer_0_0[4455:4448]};
      top_0[1] = {1'b0,layer_1_0[4463:4456]} - {1'b0, layer_0_0[4463:4456]};
      top_0[2] = {1'b0,layer_1_0[4471:4464]} - {1'b0, layer_0_0[4471:4464]};
      top_1[0] = {1'b0,layer_1_1[4455:4448]} - {1'b0, layer_0_1[4455:4448]};
      top_1[1] = {1'b0,layer_1_1[4463:4456]} - {1'b0, layer_0_1[4463:4456]};
      top_1[2] = {1'b0,layer_1_1[4471:4464]} - {1'b0, layer_0_1[4471:4464]};
      top_2[0] = {1'b0,layer_1_2[4455:4448]} - {1'b0, layer_0_2[4455:4448]};
      top_2[1] = {1'b0,layer_1_2[4463:4456]} - {1'b0, layer_0_2[4463:4456]};
      top_2[2] = {1'b0,layer_1_2[4471:4464]} - {1'b0, layer_0_2[4471:4464]};
      mid_0[0] = {1'b0,layer_2_0[4455:4448]} - {1'b0, layer_1_0[4455:4448]};
      mid_0[1] = {1'b0,layer_2_0[4463:4456]} - {1'b0, layer_1_0[4463:4456]};
      mid_0[2] = {1'b0,layer_2_0[4471:4464]} - {1'b0, layer_1_0[4471:4464]};
      mid_1[0] = {1'b0,layer_2_1[4455:4448]} - {1'b0, layer_1_1[4455:4448]};
      mid_1[1] = {1'b0,layer_2_1[4463:4456]} - {1'b0, layer_1_1[4463:4456]};
      mid_1[2] = {1'b0,layer_2_1[4471:4464]} - {1'b0, layer_1_1[4471:4464]};
      mid_2[0] = {1'b0,layer_2_2[4455:4448]} - {1'b0, layer_1_2[4455:4448]};
      mid_2[1] = {1'b0,layer_2_2[4463:4456]} - {1'b0, layer_1_2[4463:4456]};
      mid_2[2] = {1'b0,layer_2_2[4471:4464]} - {1'b0, layer_1_2[4471:4464]};
      btm_0[0] = {1'b0,layer_3_0[4455:4448]} - {1'b0, layer_2_0[4455:4448]};
      btm_0[1] = {1'b0,layer_3_0[4463:4456]} - {1'b0, layer_2_0[4463:4456]};
      btm_0[2] = {1'b0,layer_3_0[4471:4464]} - {1'b0, layer_2_0[4471:4464]};
      btm_1[0] = {1'b0,layer_3_1[4455:4448]} - {1'b0, layer_2_1[4455:4448]};
      btm_1[1] = {1'b0,layer_3_1[4463:4456]} - {1'b0, layer_2_1[4463:4456]};
      btm_1[2] = {1'b0,layer_3_1[4471:4464]} - {1'b0, layer_2_1[4471:4464]};
      btm_2[0] = {1'b0,layer_3_2[4455:4448]} - {1'b0, layer_2_2[4455:4448]};
      btm_2[1] = {1'b0,layer_3_2[4463:4456]} - {1'b0, layer_2_2[4463:4456]};
      btm_2[2] = {1'b0,layer_3_2[4471:4464]} - {1'b0, layer_2_2[4471:4464]};
    end
    'd558: begin
      top_0[0] = {1'b0,layer_1_0[4463:4456]} - {1'b0, layer_0_0[4463:4456]};
      top_0[1] = {1'b0,layer_1_0[4471:4464]} - {1'b0, layer_0_0[4471:4464]};
      top_0[2] = {1'b0,layer_1_0[4479:4472]} - {1'b0, layer_0_0[4479:4472]};
      top_1[0] = {1'b0,layer_1_1[4463:4456]} - {1'b0, layer_0_1[4463:4456]};
      top_1[1] = {1'b0,layer_1_1[4471:4464]} - {1'b0, layer_0_1[4471:4464]};
      top_1[2] = {1'b0,layer_1_1[4479:4472]} - {1'b0, layer_0_1[4479:4472]};
      top_2[0] = {1'b0,layer_1_2[4463:4456]} - {1'b0, layer_0_2[4463:4456]};
      top_2[1] = {1'b0,layer_1_2[4471:4464]} - {1'b0, layer_0_2[4471:4464]};
      top_2[2] = {1'b0,layer_1_2[4479:4472]} - {1'b0, layer_0_2[4479:4472]};
      mid_0[0] = {1'b0,layer_2_0[4463:4456]} - {1'b0, layer_1_0[4463:4456]};
      mid_0[1] = {1'b0,layer_2_0[4471:4464]} - {1'b0, layer_1_0[4471:4464]};
      mid_0[2] = {1'b0,layer_2_0[4479:4472]} - {1'b0, layer_1_0[4479:4472]};
      mid_1[0] = {1'b0,layer_2_1[4463:4456]} - {1'b0, layer_1_1[4463:4456]};
      mid_1[1] = {1'b0,layer_2_1[4471:4464]} - {1'b0, layer_1_1[4471:4464]};
      mid_1[2] = {1'b0,layer_2_1[4479:4472]} - {1'b0, layer_1_1[4479:4472]};
      mid_2[0] = {1'b0,layer_2_2[4463:4456]} - {1'b0, layer_1_2[4463:4456]};
      mid_2[1] = {1'b0,layer_2_2[4471:4464]} - {1'b0, layer_1_2[4471:4464]};
      mid_2[2] = {1'b0,layer_2_2[4479:4472]} - {1'b0, layer_1_2[4479:4472]};
      btm_0[0] = {1'b0,layer_3_0[4463:4456]} - {1'b0, layer_2_0[4463:4456]};
      btm_0[1] = {1'b0,layer_3_0[4471:4464]} - {1'b0, layer_2_0[4471:4464]};
      btm_0[2] = {1'b0,layer_3_0[4479:4472]} - {1'b0, layer_2_0[4479:4472]};
      btm_1[0] = {1'b0,layer_3_1[4463:4456]} - {1'b0, layer_2_1[4463:4456]};
      btm_1[1] = {1'b0,layer_3_1[4471:4464]} - {1'b0, layer_2_1[4471:4464]};
      btm_1[2] = {1'b0,layer_3_1[4479:4472]} - {1'b0, layer_2_1[4479:4472]};
      btm_2[0] = {1'b0,layer_3_2[4463:4456]} - {1'b0, layer_2_2[4463:4456]};
      btm_2[1] = {1'b0,layer_3_2[4471:4464]} - {1'b0, layer_2_2[4471:4464]};
      btm_2[2] = {1'b0,layer_3_2[4479:4472]} - {1'b0, layer_2_2[4479:4472]};
    end
    'd559: begin
      top_0[0] = {1'b0,layer_1_0[4471:4464]} - {1'b0, layer_0_0[4471:4464]};
      top_0[1] = {1'b0,layer_1_0[4479:4472]} - {1'b0, layer_0_0[4479:4472]};
      top_0[2] = {1'b0,layer_1_0[4487:4480]} - {1'b0, layer_0_0[4487:4480]};
      top_1[0] = {1'b0,layer_1_1[4471:4464]} - {1'b0, layer_0_1[4471:4464]};
      top_1[1] = {1'b0,layer_1_1[4479:4472]} - {1'b0, layer_0_1[4479:4472]};
      top_1[2] = {1'b0,layer_1_1[4487:4480]} - {1'b0, layer_0_1[4487:4480]};
      top_2[0] = {1'b0,layer_1_2[4471:4464]} - {1'b0, layer_0_2[4471:4464]};
      top_2[1] = {1'b0,layer_1_2[4479:4472]} - {1'b0, layer_0_2[4479:4472]};
      top_2[2] = {1'b0,layer_1_2[4487:4480]} - {1'b0, layer_0_2[4487:4480]};
      mid_0[0] = {1'b0,layer_2_0[4471:4464]} - {1'b0, layer_1_0[4471:4464]};
      mid_0[1] = {1'b0,layer_2_0[4479:4472]} - {1'b0, layer_1_0[4479:4472]};
      mid_0[2] = {1'b0,layer_2_0[4487:4480]} - {1'b0, layer_1_0[4487:4480]};
      mid_1[0] = {1'b0,layer_2_1[4471:4464]} - {1'b0, layer_1_1[4471:4464]};
      mid_1[1] = {1'b0,layer_2_1[4479:4472]} - {1'b0, layer_1_1[4479:4472]};
      mid_1[2] = {1'b0,layer_2_1[4487:4480]} - {1'b0, layer_1_1[4487:4480]};
      mid_2[0] = {1'b0,layer_2_2[4471:4464]} - {1'b0, layer_1_2[4471:4464]};
      mid_2[1] = {1'b0,layer_2_2[4479:4472]} - {1'b0, layer_1_2[4479:4472]};
      mid_2[2] = {1'b0,layer_2_2[4487:4480]} - {1'b0, layer_1_2[4487:4480]};
      btm_0[0] = {1'b0,layer_3_0[4471:4464]} - {1'b0, layer_2_0[4471:4464]};
      btm_0[1] = {1'b0,layer_3_0[4479:4472]} - {1'b0, layer_2_0[4479:4472]};
      btm_0[2] = {1'b0,layer_3_0[4487:4480]} - {1'b0, layer_2_0[4487:4480]};
      btm_1[0] = {1'b0,layer_3_1[4471:4464]} - {1'b0, layer_2_1[4471:4464]};
      btm_1[1] = {1'b0,layer_3_1[4479:4472]} - {1'b0, layer_2_1[4479:4472]};
      btm_1[2] = {1'b0,layer_3_1[4487:4480]} - {1'b0, layer_2_1[4487:4480]};
      btm_2[0] = {1'b0,layer_3_2[4471:4464]} - {1'b0, layer_2_2[4471:4464]};
      btm_2[1] = {1'b0,layer_3_2[4479:4472]} - {1'b0, layer_2_2[4479:4472]};
      btm_2[2] = {1'b0,layer_3_2[4487:4480]} - {1'b0, layer_2_2[4487:4480]};
    end
    'd560: begin
      top_0[0] = {1'b0,layer_1_0[4479:4472]} - {1'b0, layer_0_0[4479:4472]};
      top_0[1] = {1'b0,layer_1_0[4487:4480]} - {1'b0, layer_0_0[4487:4480]};
      top_0[2] = {1'b0,layer_1_0[4495:4488]} - {1'b0, layer_0_0[4495:4488]};
      top_1[0] = {1'b0,layer_1_1[4479:4472]} - {1'b0, layer_0_1[4479:4472]};
      top_1[1] = {1'b0,layer_1_1[4487:4480]} - {1'b0, layer_0_1[4487:4480]};
      top_1[2] = {1'b0,layer_1_1[4495:4488]} - {1'b0, layer_0_1[4495:4488]};
      top_2[0] = {1'b0,layer_1_2[4479:4472]} - {1'b0, layer_0_2[4479:4472]};
      top_2[1] = {1'b0,layer_1_2[4487:4480]} - {1'b0, layer_0_2[4487:4480]};
      top_2[2] = {1'b0,layer_1_2[4495:4488]} - {1'b0, layer_0_2[4495:4488]};
      mid_0[0] = {1'b0,layer_2_0[4479:4472]} - {1'b0, layer_1_0[4479:4472]};
      mid_0[1] = {1'b0,layer_2_0[4487:4480]} - {1'b0, layer_1_0[4487:4480]};
      mid_0[2] = {1'b0,layer_2_0[4495:4488]} - {1'b0, layer_1_0[4495:4488]};
      mid_1[0] = {1'b0,layer_2_1[4479:4472]} - {1'b0, layer_1_1[4479:4472]};
      mid_1[1] = {1'b0,layer_2_1[4487:4480]} - {1'b0, layer_1_1[4487:4480]};
      mid_1[2] = {1'b0,layer_2_1[4495:4488]} - {1'b0, layer_1_1[4495:4488]};
      mid_2[0] = {1'b0,layer_2_2[4479:4472]} - {1'b0, layer_1_2[4479:4472]};
      mid_2[1] = {1'b0,layer_2_2[4487:4480]} - {1'b0, layer_1_2[4487:4480]};
      mid_2[2] = {1'b0,layer_2_2[4495:4488]} - {1'b0, layer_1_2[4495:4488]};
      btm_0[0] = {1'b0,layer_3_0[4479:4472]} - {1'b0, layer_2_0[4479:4472]};
      btm_0[1] = {1'b0,layer_3_0[4487:4480]} - {1'b0, layer_2_0[4487:4480]};
      btm_0[2] = {1'b0,layer_3_0[4495:4488]} - {1'b0, layer_2_0[4495:4488]};
      btm_1[0] = {1'b0,layer_3_1[4479:4472]} - {1'b0, layer_2_1[4479:4472]};
      btm_1[1] = {1'b0,layer_3_1[4487:4480]} - {1'b0, layer_2_1[4487:4480]};
      btm_1[2] = {1'b0,layer_3_1[4495:4488]} - {1'b0, layer_2_1[4495:4488]};
      btm_2[0] = {1'b0,layer_3_2[4479:4472]} - {1'b0, layer_2_2[4479:4472]};
      btm_2[1] = {1'b0,layer_3_2[4487:4480]} - {1'b0, layer_2_2[4487:4480]};
      btm_2[2] = {1'b0,layer_3_2[4495:4488]} - {1'b0, layer_2_2[4495:4488]};
    end
    'd561: begin
      top_0[0] = {1'b0,layer_1_0[4487:4480]} - {1'b0, layer_0_0[4487:4480]};
      top_0[1] = {1'b0,layer_1_0[4495:4488]} - {1'b0, layer_0_0[4495:4488]};
      top_0[2] = {1'b0,layer_1_0[4503:4496]} - {1'b0, layer_0_0[4503:4496]};
      top_1[0] = {1'b0,layer_1_1[4487:4480]} - {1'b0, layer_0_1[4487:4480]};
      top_1[1] = {1'b0,layer_1_1[4495:4488]} - {1'b0, layer_0_1[4495:4488]};
      top_1[2] = {1'b0,layer_1_1[4503:4496]} - {1'b0, layer_0_1[4503:4496]};
      top_2[0] = {1'b0,layer_1_2[4487:4480]} - {1'b0, layer_0_2[4487:4480]};
      top_2[1] = {1'b0,layer_1_2[4495:4488]} - {1'b0, layer_0_2[4495:4488]};
      top_2[2] = {1'b0,layer_1_2[4503:4496]} - {1'b0, layer_0_2[4503:4496]};
      mid_0[0] = {1'b0,layer_2_0[4487:4480]} - {1'b0, layer_1_0[4487:4480]};
      mid_0[1] = {1'b0,layer_2_0[4495:4488]} - {1'b0, layer_1_0[4495:4488]};
      mid_0[2] = {1'b0,layer_2_0[4503:4496]} - {1'b0, layer_1_0[4503:4496]};
      mid_1[0] = {1'b0,layer_2_1[4487:4480]} - {1'b0, layer_1_1[4487:4480]};
      mid_1[1] = {1'b0,layer_2_1[4495:4488]} - {1'b0, layer_1_1[4495:4488]};
      mid_1[2] = {1'b0,layer_2_1[4503:4496]} - {1'b0, layer_1_1[4503:4496]};
      mid_2[0] = {1'b0,layer_2_2[4487:4480]} - {1'b0, layer_1_2[4487:4480]};
      mid_2[1] = {1'b0,layer_2_2[4495:4488]} - {1'b0, layer_1_2[4495:4488]};
      mid_2[2] = {1'b0,layer_2_2[4503:4496]} - {1'b0, layer_1_2[4503:4496]};
      btm_0[0] = {1'b0,layer_3_0[4487:4480]} - {1'b0, layer_2_0[4487:4480]};
      btm_0[1] = {1'b0,layer_3_0[4495:4488]} - {1'b0, layer_2_0[4495:4488]};
      btm_0[2] = {1'b0,layer_3_0[4503:4496]} - {1'b0, layer_2_0[4503:4496]};
      btm_1[0] = {1'b0,layer_3_1[4487:4480]} - {1'b0, layer_2_1[4487:4480]};
      btm_1[1] = {1'b0,layer_3_1[4495:4488]} - {1'b0, layer_2_1[4495:4488]};
      btm_1[2] = {1'b0,layer_3_1[4503:4496]} - {1'b0, layer_2_1[4503:4496]};
      btm_2[0] = {1'b0,layer_3_2[4487:4480]} - {1'b0, layer_2_2[4487:4480]};
      btm_2[1] = {1'b0,layer_3_2[4495:4488]} - {1'b0, layer_2_2[4495:4488]};
      btm_2[2] = {1'b0,layer_3_2[4503:4496]} - {1'b0, layer_2_2[4503:4496]};
    end
    'd562: begin
      top_0[0] = {1'b0,layer_1_0[4495:4488]} - {1'b0, layer_0_0[4495:4488]};
      top_0[1] = {1'b0,layer_1_0[4503:4496]} - {1'b0, layer_0_0[4503:4496]};
      top_0[2] = {1'b0,layer_1_0[4511:4504]} - {1'b0, layer_0_0[4511:4504]};
      top_1[0] = {1'b0,layer_1_1[4495:4488]} - {1'b0, layer_0_1[4495:4488]};
      top_1[1] = {1'b0,layer_1_1[4503:4496]} - {1'b0, layer_0_1[4503:4496]};
      top_1[2] = {1'b0,layer_1_1[4511:4504]} - {1'b0, layer_0_1[4511:4504]};
      top_2[0] = {1'b0,layer_1_2[4495:4488]} - {1'b0, layer_0_2[4495:4488]};
      top_2[1] = {1'b0,layer_1_2[4503:4496]} - {1'b0, layer_0_2[4503:4496]};
      top_2[2] = {1'b0,layer_1_2[4511:4504]} - {1'b0, layer_0_2[4511:4504]};
      mid_0[0] = {1'b0,layer_2_0[4495:4488]} - {1'b0, layer_1_0[4495:4488]};
      mid_0[1] = {1'b0,layer_2_0[4503:4496]} - {1'b0, layer_1_0[4503:4496]};
      mid_0[2] = {1'b0,layer_2_0[4511:4504]} - {1'b0, layer_1_0[4511:4504]};
      mid_1[0] = {1'b0,layer_2_1[4495:4488]} - {1'b0, layer_1_1[4495:4488]};
      mid_1[1] = {1'b0,layer_2_1[4503:4496]} - {1'b0, layer_1_1[4503:4496]};
      mid_1[2] = {1'b0,layer_2_1[4511:4504]} - {1'b0, layer_1_1[4511:4504]};
      mid_2[0] = {1'b0,layer_2_2[4495:4488]} - {1'b0, layer_1_2[4495:4488]};
      mid_2[1] = {1'b0,layer_2_2[4503:4496]} - {1'b0, layer_1_2[4503:4496]};
      mid_2[2] = {1'b0,layer_2_2[4511:4504]} - {1'b0, layer_1_2[4511:4504]};
      btm_0[0] = {1'b0,layer_3_0[4495:4488]} - {1'b0, layer_2_0[4495:4488]};
      btm_0[1] = {1'b0,layer_3_0[4503:4496]} - {1'b0, layer_2_0[4503:4496]};
      btm_0[2] = {1'b0,layer_3_0[4511:4504]} - {1'b0, layer_2_0[4511:4504]};
      btm_1[0] = {1'b0,layer_3_1[4495:4488]} - {1'b0, layer_2_1[4495:4488]};
      btm_1[1] = {1'b0,layer_3_1[4503:4496]} - {1'b0, layer_2_1[4503:4496]};
      btm_1[2] = {1'b0,layer_3_1[4511:4504]} - {1'b0, layer_2_1[4511:4504]};
      btm_2[0] = {1'b0,layer_3_2[4495:4488]} - {1'b0, layer_2_2[4495:4488]};
      btm_2[1] = {1'b0,layer_3_2[4503:4496]} - {1'b0, layer_2_2[4503:4496]};
      btm_2[2] = {1'b0,layer_3_2[4511:4504]} - {1'b0, layer_2_2[4511:4504]};
    end
    'd563: begin
      top_0[0] = {1'b0,layer_1_0[4503:4496]} - {1'b0, layer_0_0[4503:4496]};
      top_0[1] = {1'b0,layer_1_0[4511:4504]} - {1'b0, layer_0_0[4511:4504]};
      top_0[2] = {1'b0,layer_1_0[4519:4512]} - {1'b0, layer_0_0[4519:4512]};
      top_1[0] = {1'b0,layer_1_1[4503:4496]} - {1'b0, layer_0_1[4503:4496]};
      top_1[1] = {1'b0,layer_1_1[4511:4504]} - {1'b0, layer_0_1[4511:4504]};
      top_1[2] = {1'b0,layer_1_1[4519:4512]} - {1'b0, layer_0_1[4519:4512]};
      top_2[0] = {1'b0,layer_1_2[4503:4496]} - {1'b0, layer_0_2[4503:4496]};
      top_2[1] = {1'b0,layer_1_2[4511:4504]} - {1'b0, layer_0_2[4511:4504]};
      top_2[2] = {1'b0,layer_1_2[4519:4512]} - {1'b0, layer_0_2[4519:4512]};
      mid_0[0] = {1'b0,layer_2_0[4503:4496]} - {1'b0, layer_1_0[4503:4496]};
      mid_0[1] = {1'b0,layer_2_0[4511:4504]} - {1'b0, layer_1_0[4511:4504]};
      mid_0[2] = {1'b0,layer_2_0[4519:4512]} - {1'b0, layer_1_0[4519:4512]};
      mid_1[0] = {1'b0,layer_2_1[4503:4496]} - {1'b0, layer_1_1[4503:4496]};
      mid_1[1] = {1'b0,layer_2_1[4511:4504]} - {1'b0, layer_1_1[4511:4504]};
      mid_1[2] = {1'b0,layer_2_1[4519:4512]} - {1'b0, layer_1_1[4519:4512]};
      mid_2[0] = {1'b0,layer_2_2[4503:4496]} - {1'b0, layer_1_2[4503:4496]};
      mid_2[1] = {1'b0,layer_2_2[4511:4504]} - {1'b0, layer_1_2[4511:4504]};
      mid_2[2] = {1'b0,layer_2_2[4519:4512]} - {1'b0, layer_1_2[4519:4512]};
      btm_0[0] = {1'b0,layer_3_0[4503:4496]} - {1'b0, layer_2_0[4503:4496]};
      btm_0[1] = {1'b0,layer_3_0[4511:4504]} - {1'b0, layer_2_0[4511:4504]};
      btm_0[2] = {1'b0,layer_3_0[4519:4512]} - {1'b0, layer_2_0[4519:4512]};
      btm_1[0] = {1'b0,layer_3_1[4503:4496]} - {1'b0, layer_2_1[4503:4496]};
      btm_1[1] = {1'b0,layer_3_1[4511:4504]} - {1'b0, layer_2_1[4511:4504]};
      btm_1[2] = {1'b0,layer_3_1[4519:4512]} - {1'b0, layer_2_1[4519:4512]};
      btm_2[0] = {1'b0,layer_3_2[4503:4496]} - {1'b0, layer_2_2[4503:4496]};
      btm_2[1] = {1'b0,layer_3_2[4511:4504]} - {1'b0, layer_2_2[4511:4504]};
      btm_2[2] = {1'b0,layer_3_2[4519:4512]} - {1'b0, layer_2_2[4519:4512]};
    end
    'd564: begin
      top_0[0] = {1'b0,layer_1_0[4511:4504]} - {1'b0, layer_0_0[4511:4504]};
      top_0[1] = {1'b0,layer_1_0[4519:4512]} - {1'b0, layer_0_0[4519:4512]};
      top_0[2] = {1'b0,layer_1_0[4527:4520]} - {1'b0, layer_0_0[4527:4520]};
      top_1[0] = {1'b0,layer_1_1[4511:4504]} - {1'b0, layer_0_1[4511:4504]};
      top_1[1] = {1'b0,layer_1_1[4519:4512]} - {1'b0, layer_0_1[4519:4512]};
      top_1[2] = {1'b0,layer_1_1[4527:4520]} - {1'b0, layer_0_1[4527:4520]};
      top_2[0] = {1'b0,layer_1_2[4511:4504]} - {1'b0, layer_0_2[4511:4504]};
      top_2[1] = {1'b0,layer_1_2[4519:4512]} - {1'b0, layer_0_2[4519:4512]};
      top_2[2] = {1'b0,layer_1_2[4527:4520]} - {1'b0, layer_0_2[4527:4520]};
      mid_0[0] = {1'b0,layer_2_0[4511:4504]} - {1'b0, layer_1_0[4511:4504]};
      mid_0[1] = {1'b0,layer_2_0[4519:4512]} - {1'b0, layer_1_0[4519:4512]};
      mid_0[2] = {1'b0,layer_2_0[4527:4520]} - {1'b0, layer_1_0[4527:4520]};
      mid_1[0] = {1'b0,layer_2_1[4511:4504]} - {1'b0, layer_1_1[4511:4504]};
      mid_1[1] = {1'b0,layer_2_1[4519:4512]} - {1'b0, layer_1_1[4519:4512]};
      mid_1[2] = {1'b0,layer_2_1[4527:4520]} - {1'b0, layer_1_1[4527:4520]};
      mid_2[0] = {1'b0,layer_2_2[4511:4504]} - {1'b0, layer_1_2[4511:4504]};
      mid_2[1] = {1'b0,layer_2_2[4519:4512]} - {1'b0, layer_1_2[4519:4512]};
      mid_2[2] = {1'b0,layer_2_2[4527:4520]} - {1'b0, layer_1_2[4527:4520]};
      btm_0[0] = {1'b0,layer_3_0[4511:4504]} - {1'b0, layer_2_0[4511:4504]};
      btm_0[1] = {1'b0,layer_3_0[4519:4512]} - {1'b0, layer_2_0[4519:4512]};
      btm_0[2] = {1'b0,layer_3_0[4527:4520]} - {1'b0, layer_2_0[4527:4520]};
      btm_1[0] = {1'b0,layer_3_1[4511:4504]} - {1'b0, layer_2_1[4511:4504]};
      btm_1[1] = {1'b0,layer_3_1[4519:4512]} - {1'b0, layer_2_1[4519:4512]};
      btm_1[2] = {1'b0,layer_3_1[4527:4520]} - {1'b0, layer_2_1[4527:4520]};
      btm_2[0] = {1'b0,layer_3_2[4511:4504]} - {1'b0, layer_2_2[4511:4504]};
      btm_2[1] = {1'b0,layer_3_2[4519:4512]} - {1'b0, layer_2_2[4519:4512]};
      btm_2[2] = {1'b0,layer_3_2[4527:4520]} - {1'b0, layer_2_2[4527:4520]};
    end
    'd565: begin
      top_0[0] = {1'b0,layer_1_0[4519:4512]} - {1'b0, layer_0_0[4519:4512]};
      top_0[1] = {1'b0,layer_1_0[4527:4520]} - {1'b0, layer_0_0[4527:4520]};
      top_0[2] = {1'b0,layer_1_0[4535:4528]} - {1'b0, layer_0_0[4535:4528]};
      top_1[0] = {1'b0,layer_1_1[4519:4512]} - {1'b0, layer_0_1[4519:4512]};
      top_1[1] = {1'b0,layer_1_1[4527:4520]} - {1'b0, layer_0_1[4527:4520]};
      top_1[2] = {1'b0,layer_1_1[4535:4528]} - {1'b0, layer_0_1[4535:4528]};
      top_2[0] = {1'b0,layer_1_2[4519:4512]} - {1'b0, layer_0_2[4519:4512]};
      top_2[1] = {1'b0,layer_1_2[4527:4520]} - {1'b0, layer_0_2[4527:4520]};
      top_2[2] = {1'b0,layer_1_2[4535:4528]} - {1'b0, layer_0_2[4535:4528]};
      mid_0[0] = {1'b0,layer_2_0[4519:4512]} - {1'b0, layer_1_0[4519:4512]};
      mid_0[1] = {1'b0,layer_2_0[4527:4520]} - {1'b0, layer_1_0[4527:4520]};
      mid_0[2] = {1'b0,layer_2_0[4535:4528]} - {1'b0, layer_1_0[4535:4528]};
      mid_1[0] = {1'b0,layer_2_1[4519:4512]} - {1'b0, layer_1_1[4519:4512]};
      mid_1[1] = {1'b0,layer_2_1[4527:4520]} - {1'b0, layer_1_1[4527:4520]};
      mid_1[2] = {1'b0,layer_2_1[4535:4528]} - {1'b0, layer_1_1[4535:4528]};
      mid_2[0] = {1'b0,layer_2_2[4519:4512]} - {1'b0, layer_1_2[4519:4512]};
      mid_2[1] = {1'b0,layer_2_2[4527:4520]} - {1'b0, layer_1_2[4527:4520]};
      mid_2[2] = {1'b0,layer_2_2[4535:4528]} - {1'b0, layer_1_2[4535:4528]};
      btm_0[0] = {1'b0,layer_3_0[4519:4512]} - {1'b0, layer_2_0[4519:4512]};
      btm_0[1] = {1'b0,layer_3_0[4527:4520]} - {1'b0, layer_2_0[4527:4520]};
      btm_0[2] = {1'b0,layer_3_0[4535:4528]} - {1'b0, layer_2_0[4535:4528]};
      btm_1[0] = {1'b0,layer_3_1[4519:4512]} - {1'b0, layer_2_1[4519:4512]};
      btm_1[1] = {1'b0,layer_3_1[4527:4520]} - {1'b0, layer_2_1[4527:4520]};
      btm_1[2] = {1'b0,layer_3_1[4535:4528]} - {1'b0, layer_2_1[4535:4528]};
      btm_2[0] = {1'b0,layer_3_2[4519:4512]} - {1'b0, layer_2_2[4519:4512]};
      btm_2[1] = {1'b0,layer_3_2[4527:4520]} - {1'b0, layer_2_2[4527:4520]};
      btm_2[2] = {1'b0,layer_3_2[4535:4528]} - {1'b0, layer_2_2[4535:4528]};
    end
    'd566: begin
      top_0[0] = {1'b0,layer_1_0[4527:4520]} - {1'b0, layer_0_0[4527:4520]};
      top_0[1] = {1'b0,layer_1_0[4535:4528]} - {1'b0, layer_0_0[4535:4528]};
      top_0[2] = {1'b0,layer_1_0[4543:4536]} - {1'b0, layer_0_0[4543:4536]};
      top_1[0] = {1'b0,layer_1_1[4527:4520]} - {1'b0, layer_0_1[4527:4520]};
      top_1[1] = {1'b0,layer_1_1[4535:4528]} - {1'b0, layer_0_1[4535:4528]};
      top_1[2] = {1'b0,layer_1_1[4543:4536]} - {1'b0, layer_0_1[4543:4536]};
      top_2[0] = {1'b0,layer_1_2[4527:4520]} - {1'b0, layer_0_2[4527:4520]};
      top_2[1] = {1'b0,layer_1_2[4535:4528]} - {1'b0, layer_0_2[4535:4528]};
      top_2[2] = {1'b0,layer_1_2[4543:4536]} - {1'b0, layer_0_2[4543:4536]};
      mid_0[0] = {1'b0,layer_2_0[4527:4520]} - {1'b0, layer_1_0[4527:4520]};
      mid_0[1] = {1'b0,layer_2_0[4535:4528]} - {1'b0, layer_1_0[4535:4528]};
      mid_0[2] = {1'b0,layer_2_0[4543:4536]} - {1'b0, layer_1_0[4543:4536]};
      mid_1[0] = {1'b0,layer_2_1[4527:4520]} - {1'b0, layer_1_1[4527:4520]};
      mid_1[1] = {1'b0,layer_2_1[4535:4528]} - {1'b0, layer_1_1[4535:4528]};
      mid_1[2] = {1'b0,layer_2_1[4543:4536]} - {1'b0, layer_1_1[4543:4536]};
      mid_2[0] = {1'b0,layer_2_2[4527:4520]} - {1'b0, layer_1_2[4527:4520]};
      mid_2[1] = {1'b0,layer_2_2[4535:4528]} - {1'b0, layer_1_2[4535:4528]};
      mid_2[2] = {1'b0,layer_2_2[4543:4536]} - {1'b0, layer_1_2[4543:4536]};
      btm_0[0] = {1'b0,layer_3_0[4527:4520]} - {1'b0, layer_2_0[4527:4520]};
      btm_0[1] = {1'b0,layer_3_0[4535:4528]} - {1'b0, layer_2_0[4535:4528]};
      btm_0[2] = {1'b0,layer_3_0[4543:4536]} - {1'b0, layer_2_0[4543:4536]};
      btm_1[0] = {1'b0,layer_3_1[4527:4520]} - {1'b0, layer_2_1[4527:4520]};
      btm_1[1] = {1'b0,layer_3_1[4535:4528]} - {1'b0, layer_2_1[4535:4528]};
      btm_1[2] = {1'b0,layer_3_1[4543:4536]} - {1'b0, layer_2_1[4543:4536]};
      btm_2[0] = {1'b0,layer_3_2[4527:4520]} - {1'b0, layer_2_2[4527:4520]};
      btm_2[1] = {1'b0,layer_3_2[4535:4528]} - {1'b0, layer_2_2[4535:4528]};
      btm_2[2] = {1'b0,layer_3_2[4543:4536]} - {1'b0, layer_2_2[4543:4536]};
    end
    'd567: begin
      top_0[0] = {1'b0,layer_1_0[4535:4528]} - {1'b0, layer_0_0[4535:4528]};
      top_0[1] = {1'b0,layer_1_0[4543:4536]} - {1'b0, layer_0_0[4543:4536]};
      top_0[2] = {1'b0,layer_1_0[4551:4544]} - {1'b0, layer_0_0[4551:4544]};
      top_1[0] = {1'b0,layer_1_1[4535:4528]} - {1'b0, layer_0_1[4535:4528]};
      top_1[1] = {1'b0,layer_1_1[4543:4536]} - {1'b0, layer_0_1[4543:4536]};
      top_1[2] = {1'b0,layer_1_1[4551:4544]} - {1'b0, layer_0_1[4551:4544]};
      top_2[0] = {1'b0,layer_1_2[4535:4528]} - {1'b0, layer_0_2[4535:4528]};
      top_2[1] = {1'b0,layer_1_2[4543:4536]} - {1'b0, layer_0_2[4543:4536]};
      top_2[2] = {1'b0,layer_1_2[4551:4544]} - {1'b0, layer_0_2[4551:4544]};
      mid_0[0] = {1'b0,layer_2_0[4535:4528]} - {1'b0, layer_1_0[4535:4528]};
      mid_0[1] = {1'b0,layer_2_0[4543:4536]} - {1'b0, layer_1_0[4543:4536]};
      mid_0[2] = {1'b0,layer_2_0[4551:4544]} - {1'b0, layer_1_0[4551:4544]};
      mid_1[0] = {1'b0,layer_2_1[4535:4528]} - {1'b0, layer_1_1[4535:4528]};
      mid_1[1] = {1'b0,layer_2_1[4543:4536]} - {1'b0, layer_1_1[4543:4536]};
      mid_1[2] = {1'b0,layer_2_1[4551:4544]} - {1'b0, layer_1_1[4551:4544]};
      mid_2[0] = {1'b0,layer_2_2[4535:4528]} - {1'b0, layer_1_2[4535:4528]};
      mid_2[1] = {1'b0,layer_2_2[4543:4536]} - {1'b0, layer_1_2[4543:4536]};
      mid_2[2] = {1'b0,layer_2_2[4551:4544]} - {1'b0, layer_1_2[4551:4544]};
      btm_0[0] = {1'b0,layer_3_0[4535:4528]} - {1'b0, layer_2_0[4535:4528]};
      btm_0[1] = {1'b0,layer_3_0[4543:4536]} - {1'b0, layer_2_0[4543:4536]};
      btm_0[2] = {1'b0,layer_3_0[4551:4544]} - {1'b0, layer_2_0[4551:4544]};
      btm_1[0] = {1'b0,layer_3_1[4535:4528]} - {1'b0, layer_2_1[4535:4528]};
      btm_1[1] = {1'b0,layer_3_1[4543:4536]} - {1'b0, layer_2_1[4543:4536]};
      btm_1[2] = {1'b0,layer_3_1[4551:4544]} - {1'b0, layer_2_1[4551:4544]};
      btm_2[0] = {1'b0,layer_3_2[4535:4528]} - {1'b0, layer_2_2[4535:4528]};
      btm_2[1] = {1'b0,layer_3_2[4543:4536]} - {1'b0, layer_2_2[4543:4536]};
      btm_2[2] = {1'b0,layer_3_2[4551:4544]} - {1'b0, layer_2_2[4551:4544]};
    end
    'd568: begin
      top_0[0] = {1'b0,layer_1_0[4543:4536]} - {1'b0, layer_0_0[4543:4536]};
      top_0[1] = {1'b0,layer_1_0[4551:4544]} - {1'b0, layer_0_0[4551:4544]};
      top_0[2] = {1'b0,layer_1_0[4559:4552]} - {1'b0, layer_0_0[4559:4552]};
      top_1[0] = {1'b0,layer_1_1[4543:4536]} - {1'b0, layer_0_1[4543:4536]};
      top_1[1] = {1'b0,layer_1_1[4551:4544]} - {1'b0, layer_0_1[4551:4544]};
      top_1[2] = {1'b0,layer_1_1[4559:4552]} - {1'b0, layer_0_1[4559:4552]};
      top_2[0] = {1'b0,layer_1_2[4543:4536]} - {1'b0, layer_0_2[4543:4536]};
      top_2[1] = {1'b0,layer_1_2[4551:4544]} - {1'b0, layer_0_2[4551:4544]};
      top_2[2] = {1'b0,layer_1_2[4559:4552]} - {1'b0, layer_0_2[4559:4552]};
      mid_0[0] = {1'b0,layer_2_0[4543:4536]} - {1'b0, layer_1_0[4543:4536]};
      mid_0[1] = {1'b0,layer_2_0[4551:4544]} - {1'b0, layer_1_0[4551:4544]};
      mid_0[2] = {1'b0,layer_2_0[4559:4552]} - {1'b0, layer_1_0[4559:4552]};
      mid_1[0] = {1'b0,layer_2_1[4543:4536]} - {1'b0, layer_1_1[4543:4536]};
      mid_1[1] = {1'b0,layer_2_1[4551:4544]} - {1'b0, layer_1_1[4551:4544]};
      mid_1[2] = {1'b0,layer_2_1[4559:4552]} - {1'b0, layer_1_1[4559:4552]};
      mid_2[0] = {1'b0,layer_2_2[4543:4536]} - {1'b0, layer_1_2[4543:4536]};
      mid_2[1] = {1'b0,layer_2_2[4551:4544]} - {1'b0, layer_1_2[4551:4544]};
      mid_2[2] = {1'b0,layer_2_2[4559:4552]} - {1'b0, layer_1_2[4559:4552]};
      btm_0[0] = {1'b0,layer_3_0[4543:4536]} - {1'b0, layer_2_0[4543:4536]};
      btm_0[1] = {1'b0,layer_3_0[4551:4544]} - {1'b0, layer_2_0[4551:4544]};
      btm_0[2] = {1'b0,layer_3_0[4559:4552]} - {1'b0, layer_2_0[4559:4552]};
      btm_1[0] = {1'b0,layer_3_1[4543:4536]} - {1'b0, layer_2_1[4543:4536]};
      btm_1[1] = {1'b0,layer_3_1[4551:4544]} - {1'b0, layer_2_1[4551:4544]};
      btm_1[2] = {1'b0,layer_3_1[4559:4552]} - {1'b0, layer_2_1[4559:4552]};
      btm_2[0] = {1'b0,layer_3_2[4543:4536]} - {1'b0, layer_2_2[4543:4536]};
      btm_2[1] = {1'b0,layer_3_2[4551:4544]} - {1'b0, layer_2_2[4551:4544]};
      btm_2[2] = {1'b0,layer_3_2[4559:4552]} - {1'b0, layer_2_2[4559:4552]};
    end
    'd569: begin
      top_0[0] = {1'b0,layer_1_0[4551:4544]} - {1'b0, layer_0_0[4551:4544]};
      top_0[1] = {1'b0,layer_1_0[4559:4552]} - {1'b0, layer_0_0[4559:4552]};
      top_0[2] = {1'b0,layer_1_0[4567:4560]} - {1'b0, layer_0_0[4567:4560]};
      top_1[0] = {1'b0,layer_1_1[4551:4544]} - {1'b0, layer_0_1[4551:4544]};
      top_1[1] = {1'b0,layer_1_1[4559:4552]} - {1'b0, layer_0_1[4559:4552]};
      top_1[2] = {1'b0,layer_1_1[4567:4560]} - {1'b0, layer_0_1[4567:4560]};
      top_2[0] = {1'b0,layer_1_2[4551:4544]} - {1'b0, layer_0_2[4551:4544]};
      top_2[1] = {1'b0,layer_1_2[4559:4552]} - {1'b0, layer_0_2[4559:4552]};
      top_2[2] = {1'b0,layer_1_2[4567:4560]} - {1'b0, layer_0_2[4567:4560]};
      mid_0[0] = {1'b0,layer_2_0[4551:4544]} - {1'b0, layer_1_0[4551:4544]};
      mid_0[1] = {1'b0,layer_2_0[4559:4552]} - {1'b0, layer_1_0[4559:4552]};
      mid_0[2] = {1'b0,layer_2_0[4567:4560]} - {1'b0, layer_1_0[4567:4560]};
      mid_1[0] = {1'b0,layer_2_1[4551:4544]} - {1'b0, layer_1_1[4551:4544]};
      mid_1[1] = {1'b0,layer_2_1[4559:4552]} - {1'b0, layer_1_1[4559:4552]};
      mid_1[2] = {1'b0,layer_2_1[4567:4560]} - {1'b0, layer_1_1[4567:4560]};
      mid_2[0] = {1'b0,layer_2_2[4551:4544]} - {1'b0, layer_1_2[4551:4544]};
      mid_2[1] = {1'b0,layer_2_2[4559:4552]} - {1'b0, layer_1_2[4559:4552]};
      mid_2[2] = {1'b0,layer_2_2[4567:4560]} - {1'b0, layer_1_2[4567:4560]};
      btm_0[0] = {1'b0,layer_3_0[4551:4544]} - {1'b0, layer_2_0[4551:4544]};
      btm_0[1] = {1'b0,layer_3_0[4559:4552]} - {1'b0, layer_2_0[4559:4552]};
      btm_0[2] = {1'b0,layer_3_0[4567:4560]} - {1'b0, layer_2_0[4567:4560]};
      btm_1[0] = {1'b0,layer_3_1[4551:4544]} - {1'b0, layer_2_1[4551:4544]};
      btm_1[1] = {1'b0,layer_3_1[4559:4552]} - {1'b0, layer_2_1[4559:4552]};
      btm_1[2] = {1'b0,layer_3_1[4567:4560]} - {1'b0, layer_2_1[4567:4560]};
      btm_2[0] = {1'b0,layer_3_2[4551:4544]} - {1'b0, layer_2_2[4551:4544]};
      btm_2[1] = {1'b0,layer_3_2[4559:4552]} - {1'b0, layer_2_2[4559:4552]};
      btm_2[2] = {1'b0,layer_3_2[4567:4560]} - {1'b0, layer_2_2[4567:4560]};
    end
    'd570: begin
      top_0[0] = {1'b0,layer_1_0[4559:4552]} - {1'b0, layer_0_0[4559:4552]};
      top_0[1] = {1'b0,layer_1_0[4567:4560]} - {1'b0, layer_0_0[4567:4560]};
      top_0[2] = {1'b0,layer_1_0[4575:4568]} - {1'b0, layer_0_0[4575:4568]};
      top_1[0] = {1'b0,layer_1_1[4559:4552]} - {1'b0, layer_0_1[4559:4552]};
      top_1[1] = {1'b0,layer_1_1[4567:4560]} - {1'b0, layer_0_1[4567:4560]};
      top_1[2] = {1'b0,layer_1_1[4575:4568]} - {1'b0, layer_0_1[4575:4568]};
      top_2[0] = {1'b0,layer_1_2[4559:4552]} - {1'b0, layer_0_2[4559:4552]};
      top_2[1] = {1'b0,layer_1_2[4567:4560]} - {1'b0, layer_0_2[4567:4560]};
      top_2[2] = {1'b0,layer_1_2[4575:4568]} - {1'b0, layer_0_2[4575:4568]};
      mid_0[0] = {1'b0,layer_2_0[4559:4552]} - {1'b0, layer_1_0[4559:4552]};
      mid_0[1] = {1'b0,layer_2_0[4567:4560]} - {1'b0, layer_1_0[4567:4560]};
      mid_0[2] = {1'b0,layer_2_0[4575:4568]} - {1'b0, layer_1_0[4575:4568]};
      mid_1[0] = {1'b0,layer_2_1[4559:4552]} - {1'b0, layer_1_1[4559:4552]};
      mid_1[1] = {1'b0,layer_2_1[4567:4560]} - {1'b0, layer_1_1[4567:4560]};
      mid_1[2] = {1'b0,layer_2_1[4575:4568]} - {1'b0, layer_1_1[4575:4568]};
      mid_2[0] = {1'b0,layer_2_2[4559:4552]} - {1'b0, layer_1_2[4559:4552]};
      mid_2[1] = {1'b0,layer_2_2[4567:4560]} - {1'b0, layer_1_2[4567:4560]};
      mid_2[2] = {1'b0,layer_2_2[4575:4568]} - {1'b0, layer_1_2[4575:4568]};
      btm_0[0] = {1'b0,layer_3_0[4559:4552]} - {1'b0, layer_2_0[4559:4552]};
      btm_0[1] = {1'b0,layer_3_0[4567:4560]} - {1'b0, layer_2_0[4567:4560]};
      btm_0[2] = {1'b0,layer_3_0[4575:4568]} - {1'b0, layer_2_0[4575:4568]};
      btm_1[0] = {1'b0,layer_3_1[4559:4552]} - {1'b0, layer_2_1[4559:4552]};
      btm_1[1] = {1'b0,layer_3_1[4567:4560]} - {1'b0, layer_2_1[4567:4560]};
      btm_1[2] = {1'b0,layer_3_1[4575:4568]} - {1'b0, layer_2_1[4575:4568]};
      btm_2[0] = {1'b0,layer_3_2[4559:4552]} - {1'b0, layer_2_2[4559:4552]};
      btm_2[1] = {1'b0,layer_3_2[4567:4560]} - {1'b0, layer_2_2[4567:4560]};
      btm_2[2] = {1'b0,layer_3_2[4575:4568]} - {1'b0, layer_2_2[4575:4568]};
    end
    'd571: begin
      top_0[0] = {1'b0,layer_1_0[4567:4560]} - {1'b0, layer_0_0[4567:4560]};
      top_0[1] = {1'b0,layer_1_0[4575:4568]} - {1'b0, layer_0_0[4575:4568]};
      top_0[2] = {1'b0,layer_1_0[4583:4576]} - {1'b0, layer_0_0[4583:4576]};
      top_1[0] = {1'b0,layer_1_1[4567:4560]} - {1'b0, layer_0_1[4567:4560]};
      top_1[1] = {1'b0,layer_1_1[4575:4568]} - {1'b0, layer_0_1[4575:4568]};
      top_1[2] = {1'b0,layer_1_1[4583:4576]} - {1'b0, layer_0_1[4583:4576]};
      top_2[0] = {1'b0,layer_1_2[4567:4560]} - {1'b0, layer_0_2[4567:4560]};
      top_2[1] = {1'b0,layer_1_2[4575:4568]} - {1'b0, layer_0_2[4575:4568]};
      top_2[2] = {1'b0,layer_1_2[4583:4576]} - {1'b0, layer_0_2[4583:4576]};
      mid_0[0] = {1'b0,layer_2_0[4567:4560]} - {1'b0, layer_1_0[4567:4560]};
      mid_0[1] = {1'b0,layer_2_0[4575:4568]} - {1'b0, layer_1_0[4575:4568]};
      mid_0[2] = {1'b0,layer_2_0[4583:4576]} - {1'b0, layer_1_0[4583:4576]};
      mid_1[0] = {1'b0,layer_2_1[4567:4560]} - {1'b0, layer_1_1[4567:4560]};
      mid_1[1] = {1'b0,layer_2_1[4575:4568]} - {1'b0, layer_1_1[4575:4568]};
      mid_1[2] = {1'b0,layer_2_1[4583:4576]} - {1'b0, layer_1_1[4583:4576]};
      mid_2[0] = {1'b0,layer_2_2[4567:4560]} - {1'b0, layer_1_2[4567:4560]};
      mid_2[1] = {1'b0,layer_2_2[4575:4568]} - {1'b0, layer_1_2[4575:4568]};
      mid_2[2] = {1'b0,layer_2_2[4583:4576]} - {1'b0, layer_1_2[4583:4576]};
      btm_0[0] = {1'b0,layer_3_0[4567:4560]} - {1'b0, layer_2_0[4567:4560]};
      btm_0[1] = {1'b0,layer_3_0[4575:4568]} - {1'b0, layer_2_0[4575:4568]};
      btm_0[2] = {1'b0,layer_3_0[4583:4576]} - {1'b0, layer_2_0[4583:4576]};
      btm_1[0] = {1'b0,layer_3_1[4567:4560]} - {1'b0, layer_2_1[4567:4560]};
      btm_1[1] = {1'b0,layer_3_1[4575:4568]} - {1'b0, layer_2_1[4575:4568]};
      btm_1[2] = {1'b0,layer_3_1[4583:4576]} - {1'b0, layer_2_1[4583:4576]};
      btm_2[0] = {1'b0,layer_3_2[4567:4560]} - {1'b0, layer_2_2[4567:4560]};
      btm_2[1] = {1'b0,layer_3_2[4575:4568]} - {1'b0, layer_2_2[4575:4568]};
      btm_2[2] = {1'b0,layer_3_2[4583:4576]} - {1'b0, layer_2_2[4583:4576]};
    end
    'd572: begin
      top_0[0] = {1'b0,layer_1_0[4575:4568]} - {1'b0, layer_0_0[4575:4568]};
      top_0[1] = {1'b0,layer_1_0[4583:4576]} - {1'b0, layer_0_0[4583:4576]};
      top_0[2] = {1'b0,layer_1_0[4591:4584]} - {1'b0, layer_0_0[4591:4584]};
      top_1[0] = {1'b0,layer_1_1[4575:4568]} - {1'b0, layer_0_1[4575:4568]};
      top_1[1] = {1'b0,layer_1_1[4583:4576]} - {1'b0, layer_0_1[4583:4576]};
      top_1[2] = {1'b0,layer_1_1[4591:4584]} - {1'b0, layer_0_1[4591:4584]};
      top_2[0] = {1'b0,layer_1_2[4575:4568]} - {1'b0, layer_0_2[4575:4568]};
      top_2[1] = {1'b0,layer_1_2[4583:4576]} - {1'b0, layer_0_2[4583:4576]};
      top_2[2] = {1'b0,layer_1_2[4591:4584]} - {1'b0, layer_0_2[4591:4584]};
      mid_0[0] = {1'b0,layer_2_0[4575:4568]} - {1'b0, layer_1_0[4575:4568]};
      mid_0[1] = {1'b0,layer_2_0[4583:4576]} - {1'b0, layer_1_0[4583:4576]};
      mid_0[2] = {1'b0,layer_2_0[4591:4584]} - {1'b0, layer_1_0[4591:4584]};
      mid_1[0] = {1'b0,layer_2_1[4575:4568]} - {1'b0, layer_1_1[4575:4568]};
      mid_1[1] = {1'b0,layer_2_1[4583:4576]} - {1'b0, layer_1_1[4583:4576]};
      mid_1[2] = {1'b0,layer_2_1[4591:4584]} - {1'b0, layer_1_1[4591:4584]};
      mid_2[0] = {1'b0,layer_2_2[4575:4568]} - {1'b0, layer_1_2[4575:4568]};
      mid_2[1] = {1'b0,layer_2_2[4583:4576]} - {1'b0, layer_1_2[4583:4576]};
      mid_2[2] = {1'b0,layer_2_2[4591:4584]} - {1'b0, layer_1_2[4591:4584]};
      btm_0[0] = {1'b0,layer_3_0[4575:4568]} - {1'b0, layer_2_0[4575:4568]};
      btm_0[1] = {1'b0,layer_3_0[4583:4576]} - {1'b0, layer_2_0[4583:4576]};
      btm_0[2] = {1'b0,layer_3_0[4591:4584]} - {1'b0, layer_2_0[4591:4584]};
      btm_1[0] = {1'b0,layer_3_1[4575:4568]} - {1'b0, layer_2_1[4575:4568]};
      btm_1[1] = {1'b0,layer_3_1[4583:4576]} - {1'b0, layer_2_1[4583:4576]};
      btm_1[2] = {1'b0,layer_3_1[4591:4584]} - {1'b0, layer_2_1[4591:4584]};
      btm_2[0] = {1'b0,layer_3_2[4575:4568]} - {1'b0, layer_2_2[4575:4568]};
      btm_2[1] = {1'b0,layer_3_2[4583:4576]} - {1'b0, layer_2_2[4583:4576]};
      btm_2[2] = {1'b0,layer_3_2[4591:4584]} - {1'b0, layer_2_2[4591:4584]};
    end
    'd573: begin
      top_0[0] = {1'b0,layer_1_0[4583:4576]} - {1'b0, layer_0_0[4583:4576]};
      top_0[1] = {1'b0,layer_1_0[4591:4584]} - {1'b0, layer_0_0[4591:4584]};
      top_0[2] = {1'b0,layer_1_0[4599:4592]} - {1'b0, layer_0_0[4599:4592]};
      top_1[0] = {1'b0,layer_1_1[4583:4576]} - {1'b0, layer_0_1[4583:4576]};
      top_1[1] = {1'b0,layer_1_1[4591:4584]} - {1'b0, layer_0_1[4591:4584]};
      top_1[2] = {1'b0,layer_1_1[4599:4592]} - {1'b0, layer_0_1[4599:4592]};
      top_2[0] = {1'b0,layer_1_2[4583:4576]} - {1'b0, layer_0_2[4583:4576]};
      top_2[1] = {1'b0,layer_1_2[4591:4584]} - {1'b0, layer_0_2[4591:4584]};
      top_2[2] = {1'b0,layer_1_2[4599:4592]} - {1'b0, layer_0_2[4599:4592]};
      mid_0[0] = {1'b0,layer_2_0[4583:4576]} - {1'b0, layer_1_0[4583:4576]};
      mid_0[1] = {1'b0,layer_2_0[4591:4584]} - {1'b0, layer_1_0[4591:4584]};
      mid_0[2] = {1'b0,layer_2_0[4599:4592]} - {1'b0, layer_1_0[4599:4592]};
      mid_1[0] = {1'b0,layer_2_1[4583:4576]} - {1'b0, layer_1_1[4583:4576]};
      mid_1[1] = {1'b0,layer_2_1[4591:4584]} - {1'b0, layer_1_1[4591:4584]};
      mid_1[2] = {1'b0,layer_2_1[4599:4592]} - {1'b0, layer_1_1[4599:4592]};
      mid_2[0] = {1'b0,layer_2_2[4583:4576]} - {1'b0, layer_1_2[4583:4576]};
      mid_2[1] = {1'b0,layer_2_2[4591:4584]} - {1'b0, layer_1_2[4591:4584]};
      mid_2[2] = {1'b0,layer_2_2[4599:4592]} - {1'b0, layer_1_2[4599:4592]};
      btm_0[0] = {1'b0,layer_3_0[4583:4576]} - {1'b0, layer_2_0[4583:4576]};
      btm_0[1] = {1'b0,layer_3_0[4591:4584]} - {1'b0, layer_2_0[4591:4584]};
      btm_0[2] = {1'b0,layer_3_0[4599:4592]} - {1'b0, layer_2_0[4599:4592]};
      btm_1[0] = {1'b0,layer_3_1[4583:4576]} - {1'b0, layer_2_1[4583:4576]};
      btm_1[1] = {1'b0,layer_3_1[4591:4584]} - {1'b0, layer_2_1[4591:4584]};
      btm_1[2] = {1'b0,layer_3_1[4599:4592]} - {1'b0, layer_2_1[4599:4592]};
      btm_2[0] = {1'b0,layer_3_2[4583:4576]} - {1'b0, layer_2_2[4583:4576]};
      btm_2[1] = {1'b0,layer_3_2[4591:4584]} - {1'b0, layer_2_2[4591:4584]};
      btm_2[2] = {1'b0,layer_3_2[4599:4592]} - {1'b0, layer_2_2[4599:4592]};
    end
    'd574: begin
      top_0[0] = {1'b0,layer_1_0[4591:4584]} - {1'b0, layer_0_0[4591:4584]};
      top_0[1] = {1'b0,layer_1_0[4599:4592]} - {1'b0, layer_0_0[4599:4592]};
      top_0[2] = {1'b0,layer_1_0[4607:4600]} - {1'b0, layer_0_0[4607:4600]};
      top_1[0] = {1'b0,layer_1_1[4591:4584]} - {1'b0, layer_0_1[4591:4584]};
      top_1[1] = {1'b0,layer_1_1[4599:4592]} - {1'b0, layer_0_1[4599:4592]};
      top_1[2] = {1'b0,layer_1_1[4607:4600]} - {1'b0, layer_0_1[4607:4600]};
      top_2[0] = {1'b0,layer_1_2[4591:4584]} - {1'b0, layer_0_2[4591:4584]};
      top_2[1] = {1'b0,layer_1_2[4599:4592]} - {1'b0, layer_0_2[4599:4592]};
      top_2[2] = {1'b0,layer_1_2[4607:4600]} - {1'b0, layer_0_2[4607:4600]};
      mid_0[0] = {1'b0,layer_2_0[4591:4584]} - {1'b0, layer_1_0[4591:4584]};
      mid_0[1] = {1'b0,layer_2_0[4599:4592]} - {1'b0, layer_1_0[4599:4592]};
      mid_0[2] = {1'b0,layer_2_0[4607:4600]} - {1'b0, layer_1_0[4607:4600]};
      mid_1[0] = {1'b0,layer_2_1[4591:4584]} - {1'b0, layer_1_1[4591:4584]};
      mid_1[1] = {1'b0,layer_2_1[4599:4592]} - {1'b0, layer_1_1[4599:4592]};
      mid_1[2] = {1'b0,layer_2_1[4607:4600]} - {1'b0, layer_1_1[4607:4600]};
      mid_2[0] = {1'b0,layer_2_2[4591:4584]} - {1'b0, layer_1_2[4591:4584]};
      mid_2[1] = {1'b0,layer_2_2[4599:4592]} - {1'b0, layer_1_2[4599:4592]};
      mid_2[2] = {1'b0,layer_2_2[4607:4600]} - {1'b0, layer_1_2[4607:4600]};
      btm_0[0] = {1'b0,layer_3_0[4591:4584]} - {1'b0, layer_2_0[4591:4584]};
      btm_0[1] = {1'b0,layer_3_0[4599:4592]} - {1'b0, layer_2_0[4599:4592]};
      btm_0[2] = {1'b0,layer_3_0[4607:4600]} - {1'b0, layer_2_0[4607:4600]};
      btm_1[0] = {1'b0,layer_3_1[4591:4584]} - {1'b0, layer_2_1[4591:4584]};
      btm_1[1] = {1'b0,layer_3_1[4599:4592]} - {1'b0, layer_2_1[4599:4592]};
      btm_1[2] = {1'b0,layer_3_1[4607:4600]} - {1'b0, layer_2_1[4607:4600]};
      btm_2[0] = {1'b0,layer_3_2[4591:4584]} - {1'b0, layer_2_2[4591:4584]};
      btm_2[1] = {1'b0,layer_3_2[4599:4592]} - {1'b0, layer_2_2[4599:4592]};
      btm_2[2] = {1'b0,layer_3_2[4607:4600]} - {1'b0, layer_2_2[4607:4600]};
    end
    'd575: begin
      top_0[0] = {1'b0,layer_1_0[4599:4592]} - {1'b0, layer_0_0[4599:4592]};
      top_0[1] = {1'b0,layer_1_0[4607:4600]} - {1'b0, layer_0_0[4607:4600]};
      top_0[2] = {1'b0,layer_1_0[4615:4608]} - {1'b0, layer_0_0[4615:4608]};
      top_1[0] = {1'b0,layer_1_1[4599:4592]} - {1'b0, layer_0_1[4599:4592]};
      top_1[1] = {1'b0,layer_1_1[4607:4600]} - {1'b0, layer_0_1[4607:4600]};
      top_1[2] = {1'b0,layer_1_1[4615:4608]} - {1'b0, layer_0_1[4615:4608]};
      top_2[0] = {1'b0,layer_1_2[4599:4592]} - {1'b0, layer_0_2[4599:4592]};
      top_2[1] = {1'b0,layer_1_2[4607:4600]} - {1'b0, layer_0_2[4607:4600]};
      top_2[2] = {1'b0,layer_1_2[4615:4608]} - {1'b0, layer_0_2[4615:4608]};
      mid_0[0] = {1'b0,layer_2_0[4599:4592]} - {1'b0, layer_1_0[4599:4592]};
      mid_0[1] = {1'b0,layer_2_0[4607:4600]} - {1'b0, layer_1_0[4607:4600]};
      mid_0[2] = {1'b0,layer_2_0[4615:4608]} - {1'b0, layer_1_0[4615:4608]};
      mid_1[0] = {1'b0,layer_2_1[4599:4592]} - {1'b0, layer_1_1[4599:4592]};
      mid_1[1] = {1'b0,layer_2_1[4607:4600]} - {1'b0, layer_1_1[4607:4600]};
      mid_1[2] = {1'b0,layer_2_1[4615:4608]} - {1'b0, layer_1_1[4615:4608]};
      mid_2[0] = {1'b0,layer_2_2[4599:4592]} - {1'b0, layer_1_2[4599:4592]};
      mid_2[1] = {1'b0,layer_2_2[4607:4600]} - {1'b0, layer_1_2[4607:4600]};
      mid_2[2] = {1'b0,layer_2_2[4615:4608]} - {1'b0, layer_1_2[4615:4608]};
      btm_0[0] = {1'b0,layer_3_0[4599:4592]} - {1'b0, layer_2_0[4599:4592]};
      btm_0[1] = {1'b0,layer_3_0[4607:4600]} - {1'b0, layer_2_0[4607:4600]};
      btm_0[2] = {1'b0,layer_3_0[4615:4608]} - {1'b0, layer_2_0[4615:4608]};
      btm_1[0] = {1'b0,layer_3_1[4599:4592]} - {1'b0, layer_2_1[4599:4592]};
      btm_1[1] = {1'b0,layer_3_1[4607:4600]} - {1'b0, layer_2_1[4607:4600]};
      btm_1[2] = {1'b0,layer_3_1[4615:4608]} - {1'b0, layer_2_1[4615:4608]};
      btm_2[0] = {1'b0,layer_3_2[4599:4592]} - {1'b0, layer_2_2[4599:4592]};
      btm_2[1] = {1'b0,layer_3_2[4607:4600]} - {1'b0, layer_2_2[4607:4600]};
      btm_2[2] = {1'b0,layer_3_2[4615:4608]} - {1'b0, layer_2_2[4615:4608]};
    end
    'd576: begin
      top_0[0] = {1'b0,layer_1_0[4607:4600]} - {1'b0, layer_0_0[4607:4600]};
      top_0[1] = {1'b0,layer_1_0[4615:4608]} - {1'b0, layer_0_0[4615:4608]};
      top_0[2] = {1'b0,layer_1_0[4623:4616]} - {1'b0, layer_0_0[4623:4616]};
      top_1[0] = {1'b0,layer_1_1[4607:4600]} - {1'b0, layer_0_1[4607:4600]};
      top_1[1] = {1'b0,layer_1_1[4615:4608]} - {1'b0, layer_0_1[4615:4608]};
      top_1[2] = {1'b0,layer_1_1[4623:4616]} - {1'b0, layer_0_1[4623:4616]};
      top_2[0] = {1'b0,layer_1_2[4607:4600]} - {1'b0, layer_0_2[4607:4600]};
      top_2[1] = {1'b0,layer_1_2[4615:4608]} - {1'b0, layer_0_2[4615:4608]};
      top_2[2] = {1'b0,layer_1_2[4623:4616]} - {1'b0, layer_0_2[4623:4616]};
      mid_0[0] = {1'b0,layer_2_0[4607:4600]} - {1'b0, layer_1_0[4607:4600]};
      mid_0[1] = {1'b0,layer_2_0[4615:4608]} - {1'b0, layer_1_0[4615:4608]};
      mid_0[2] = {1'b0,layer_2_0[4623:4616]} - {1'b0, layer_1_0[4623:4616]};
      mid_1[0] = {1'b0,layer_2_1[4607:4600]} - {1'b0, layer_1_1[4607:4600]};
      mid_1[1] = {1'b0,layer_2_1[4615:4608]} - {1'b0, layer_1_1[4615:4608]};
      mid_1[2] = {1'b0,layer_2_1[4623:4616]} - {1'b0, layer_1_1[4623:4616]};
      mid_2[0] = {1'b0,layer_2_2[4607:4600]} - {1'b0, layer_1_2[4607:4600]};
      mid_2[1] = {1'b0,layer_2_2[4615:4608]} - {1'b0, layer_1_2[4615:4608]};
      mid_2[2] = {1'b0,layer_2_2[4623:4616]} - {1'b0, layer_1_2[4623:4616]};
      btm_0[0] = {1'b0,layer_3_0[4607:4600]} - {1'b0, layer_2_0[4607:4600]};
      btm_0[1] = {1'b0,layer_3_0[4615:4608]} - {1'b0, layer_2_0[4615:4608]};
      btm_0[2] = {1'b0,layer_3_0[4623:4616]} - {1'b0, layer_2_0[4623:4616]};
      btm_1[0] = {1'b0,layer_3_1[4607:4600]} - {1'b0, layer_2_1[4607:4600]};
      btm_1[1] = {1'b0,layer_3_1[4615:4608]} - {1'b0, layer_2_1[4615:4608]};
      btm_1[2] = {1'b0,layer_3_1[4623:4616]} - {1'b0, layer_2_1[4623:4616]};
      btm_2[0] = {1'b0,layer_3_2[4607:4600]} - {1'b0, layer_2_2[4607:4600]};
      btm_2[1] = {1'b0,layer_3_2[4615:4608]} - {1'b0, layer_2_2[4615:4608]};
      btm_2[2] = {1'b0,layer_3_2[4623:4616]} - {1'b0, layer_2_2[4623:4616]};
    end
    'd577: begin
      top_0[0] = {1'b0,layer_1_0[4615:4608]} - {1'b0, layer_0_0[4615:4608]};
      top_0[1] = {1'b0,layer_1_0[4623:4616]} - {1'b0, layer_0_0[4623:4616]};
      top_0[2] = {1'b0,layer_1_0[4631:4624]} - {1'b0, layer_0_0[4631:4624]};
      top_1[0] = {1'b0,layer_1_1[4615:4608]} - {1'b0, layer_0_1[4615:4608]};
      top_1[1] = {1'b0,layer_1_1[4623:4616]} - {1'b0, layer_0_1[4623:4616]};
      top_1[2] = {1'b0,layer_1_1[4631:4624]} - {1'b0, layer_0_1[4631:4624]};
      top_2[0] = {1'b0,layer_1_2[4615:4608]} - {1'b0, layer_0_2[4615:4608]};
      top_2[1] = {1'b0,layer_1_2[4623:4616]} - {1'b0, layer_0_2[4623:4616]};
      top_2[2] = {1'b0,layer_1_2[4631:4624]} - {1'b0, layer_0_2[4631:4624]};
      mid_0[0] = {1'b0,layer_2_0[4615:4608]} - {1'b0, layer_1_0[4615:4608]};
      mid_0[1] = {1'b0,layer_2_0[4623:4616]} - {1'b0, layer_1_0[4623:4616]};
      mid_0[2] = {1'b0,layer_2_0[4631:4624]} - {1'b0, layer_1_0[4631:4624]};
      mid_1[0] = {1'b0,layer_2_1[4615:4608]} - {1'b0, layer_1_1[4615:4608]};
      mid_1[1] = {1'b0,layer_2_1[4623:4616]} - {1'b0, layer_1_1[4623:4616]};
      mid_1[2] = {1'b0,layer_2_1[4631:4624]} - {1'b0, layer_1_1[4631:4624]};
      mid_2[0] = {1'b0,layer_2_2[4615:4608]} - {1'b0, layer_1_2[4615:4608]};
      mid_2[1] = {1'b0,layer_2_2[4623:4616]} - {1'b0, layer_1_2[4623:4616]};
      mid_2[2] = {1'b0,layer_2_2[4631:4624]} - {1'b0, layer_1_2[4631:4624]};
      btm_0[0] = {1'b0,layer_3_0[4615:4608]} - {1'b0, layer_2_0[4615:4608]};
      btm_0[1] = {1'b0,layer_3_0[4623:4616]} - {1'b0, layer_2_0[4623:4616]};
      btm_0[2] = {1'b0,layer_3_0[4631:4624]} - {1'b0, layer_2_0[4631:4624]};
      btm_1[0] = {1'b0,layer_3_1[4615:4608]} - {1'b0, layer_2_1[4615:4608]};
      btm_1[1] = {1'b0,layer_3_1[4623:4616]} - {1'b0, layer_2_1[4623:4616]};
      btm_1[2] = {1'b0,layer_3_1[4631:4624]} - {1'b0, layer_2_1[4631:4624]};
      btm_2[0] = {1'b0,layer_3_2[4615:4608]} - {1'b0, layer_2_2[4615:4608]};
      btm_2[1] = {1'b0,layer_3_2[4623:4616]} - {1'b0, layer_2_2[4623:4616]};
      btm_2[2] = {1'b0,layer_3_2[4631:4624]} - {1'b0, layer_2_2[4631:4624]};
    end
    'd578: begin
      top_0[0] = {1'b0,layer_1_0[4623:4616]} - {1'b0, layer_0_0[4623:4616]};
      top_0[1] = {1'b0,layer_1_0[4631:4624]} - {1'b0, layer_0_0[4631:4624]};
      top_0[2] = {1'b0,layer_1_0[4639:4632]} - {1'b0, layer_0_0[4639:4632]};
      top_1[0] = {1'b0,layer_1_1[4623:4616]} - {1'b0, layer_0_1[4623:4616]};
      top_1[1] = {1'b0,layer_1_1[4631:4624]} - {1'b0, layer_0_1[4631:4624]};
      top_1[2] = {1'b0,layer_1_1[4639:4632]} - {1'b0, layer_0_1[4639:4632]};
      top_2[0] = {1'b0,layer_1_2[4623:4616]} - {1'b0, layer_0_2[4623:4616]};
      top_2[1] = {1'b0,layer_1_2[4631:4624]} - {1'b0, layer_0_2[4631:4624]};
      top_2[2] = {1'b0,layer_1_2[4639:4632]} - {1'b0, layer_0_2[4639:4632]};
      mid_0[0] = {1'b0,layer_2_0[4623:4616]} - {1'b0, layer_1_0[4623:4616]};
      mid_0[1] = {1'b0,layer_2_0[4631:4624]} - {1'b0, layer_1_0[4631:4624]};
      mid_0[2] = {1'b0,layer_2_0[4639:4632]} - {1'b0, layer_1_0[4639:4632]};
      mid_1[0] = {1'b0,layer_2_1[4623:4616]} - {1'b0, layer_1_1[4623:4616]};
      mid_1[1] = {1'b0,layer_2_1[4631:4624]} - {1'b0, layer_1_1[4631:4624]};
      mid_1[2] = {1'b0,layer_2_1[4639:4632]} - {1'b0, layer_1_1[4639:4632]};
      mid_2[0] = {1'b0,layer_2_2[4623:4616]} - {1'b0, layer_1_2[4623:4616]};
      mid_2[1] = {1'b0,layer_2_2[4631:4624]} - {1'b0, layer_1_2[4631:4624]};
      mid_2[2] = {1'b0,layer_2_2[4639:4632]} - {1'b0, layer_1_2[4639:4632]};
      btm_0[0] = {1'b0,layer_3_0[4623:4616]} - {1'b0, layer_2_0[4623:4616]};
      btm_0[1] = {1'b0,layer_3_0[4631:4624]} - {1'b0, layer_2_0[4631:4624]};
      btm_0[2] = {1'b0,layer_3_0[4639:4632]} - {1'b0, layer_2_0[4639:4632]};
      btm_1[0] = {1'b0,layer_3_1[4623:4616]} - {1'b0, layer_2_1[4623:4616]};
      btm_1[1] = {1'b0,layer_3_1[4631:4624]} - {1'b0, layer_2_1[4631:4624]};
      btm_1[2] = {1'b0,layer_3_1[4639:4632]} - {1'b0, layer_2_1[4639:4632]};
      btm_2[0] = {1'b0,layer_3_2[4623:4616]} - {1'b0, layer_2_2[4623:4616]};
      btm_2[1] = {1'b0,layer_3_2[4631:4624]} - {1'b0, layer_2_2[4631:4624]};
      btm_2[2] = {1'b0,layer_3_2[4639:4632]} - {1'b0, layer_2_2[4639:4632]};
    end
    'd579: begin
      top_0[0] = {1'b0,layer_1_0[4631:4624]} - {1'b0, layer_0_0[4631:4624]};
      top_0[1] = {1'b0,layer_1_0[4639:4632]} - {1'b0, layer_0_0[4639:4632]};
      top_0[2] = {1'b0,layer_1_0[4647:4640]} - {1'b0, layer_0_0[4647:4640]};
      top_1[0] = {1'b0,layer_1_1[4631:4624]} - {1'b0, layer_0_1[4631:4624]};
      top_1[1] = {1'b0,layer_1_1[4639:4632]} - {1'b0, layer_0_1[4639:4632]};
      top_1[2] = {1'b0,layer_1_1[4647:4640]} - {1'b0, layer_0_1[4647:4640]};
      top_2[0] = {1'b0,layer_1_2[4631:4624]} - {1'b0, layer_0_2[4631:4624]};
      top_2[1] = {1'b0,layer_1_2[4639:4632]} - {1'b0, layer_0_2[4639:4632]};
      top_2[2] = {1'b0,layer_1_2[4647:4640]} - {1'b0, layer_0_2[4647:4640]};
      mid_0[0] = {1'b0,layer_2_0[4631:4624]} - {1'b0, layer_1_0[4631:4624]};
      mid_0[1] = {1'b0,layer_2_0[4639:4632]} - {1'b0, layer_1_0[4639:4632]};
      mid_0[2] = {1'b0,layer_2_0[4647:4640]} - {1'b0, layer_1_0[4647:4640]};
      mid_1[0] = {1'b0,layer_2_1[4631:4624]} - {1'b0, layer_1_1[4631:4624]};
      mid_1[1] = {1'b0,layer_2_1[4639:4632]} - {1'b0, layer_1_1[4639:4632]};
      mid_1[2] = {1'b0,layer_2_1[4647:4640]} - {1'b0, layer_1_1[4647:4640]};
      mid_2[0] = {1'b0,layer_2_2[4631:4624]} - {1'b0, layer_1_2[4631:4624]};
      mid_2[1] = {1'b0,layer_2_2[4639:4632]} - {1'b0, layer_1_2[4639:4632]};
      mid_2[2] = {1'b0,layer_2_2[4647:4640]} - {1'b0, layer_1_2[4647:4640]};
      btm_0[0] = {1'b0,layer_3_0[4631:4624]} - {1'b0, layer_2_0[4631:4624]};
      btm_0[1] = {1'b0,layer_3_0[4639:4632]} - {1'b0, layer_2_0[4639:4632]};
      btm_0[2] = {1'b0,layer_3_0[4647:4640]} - {1'b0, layer_2_0[4647:4640]};
      btm_1[0] = {1'b0,layer_3_1[4631:4624]} - {1'b0, layer_2_1[4631:4624]};
      btm_1[1] = {1'b0,layer_3_1[4639:4632]} - {1'b0, layer_2_1[4639:4632]};
      btm_1[2] = {1'b0,layer_3_1[4647:4640]} - {1'b0, layer_2_1[4647:4640]};
      btm_2[0] = {1'b0,layer_3_2[4631:4624]} - {1'b0, layer_2_2[4631:4624]};
      btm_2[1] = {1'b0,layer_3_2[4639:4632]} - {1'b0, layer_2_2[4639:4632]};
      btm_2[2] = {1'b0,layer_3_2[4647:4640]} - {1'b0, layer_2_2[4647:4640]};
    end
    'd580: begin
      top_0[0] = {1'b0,layer_1_0[4639:4632]} - {1'b0, layer_0_0[4639:4632]};
      top_0[1] = {1'b0,layer_1_0[4647:4640]} - {1'b0, layer_0_0[4647:4640]};
      top_0[2] = {1'b0,layer_1_0[4655:4648]} - {1'b0, layer_0_0[4655:4648]};
      top_1[0] = {1'b0,layer_1_1[4639:4632]} - {1'b0, layer_0_1[4639:4632]};
      top_1[1] = {1'b0,layer_1_1[4647:4640]} - {1'b0, layer_0_1[4647:4640]};
      top_1[2] = {1'b0,layer_1_1[4655:4648]} - {1'b0, layer_0_1[4655:4648]};
      top_2[0] = {1'b0,layer_1_2[4639:4632]} - {1'b0, layer_0_2[4639:4632]};
      top_2[1] = {1'b0,layer_1_2[4647:4640]} - {1'b0, layer_0_2[4647:4640]};
      top_2[2] = {1'b0,layer_1_2[4655:4648]} - {1'b0, layer_0_2[4655:4648]};
      mid_0[0] = {1'b0,layer_2_0[4639:4632]} - {1'b0, layer_1_0[4639:4632]};
      mid_0[1] = {1'b0,layer_2_0[4647:4640]} - {1'b0, layer_1_0[4647:4640]};
      mid_0[2] = {1'b0,layer_2_0[4655:4648]} - {1'b0, layer_1_0[4655:4648]};
      mid_1[0] = {1'b0,layer_2_1[4639:4632]} - {1'b0, layer_1_1[4639:4632]};
      mid_1[1] = {1'b0,layer_2_1[4647:4640]} - {1'b0, layer_1_1[4647:4640]};
      mid_1[2] = {1'b0,layer_2_1[4655:4648]} - {1'b0, layer_1_1[4655:4648]};
      mid_2[0] = {1'b0,layer_2_2[4639:4632]} - {1'b0, layer_1_2[4639:4632]};
      mid_2[1] = {1'b0,layer_2_2[4647:4640]} - {1'b0, layer_1_2[4647:4640]};
      mid_2[2] = {1'b0,layer_2_2[4655:4648]} - {1'b0, layer_1_2[4655:4648]};
      btm_0[0] = {1'b0,layer_3_0[4639:4632]} - {1'b0, layer_2_0[4639:4632]};
      btm_0[1] = {1'b0,layer_3_0[4647:4640]} - {1'b0, layer_2_0[4647:4640]};
      btm_0[2] = {1'b0,layer_3_0[4655:4648]} - {1'b0, layer_2_0[4655:4648]};
      btm_1[0] = {1'b0,layer_3_1[4639:4632]} - {1'b0, layer_2_1[4639:4632]};
      btm_1[1] = {1'b0,layer_3_1[4647:4640]} - {1'b0, layer_2_1[4647:4640]};
      btm_1[2] = {1'b0,layer_3_1[4655:4648]} - {1'b0, layer_2_1[4655:4648]};
      btm_2[0] = {1'b0,layer_3_2[4639:4632]} - {1'b0, layer_2_2[4639:4632]};
      btm_2[1] = {1'b0,layer_3_2[4647:4640]} - {1'b0, layer_2_2[4647:4640]};
      btm_2[2] = {1'b0,layer_3_2[4655:4648]} - {1'b0, layer_2_2[4655:4648]};
    end
    'd581: begin
      top_0[0] = {1'b0,layer_1_0[4647:4640]} - {1'b0, layer_0_0[4647:4640]};
      top_0[1] = {1'b0,layer_1_0[4655:4648]} - {1'b0, layer_0_0[4655:4648]};
      top_0[2] = {1'b0,layer_1_0[4663:4656]} - {1'b0, layer_0_0[4663:4656]};
      top_1[0] = {1'b0,layer_1_1[4647:4640]} - {1'b0, layer_0_1[4647:4640]};
      top_1[1] = {1'b0,layer_1_1[4655:4648]} - {1'b0, layer_0_1[4655:4648]};
      top_1[2] = {1'b0,layer_1_1[4663:4656]} - {1'b0, layer_0_1[4663:4656]};
      top_2[0] = {1'b0,layer_1_2[4647:4640]} - {1'b0, layer_0_2[4647:4640]};
      top_2[1] = {1'b0,layer_1_2[4655:4648]} - {1'b0, layer_0_2[4655:4648]};
      top_2[2] = {1'b0,layer_1_2[4663:4656]} - {1'b0, layer_0_2[4663:4656]};
      mid_0[0] = {1'b0,layer_2_0[4647:4640]} - {1'b0, layer_1_0[4647:4640]};
      mid_0[1] = {1'b0,layer_2_0[4655:4648]} - {1'b0, layer_1_0[4655:4648]};
      mid_0[2] = {1'b0,layer_2_0[4663:4656]} - {1'b0, layer_1_0[4663:4656]};
      mid_1[0] = {1'b0,layer_2_1[4647:4640]} - {1'b0, layer_1_1[4647:4640]};
      mid_1[1] = {1'b0,layer_2_1[4655:4648]} - {1'b0, layer_1_1[4655:4648]};
      mid_1[2] = {1'b0,layer_2_1[4663:4656]} - {1'b0, layer_1_1[4663:4656]};
      mid_2[0] = {1'b0,layer_2_2[4647:4640]} - {1'b0, layer_1_2[4647:4640]};
      mid_2[1] = {1'b0,layer_2_2[4655:4648]} - {1'b0, layer_1_2[4655:4648]};
      mid_2[2] = {1'b0,layer_2_2[4663:4656]} - {1'b0, layer_1_2[4663:4656]};
      btm_0[0] = {1'b0,layer_3_0[4647:4640]} - {1'b0, layer_2_0[4647:4640]};
      btm_0[1] = {1'b0,layer_3_0[4655:4648]} - {1'b0, layer_2_0[4655:4648]};
      btm_0[2] = {1'b0,layer_3_0[4663:4656]} - {1'b0, layer_2_0[4663:4656]};
      btm_1[0] = {1'b0,layer_3_1[4647:4640]} - {1'b0, layer_2_1[4647:4640]};
      btm_1[1] = {1'b0,layer_3_1[4655:4648]} - {1'b0, layer_2_1[4655:4648]};
      btm_1[2] = {1'b0,layer_3_1[4663:4656]} - {1'b0, layer_2_1[4663:4656]};
      btm_2[0] = {1'b0,layer_3_2[4647:4640]} - {1'b0, layer_2_2[4647:4640]};
      btm_2[1] = {1'b0,layer_3_2[4655:4648]} - {1'b0, layer_2_2[4655:4648]};
      btm_2[2] = {1'b0,layer_3_2[4663:4656]} - {1'b0, layer_2_2[4663:4656]};
    end
    'd582: begin
      top_0[0] = {1'b0,layer_1_0[4655:4648]} - {1'b0, layer_0_0[4655:4648]};
      top_0[1] = {1'b0,layer_1_0[4663:4656]} - {1'b0, layer_0_0[4663:4656]};
      top_0[2] = {1'b0,layer_1_0[4671:4664]} - {1'b0, layer_0_0[4671:4664]};
      top_1[0] = {1'b0,layer_1_1[4655:4648]} - {1'b0, layer_0_1[4655:4648]};
      top_1[1] = {1'b0,layer_1_1[4663:4656]} - {1'b0, layer_0_1[4663:4656]};
      top_1[2] = {1'b0,layer_1_1[4671:4664]} - {1'b0, layer_0_1[4671:4664]};
      top_2[0] = {1'b0,layer_1_2[4655:4648]} - {1'b0, layer_0_2[4655:4648]};
      top_2[1] = {1'b0,layer_1_2[4663:4656]} - {1'b0, layer_0_2[4663:4656]};
      top_2[2] = {1'b0,layer_1_2[4671:4664]} - {1'b0, layer_0_2[4671:4664]};
      mid_0[0] = {1'b0,layer_2_0[4655:4648]} - {1'b0, layer_1_0[4655:4648]};
      mid_0[1] = {1'b0,layer_2_0[4663:4656]} - {1'b0, layer_1_0[4663:4656]};
      mid_0[2] = {1'b0,layer_2_0[4671:4664]} - {1'b0, layer_1_0[4671:4664]};
      mid_1[0] = {1'b0,layer_2_1[4655:4648]} - {1'b0, layer_1_1[4655:4648]};
      mid_1[1] = {1'b0,layer_2_1[4663:4656]} - {1'b0, layer_1_1[4663:4656]};
      mid_1[2] = {1'b0,layer_2_1[4671:4664]} - {1'b0, layer_1_1[4671:4664]};
      mid_2[0] = {1'b0,layer_2_2[4655:4648]} - {1'b0, layer_1_2[4655:4648]};
      mid_2[1] = {1'b0,layer_2_2[4663:4656]} - {1'b0, layer_1_2[4663:4656]};
      mid_2[2] = {1'b0,layer_2_2[4671:4664]} - {1'b0, layer_1_2[4671:4664]};
      btm_0[0] = {1'b0,layer_3_0[4655:4648]} - {1'b0, layer_2_0[4655:4648]};
      btm_0[1] = {1'b0,layer_3_0[4663:4656]} - {1'b0, layer_2_0[4663:4656]};
      btm_0[2] = {1'b0,layer_3_0[4671:4664]} - {1'b0, layer_2_0[4671:4664]};
      btm_1[0] = {1'b0,layer_3_1[4655:4648]} - {1'b0, layer_2_1[4655:4648]};
      btm_1[1] = {1'b0,layer_3_1[4663:4656]} - {1'b0, layer_2_1[4663:4656]};
      btm_1[2] = {1'b0,layer_3_1[4671:4664]} - {1'b0, layer_2_1[4671:4664]};
      btm_2[0] = {1'b0,layer_3_2[4655:4648]} - {1'b0, layer_2_2[4655:4648]};
      btm_2[1] = {1'b0,layer_3_2[4663:4656]} - {1'b0, layer_2_2[4663:4656]};
      btm_2[2] = {1'b0,layer_3_2[4671:4664]} - {1'b0, layer_2_2[4671:4664]};
    end
    'd583: begin
      top_0[0] = {1'b0,layer_1_0[4663:4656]} - {1'b0, layer_0_0[4663:4656]};
      top_0[1] = {1'b0,layer_1_0[4671:4664]} - {1'b0, layer_0_0[4671:4664]};
      top_0[2] = {1'b0,layer_1_0[4679:4672]} - {1'b0, layer_0_0[4679:4672]};
      top_1[0] = {1'b0,layer_1_1[4663:4656]} - {1'b0, layer_0_1[4663:4656]};
      top_1[1] = {1'b0,layer_1_1[4671:4664]} - {1'b0, layer_0_1[4671:4664]};
      top_1[2] = {1'b0,layer_1_1[4679:4672]} - {1'b0, layer_0_1[4679:4672]};
      top_2[0] = {1'b0,layer_1_2[4663:4656]} - {1'b0, layer_0_2[4663:4656]};
      top_2[1] = {1'b0,layer_1_2[4671:4664]} - {1'b0, layer_0_2[4671:4664]};
      top_2[2] = {1'b0,layer_1_2[4679:4672]} - {1'b0, layer_0_2[4679:4672]};
      mid_0[0] = {1'b0,layer_2_0[4663:4656]} - {1'b0, layer_1_0[4663:4656]};
      mid_0[1] = {1'b0,layer_2_0[4671:4664]} - {1'b0, layer_1_0[4671:4664]};
      mid_0[2] = {1'b0,layer_2_0[4679:4672]} - {1'b0, layer_1_0[4679:4672]};
      mid_1[0] = {1'b0,layer_2_1[4663:4656]} - {1'b0, layer_1_1[4663:4656]};
      mid_1[1] = {1'b0,layer_2_1[4671:4664]} - {1'b0, layer_1_1[4671:4664]};
      mid_1[2] = {1'b0,layer_2_1[4679:4672]} - {1'b0, layer_1_1[4679:4672]};
      mid_2[0] = {1'b0,layer_2_2[4663:4656]} - {1'b0, layer_1_2[4663:4656]};
      mid_2[1] = {1'b0,layer_2_2[4671:4664]} - {1'b0, layer_1_2[4671:4664]};
      mid_2[2] = {1'b0,layer_2_2[4679:4672]} - {1'b0, layer_1_2[4679:4672]};
      btm_0[0] = {1'b0,layer_3_0[4663:4656]} - {1'b0, layer_2_0[4663:4656]};
      btm_0[1] = {1'b0,layer_3_0[4671:4664]} - {1'b0, layer_2_0[4671:4664]};
      btm_0[2] = {1'b0,layer_3_0[4679:4672]} - {1'b0, layer_2_0[4679:4672]};
      btm_1[0] = {1'b0,layer_3_1[4663:4656]} - {1'b0, layer_2_1[4663:4656]};
      btm_1[1] = {1'b0,layer_3_1[4671:4664]} - {1'b0, layer_2_1[4671:4664]};
      btm_1[2] = {1'b0,layer_3_1[4679:4672]} - {1'b0, layer_2_1[4679:4672]};
      btm_2[0] = {1'b0,layer_3_2[4663:4656]} - {1'b0, layer_2_2[4663:4656]};
      btm_2[1] = {1'b0,layer_3_2[4671:4664]} - {1'b0, layer_2_2[4671:4664]};
      btm_2[2] = {1'b0,layer_3_2[4679:4672]} - {1'b0, layer_2_2[4679:4672]};
    end
    'd584: begin
      top_0[0] = {1'b0,layer_1_0[4671:4664]} - {1'b0, layer_0_0[4671:4664]};
      top_0[1] = {1'b0,layer_1_0[4679:4672]} - {1'b0, layer_0_0[4679:4672]};
      top_0[2] = {1'b0,layer_1_0[4687:4680]} - {1'b0, layer_0_0[4687:4680]};
      top_1[0] = {1'b0,layer_1_1[4671:4664]} - {1'b0, layer_0_1[4671:4664]};
      top_1[1] = {1'b0,layer_1_1[4679:4672]} - {1'b0, layer_0_1[4679:4672]};
      top_1[2] = {1'b0,layer_1_1[4687:4680]} - {1'b0, layer_0_1[4687:4680]};
      top_2[0] = {1'b0,layer_1_2[4671:4664]} - {1'b0, layer_0_2[4671:4664]};
      top_2[1] = {1'b0,layer_1_2[4679:4672]} - {1'b0, layer_0_2[4679:4672]};
      top_2[2] = {1'b0,layer_1_2[4687:4680]} - {1'b0, layer_0_2[4687:4680]};
      mid_0[0] = {1'b0,layer_2_0[4671:4664]} - {1'b0, layer_1_0[4671:4664]};
      mid_0[1] = {1'b0,layer_2_0[4679:4672]} - {1'b0, layer_1_0[4679:4672]};
      mid_0[2] = {1'b0,layer_2_0[4687:4680]} - {1'b0, layer_1_0[4687:4680]};
      mid_1[0] = {1'b0,layer_2_1[4671:4664]} - {1'b0, layer_1_1[4671:4664]};
      mid_1[1] = {1'b0,layer_2_1[4679:4672]} - {1'b0, layer_1_1[4679:4672]};
      mid_1[2] = {1'b0,layer_2_1[4687:4680]} - {1'b0, layer_1_1[4687:4680]};
      mid_2[0] = {1'b0,layer_2_2[4671:4664]} - {1'b0, layer_1_2[4671:4664]};
      mid_2[1] = {1'b0,layer_2_2[4679:4672]} - {1'b0, layer_1_2[4679:4672]};
      mid_2[2] = {1'b0,layer_2_2[4687:4680]} - {1'b0, layer_1_2[4687:4680]};
      btm_0[0] = {1'b0,layer_3_0[4671:4664]} - {1'b0, layer_2_0[4671:4664]};
      btm_0[1] = {1'b0,layer_3_0[4679:4672]} - {1'b0, layer_2_0[4679:4672]};
      btm_0[2] = {1'b0,layer_3_0[4687:4680]} - {1'b0, layer_2_0[4687:4680]};
      btm_1[0] = {1'b0,layer_3_1[4671:4664]} - {1'b0, layer_2_1[4671:4664]};
      btm_1[1] = {1'b0,layer_3_1[4679:4672]} - {1'b0, layer_2_1[4679:4672]};
      btm_1[2] = {1'b0,layer_3_1[4687:4680]} - {1'b0, layer_2_1[4687:4680]};
      btm_2[0] = {1'b0,layer_3_2[4671:4664]} - {1'b0, layer_2_2[4671:4664]};
      btm_2[1] = {1'b0,layer_3_2[4679:4672]} - {1'b0, layer_2_2[4679:4672]};
      btm_2[2] = {1'b0,layer_3_2[4687:4680]} - {1'b0, layer_2_2[4687:4680]};
    end
    'd585: begin
      top_0[0] = {1'b0,layer_1_0[4679:4672]} - {1'b0, layer_0_0[4679:4672]};
      top_0[1] = {1'b0,layer_1_0[4687:4680]} - {1'b0, layer_0_0[4687:4680]};
      top_0[2] = {1'b0,layer_1_0[4695:4688]} - {1'b0, layer_0_0[4695:4688]};
      top_1[0] = {1'b0,layer_1_1[4679:4672]} - {1'b0, layer_0_1[4679:4672]};
      top_1[1] = {1'b0,layer_1_1[4687:4680]} - {1'b0, layer_0_1[4687:4680]};
      top_1[2] = {1'b0,layer_1_1[4695:4688]} - {1'b0, layer_0_1[4695:4688]};
      top_2[0] = {1'b0,layer_1_2[4679:4672]} - {1'b0, layer_0_2[4679:4672]};
      top_2[1] = {1'b0,layer_1_2[4687:4680]} - {1'b0, layer_0_2[4687:4680]};
      top_2[2] = {1'b0,layer_1_2[4695:4688]} - {1'b0, layer_0_2[4695:4688]};
      mid_0[0] = {1'b0,layer_2_0[4679:4672]} - {1'b0, layer_1_0[4679:4672]};
      mid_0[1] = {1'b0,layer_2_0[4687:4680]} - {1'b0, layer_1_0[4687:4680]};
      mid_0[2] = {1'b0,layer_2_0[4695:4688]} - {1'b0, layer_1_0[4695:4688]};
      mid_1[0] = {1'b0,layer_2_1[4679:4672]} - {1'b0, layer_1_1[4679:4672]};
      mid_1[1] = {1'b0,layer_2_1[4687:4680]} - {1'b0, layer_1_1[4687:4680]};
      mid_1[2] = {1'b0,layer_2_1[4695:4688]} - {1'b0, layer_1_1[4695:4688]};
      mid_2[0] = {1'b0,layer_2_2[4679:4672]} - {1'b0, layer_1_2[4679:4672]};
      mid_2[1] = {1'b0,layer_2_2[4687:4680]} - {1'b0, layer_1_2[4687:4680]};
      mid_2[2] = {1'b0,layer_2_2[4695:4688]} - {1'b0, layer_1_2[4695:4688]};
      btm_0[0] = {1'b0,layer_3_0[4679:4672]} - {1'b0, layer_2_0[4679:4672]};
      btm_0[1] = {1'b0,layer_3_0[4687:4680]} - {1'b0, layer_2_0[4687:4680]};
      btm_0[2] = {1'b0,layer_3_0[4695:4688]} - {1'b0, layer_2_0[4695:4688]};
      btm_1[0] = {1'b0,layer_3_1[4679:4672]} - {1'b0, layer_2_1[4679:4672]};
      btm_1[1] = {1'b0,layer_3_1[4687:4680]} - {1'b0, layer_2_1[4687:4680]};
      btm_1[2] = {1'b0,layer_3_1[4695:4688]} - {1'b0, layer_2_1[4695:4688]};
      btm_2[0] = {1'b0,layer_3_2[4679:4672]} - {1'b0, layer_2_2[4679:4672]};
      btm_2[1] = {1'b0,layer_3_2[4687:4680]} - {1'b0, layer_2_2[4687:4680]};
      btm_2[2] = {1'b0,layer_3_2[4695:4688]} - {1'b0, layer_2_2[4695:4688]};
    end
    'd586: begin
      top_0[0] = {1'b0,layer_1_0[4687:4680]} - {1'b0, layer_0_0[4687:4680]};
      top_0[1] = {1'b0,layer_1_0[4695:4688]} - {1'b0, layer_0_0[4695:4688]};
      top_0[2] = {1'b0,layer_1_0[4703:4696]} - {1'b0, layer_0_0[4703:4696]};
      top_1[0] = {1'b0,layer_1_1[4687:4680]} - {1'b0, layer_0_1[4687:4680]};
      top_1[1] = {1'b0,layer_1_1[4695:4688]} - {1'b0, layer_0_1[4695:4688]};
      top_1[2] = {1'b0,layer_1_1[4703:4696]} - {1'b0, layer_0_1[4703:4696]};
      top_2[0] = {1'b0,layer_1_2[4687:4680]} - {1'b0, layer_0_2[4687:4680]};
      top_2[1] = {1'b0,layer_1_2[4695:4688]} - {1'b0, layer_0_2[4695:4688]};
      top_2[2] = {1'b0,layer_1_2[4703:4696]} - {1'b0, layer_0_2[4703:4696]};
      mid_0[0] = {1'b0,layer_2_0[4687:4680]} - {1'b0, layer_1_0[4687:4680]};
      mid_0[1] = {1'b0,layer_2_0[4695:4688]} - {1'b0, layer_1_0[4695:4688]};
      mid_0[2] = {1'b0,layer_2_0[4703:4696]} - {1'b0, layer_1_0[4703:4696]};
      mid_1[0] = {1'b0,layer_2_1[4687:4680]} - {1'b0, layer_1_1[4687:4680]};
      mid_1[1] = {1'b0,layer_2_1[4695:4688]} - {1'b0, layer_1_1[4695:4688]};
      mid_1[2] = {1'b0,layer_2_1[4703:4696]} - {1'b0, layer_1_1[4703:4696]};
      mid_2[0] = {1'b0,layer_2_2[4687:4680]} - {1'b0, layer_1_2[4687:4680]};
      mid_2[1] = {1'b0,layer_2_2[4695:4688]} - {1'b0, layer_1_2[4695:4688]};
      mid_2[2] = {1'b0,layer_2_2[4703:4696]} - {1'b0, layer_1_2[4703:4696]};
      btm_0[0] = {1'b0,layer_3_0[4687:4680]} - {1'b0, layer_2_0[4687:4680]};
      btm_0[1] = {1'b0,layer_3_0[4695:4688]} - {1'b0, layer_2_0[4695:4688]};
      btm_0[2] = {1'b0,layer_3_0[4703:4696]} - {1'b0, layer_2_0[4703:4696]};
      btm_1[0] = {1'b0,layer_3_1[4687:4680]} - {1'b0, layer_2_1[4687:4680]};
      btm_1[1] = {1'b0,layer_3_1[4695:4688]} - {1'b0, layer_2_1[4695:4688]};
      btm_1[2] = {1'b0,layer_3_1[4703:4696]} - {1'b0, layer_2_1[4703:4696]};
      btm_2[0] = {1'b0,layer_3_2[4687:4680]} - {1'b0, layer_2_2[4687:4680]};
      btm_2[1] = {1'b0,layer_3_2[4695:4688]} - {1'b0, layer_2_2[4695:4688]};
      btm_2[2] = {1'b0,layer_3_2[4703:4696]} - {1'b0, layer_2_2[4703:4696]};
    end
    'd587: begin
      top_0[0] = {1'b0,layer_1_0[4695:4688]} - {1'b0, layer_0_0[4695:4688]};
      top_0[1] = {1'b0,layer_1_0[4703:4696]} - {1'b0, layer_0_0[4703:4696]};
      top_0[2] = {1'b0,layer_1_0[4711:4704]} - {1'b0, layer_0_0[4711:4704]};
      top_1[0] = {1'b0,layer_1_1[4695:4688]} - {1'b0, layer_0_1[4695:4688]};
      top_1[1] = {1'b0,layer_1_1[4703:4696]} - {1'b0, layer_0_1[4703:4696]};
      top_1[2] = {1'b0,layer_1_1[4711:4704]} - {1'b0, layer_0_1[4711:4704]};
      top_2[0] = {1'b0,layer_1_2[4695:4688]} - {1'b0, layer_0_2[4695:4688]};
      top_2[1] = {1'b0,layer_1_2[4703:4696]} - {1'b0, layer_0_2[4703:4696]};
      top_2[2] = {1'b0,layer_1_2[4711:4704]} - {1'b0, layer_0_2[4711:4704]};
      mid_0[0] = {1'b0,layer_2_0[4695:4688]} - {1'b0, layer_1_0[4695:4688]};
      mid_0[1] = {1'b0,layer_2_0[4703:4696]} - {1'b0, layer_1_0[4703:4696]};
      mid_0[2] = {1'b0,layer_2_0[4711:4704]} - {1'b0, layer_1_0[4711:4704]};
      mid_1[0] = {1'b0,layer_2_1[4695:4688]} - {1'b0, layer_1_1[4695:4688]};
      mid_1[1] = {1'b0,layer_2_1[4703:4696]} - {1'b0, layer_1_1[4703:4696]};
      mid_1[2] = {1'b0,layer_2_1[4711:4704]} - {1'b0, layer_1_1[4711:4704]};
      mid_2[0] = {1'b0,layer_2_2[4695:4688]} - {1'b0, layer_1_2[4695:4688]};
      mid_2[1] = {1'b0,layer_2_2[4703:4696]} - {1'b0, layer_1_2[4703:4696]};
      mid_2[2] = {1'b0,layer_2_2[4711:4704]} - {1'b0, layer_1_2[4711:4704]};
      btm_0[0] = {1'b0,layer_3_0[4695:4688]} - {1'b0, layer_2_0[4695:4688]};
      btm_0[1] = {1'b0,layer_3_0[4703:4696]} - {1'b0, layer_2_0[4703:4696]};
      btm_0[2] = {1'b0,layer_3_0[4711:4704]} - {1'b0, layer_2_0[4711:4704]};
      btm_1[0] = {1'b0,layer_3_1[4695:4688]} - {1'b0, layer_2_1[4695:4688]};
      btm_1[1] = {1'b0,layer_3_1[4703:4696]} - {1'b0, layer_2_1[4703:4696]};
      btm_1[2] = {1'b0,layer_3_1[4711:4704]} - {1'b0, layer_2_1[4711:4704]};
      btm_2[0] = {1'b0,layer_3_2[4695:4688]} - {1'b0, layer_2_2[4695:4688]};
      btm_2[1] = {1'b0,layer_3_2[4703:4696]} - {1'b0, layer_2_2[4703:4696]};
      btm_2[2] = {1'b0,layer_3_2[4711:4704]} - {1'b0, layer_2_2[4711:4704]};
    end
    'd588: begin
      top_0[0] = {1'b0,layer_1_0[4703:4696]} - {1'b0, layer_0_0[4703:4696]};
      top_0[1] = {1'b0,layer_1_0[4711:4704]} - {1'b0, layer_0_0[4711:4704]};
      top_0[2] = {1'b0,layer_1_0[4719:4712]} - {1'b0, layer_0_0[4719:4712]};
      top_1[0] = {1'b0,layer_1_1[4703:4696]} - {1'b0, layer_0_1[4703:4696]};
      top_1[1] = {1'b0,layer_1_1[4711:4704]} - {1'b0, layer_0_1[4711:4704]};
      top_1[2] = {1'b0,layer_1_1[4719:4712]} - {1'b0, layer_0_1[4719:4712]};
      top_2[0] = {1'b0,layer_1_2[4703:4696]} - {1'b0, layer_0_2[4703:4696]};
      top_2[1] = {1'b0,layer_1_2[4711:4704]} - {1'b0, layer_0_2[4711:4704]};
      top_2[2] = {1'b0,layer_1_2[4719:4712]} - {1'b0, layer_0_2[4719:4712]};
      mid_0[0] = {1'b0,layer_2_0[4703:4696]} - {1'b0, layer_1_0[4703:4696]};
      mid_0[1] = {1'b0,layer_2_0[4711:4704]} - {1'b0, layer_1_0[4711:4704]};
      mid_0[2] = {1'b0,layer_2_0[4719:4712]} - {1'b0, layer_1_0[4719:4712]};
      mid_1[0] = {1'b0,layer_2_1[4703:4696]} - {1'b0, layer_1_1[4703:4696]};
      mid_1[1] = {1'b0,layer_2_1[4711:4704]} - {1'b0, layer_1_1[4711:4704]};
      mid_1[2] = {1'b0,layer_2_1[4719:4712]} - {1'b0, layer_1_1[4719:4712]};
      mid_2[0] = {1'b0,layer_2_2[4703:4696]} - {1'b0, layer_1_2[4703:4696]};
      mid_2[1] = {1'b0,layer_2_2[4711:4704]} - {1'b0, layer_1_2[4711:4704]};
      mid_2[2] = {1'b0,layer_2_2[4719:4712]} - {1'b0, layer_1_2[4719:4712]};
      btm_0[0] = {1'b0,layer_3_0[4703:4696]} - {1'b0, layer_2_0[4703:4696]};
      btm_0[1] = {1'b0,layer_3_0[4711:4704]} - {1'b0, layer_2_0[4711:4704]};
      btm_0[2] = {1'b0,layer_3_0[4719:4712]} - {1'b0, layer_2_0[4719:4712]};
      btm_1[0] = {1'b0,layer_3_1[4703:4696]} - {1'b0, layer_2_1[4703:4696]};
      btm_1[1] = {1'b0,layer_3_1[4711:4704]} - {1'b0, layer_2_1[4711:4704]};
      btm_1[2] = {1'b0,layer_3_1[4719:4712]} - {1'b0, layer_2_1[4719:4712]};
      btm_2[0] = {1'b0,layer_3_2[4703:4696]} - {1'b0, layer_2_2[4703:4696]};
      btm_2[1] = {1'b0,layer_3_2[4711:4704]} - {1'b0, layer_2_2[4711:4704]};
      btm_2[2] = {1'b0,layer_3_2[4719:4712]} - {1'b0, layer_2_2[4719:4712]};
    end
    'd589: begin
      top_0[0] = {1'b0,layer_1_0[4711:4704]} - {1'b0, layer_0_0[4711:4704]};
      top_0[1] = {1'b0,layer_1_0[4719:4712]} - {1'b0, layer_0_0[4719:4712]};
      top_0[2] = {1'b0,layer_1_0[4727:4720]} - {1'b0, layer_0_0[4727:4720]};
      top_1[0] = {1'b0,layer_1_1[4711:4704]} - {1'b0, layer_0_1[4711:4704]};
      top_1[1] = {1'b0,layer_1_1[4719:4712]} - {1'b0, layer_0_1[4719:4712]};
      top_1[2] = {1'b0,layer_1_1[4727:4720]} - {1'b0, layer_0_1[4727:4720]};
      top_2[0] = {1'b0,layer_1_2[4711:4704]} - {1'b0, layer_0_2[4711:4704]};
      top_2[1] = {1'b0,layer_1_2[4719:4712]} - {1'b0, layer_0_2[4719:4712]};
      top_2[2] = {1'b0,layer_1_2[4727:4720]} - {1'b0, layer_0_2[4727:4720]};
      mid_0[0] = {1'b0,layer_2_0[4711:4704]} - {1'b0, layer_1_0[4711:4704]};
      mid_0[1] = {1'b0,layer_2_0[4719:4712]} - {1'b0, layer_1_0[4719:4712]};
      mid_0[2] = {1'b0,layer_2_0[4727:4720]} - {1'b0, layer_1_0[4727:4720]};
      mid_1[0] = {1'b0,layer_2_1[4711:4704]} - {1'b0, layer_1_1[4711:4704]};
      mid_1[1] = {1'b0,layer_2_1[4719:4712]} - {1'b0, layer_1_1[4719:4712]};
      mid_1[2] = {1'b0,layer_2_1[4727:4720]} - {1'b0, layer_1_1[4727:4720]};
      mid_2[0] = {1'b0,layer_2_2[4711:4704]} - {1'b0, layer_1_2[4711:4704]};
      mid_2[1] = {1'b0,layer_2_2[4719:4712]} - {1'b0, layer_1_2[4719:4712]};
      mid_2[2] = {1'b0,layer_2_2[4727:4720]} - {1'b0, layer_1_2[4727:4720]};
      btm_0[0] = {1'b0,layer_3_0[4711:4704]} - {1'b0, layer_2_0[4711:4704]};
      btm_0[1] = {1'b0,layer_3_0[4719:4712]} - {1'b0, layer_2_0[4719:4712]};
      btm_0[2] = {1'b0,layer_3_0[4727:4720]} - {1'b0, layer_2_0[4727:4720]};
      btm_1[0] = {1'b0,layer_3_1[4711:4704]} - {1'b0, layer_2_1[4711:4704]};
      btm_1[1] = {1'b0,layer_3_1[4719:4712]} - {1'b0, layer_2_1[4719:4712]};
      btm_1[2] = {1'b0,layer_3_1[4727:4720]} - {1'b0, layer_2_1[4727:4720]};
      btm_2[0] = {1'b0,layer_3_2[4711:4704]} - {1'b0, layer_2_2[4711:4704]};
      btm_2[1] = {1'b0,layer_3_2[4719:4712]} - {1'b0, layer_2_2[4719:4712]};
      btm_2[2] = {1'b0,layer_3_2[4727:4720]} - {1'b0, layer_2_2[4727:4720]};
    end
    'd590: begin
      top_0[0] = {1'b0,layer_1_0[4719:4712]} - {1'b0, layer_0_0[4719:4712]};
      top_0[1] = {1'b0,layer_1_0[4727:4720]} - {1'b0, layer_0_0[4727:4720]};
      top_0[2] = {1'b0,layer_1_0[4735:4728]} - {1'b0, layer_0_0[4735:4728]};
      top_1[0] = {1'b0,layer_1_1[4719:4712]} - {1'b0, layer_0_1[4719:4712]};
      top_1[1] = {1'b0,layer_1_1[4727:4720]} - {1'b0, layer_0_1[4727:4720]};
      top_1[2] = {1'b0,layer_1_1[4735:4728]} - {1'b0, layer_0_1[4735:4728]};
      top_2[0] = {1'b0,layer_1_2[4719:4712]} - {1'b0, layer_0_2[4719:4712]};
      top_2[1] = {1'b0,layer_1_2[4727:4720]} - {1'b0, layer_0_2[4727:4720]};
      top_2[2] = {1'b0,layer_1_2[4735:4728]} - {1'b0, layer_0_2[4735:4728]};
      mid_0[0] = {1'b0,layer_2_0[4719:4712]} - {1'b0, layer_1_0[4719:4712]};
      mid_0[1] = {1'b0,layer_2_0[4727:4720]} - {1'b0, layer_1_0[4727:4720]};
      mid_0[2] = {1'b0,layer_2_0[4735:4728]} - {1'b0, layer_1_0[4735:4728]};
      mid_1[0] = {1'b0,layer_2_1[4719:4712]} - {1'b0, layer_1_1[4719:4712]};
      mid_1[1] = {1'b0,layer_2_1[4727:4720]} - {1'b0, layer_1_1[4727:4720]};
      mid_1[2] = {1'b0,layer_2_1[4735:4728]} - {1'b0, layer_1_1[4735:4728]};
      mid_2[0] = {1'b0,layer_2_2[4719:4712]} - {1'b0, layer_1_2[4719:4712]};
      mid_2[1] = {1'b0,layer_2_2[4727:4720]} - {1'b0, layer_1_2[4727:4720]};
      mid_2[2] = {1'b0,layer_2_2[4735:4728]} - {1'b0, layer_1_2[4735:4728]};
      btm_0[0] = {1'b0,layer_3_0[4719:4712]} - {1'b0, layer_2_0[4719:4712]};
      btm_0[1] = {1'b0,layer_3_0[4727:4720]} - {1'b0, layer_2_0[4727:4720]};
      btm_0[2] = {1'b0,layer_3_0[4735:4728]} - {1'b0, layer_2_0[4735:4728]};
      btm_1[0] = {1'b0,layer_3_1[4719:4712]} - {1'b0, layer_2_1[4719:4712]};
      btm_1[1] = {1'b0,layer_3_1[4727:4720]} - {1'b0, layer_2_1[4727:4720]};
      btm_1[2] = {1'b0,layer_3_1[4735:4728]} - {1'b0, layer_2_1[4735:4728]};
      btm_2[0] = {1'b0,layer_3_2[4719:4712]} - {1'b0, layer_2_2[4719:4712]};
      btm_2[1] = {1'b0,layer_3_2[4727:4720]} - {1'b0, layer_2_2[4727:4720]};
      btm_2[2] = {1'b0,layer_3_2[4735:4728]} - {1'b0, layer_2_2[4735:4728]};
    end
    'd591: begin
      top_0[0] = {1'b0,layer_1_0[4727:4720]} - {1'b0, layer_0_0[4727:4720]};
      top_0[1] = {1'b0,layer_1_0[4735:4728]} - {1'b0, layer_0_0[4735:4728]};
      top_0[2] = {1'b0,layer_1_0[4743:4736]} - {1'b0, layer_0_0[4743:4736]};
      top_1[0] = {1'b0,layer_1_1[4727:4720]} - {1'b0, layer_0_1[4727:4720]};
      top_1[1] = {1'b0,layer_1_1[4735:4728]} - {1'b0, layer_0_1[4735:4728]};
      top_1[2] = {1'b0,layer_1_1[4743:4736]} - {1'b0, layer_0_1[4743:4736]};
      top_2[0] = {1'b0,layer_1_2[4727:4720]} - {1'b0, layer_0_2[4727:4720]};
      top_2[1] = {1'b0,layer_1_2[4735:4728]} - {1'b0, layer_0_2[4735:4728]};
      top_2[2] = {1'b0,layer_1_2[4743:4736]} - {1'b0, layer_0_2[4743:4736]};
      mid_0[0] = {1'b0,layer_2_0[4727:4720]} - {1'b0, layer_1_0[4727:4720]};
      mid_0[1] = {1'b0,layer_2_0[4735:4728]} - {1'b0, layer_1_0[4735:4728]};
      mid_0[2] = {1'b0,layer_2_0[4743:4736]} - {1'b0, layer_1_0[4743:4736]};
      mid_1[0] = {1'b0,layer_2_1[4727:4720]} - {1'b0, layer_1_1[4727:4720]};
      mid_1[1] = {1'b0,layer_2_1[4735:4728]} - {1'b0, layer_1_1[4735:4728]};
      mid_1[2] = {1'b0,layer_2_1[4743:4736]} - {1'b0, layer_1_1[4743:4736]};
      mid_2[0] = {1'b0,layer_2_2[4727:4720]} - {1'b0, layer_1_2[4727:4720]};
      mid_2[1] = {1'b0,layer_2_2[4735:4728]} - {1'b0, layer_1_2[4735:4728]};
      mid_2[2] = {1'b0,layer_2_2[4743:4736]} - {1'b0, layer_1_2[4743:4736]};
      btm_0[0] = {1'b0,layer_3_0[4727:4720]} - {1'b0, layer_2_0[4727:4720]};
      btm_0[1] = {1'b0,layer_3_0[4735:4728]} - {1'b0, layer_2_0[4735:4728]};
      btm_0[2] = {1'b0,layer_3_0[4743:4736]} - {1'b0, layer_2_0[4743:4736]};
      btm_1[0] = {1'b0,layer_3_1[4727:4720]} - {1'b0, layer_2_1[4727:4720]};
      btm_1[1] = {1'b0,layer_3_1[4735:4728]} - {1'b0, layer_2_1[4735:4728]};
      btm_1[2] = {1'b0,layer_3_1[4743:4736]} - {1'b0, layer_2_1[4743:4736]};
      btm_2[0] = {1'b0,layer_3_2[4727:4720]} - {1'b0, layer_2_2[4727:4720]};
      btm_2[1] = {1'b0,layer_3_2[4735:4728]} - {1'b0, layer_2_2[4735:4728]};
      btm_2[2] = {1'b0,layer_3_2[4743:4736]} - {1'b0, layer_2_2[4743:4736]};
    end
    'd592: begin
      top_0[0] = {1'b0,layer_1_0[4735:4728]} - {1'b0, layer_0_0[4735:4728]};
      top_0[1] = {1'b0,layer_1_0[4743:4736]} - {1'b0, layer_0_0[4743:4736]};
      top_0[2] = {1'b0,layer_1_0[4751:4744]} - {1'b0, layer_0_0[4751:4744]};
      top_1[0] = {1'b0,layer_1_1[4735:4728]} - {1'b0, layer_0_1[4735:4728]};
      top_1[1] = {1'b0,layer_1_1[4743:4736]} - {1'b0, layer_0_1[4743:4736]};
      top_1[2] = {1'b0,layer_1_1[4751:4744]} - {1'b0, layer_0_1[4751:4744]};
      top_2[0] = {1'b0,layer_1_2[4735:4728]} - {1'b0, layer_0_2[4735:4728]};
      top_2[1] = {1'b0,layer_1_2[4743:4736]} - {1'b0, layer_0_2[4743:4736]};
      top_2[2] = {1'b0,layer_1_2[4751:4744]} - {1'b0, layer_0_2[4751:4744]};
      mid_0[0] = {1'b0,layer_2_0[4735:4728]} - {1'b0, layer_1_0[4735:4728]};
      mid_0[1] = {1'b0,layer_2_0[4743:4736]} - {1'b0, layer_1_0[4743:4736]};
      mid_0[2] = {1'b0,layer_2_0[4751:4744]} - {1'b0, layer_1_0[4751:4744]};
      mid_1[0] = {1'b0,layer_2_1[4735:4728]} - {1'b0, layer_1_1[4735:4728]};
      mid_1[1] = {1'b0,layer_2_1[4743:4736]} - {1'b0, layer_1_1[4743:4736]};
      mid_1[2] = {1'b0,layer_2_1[4751:4744]} - {1'b0, layer_1_1[4751:4744]};
      mid_2[0] = {1'b0,layer_2_2[4735:4728]} - {1'b0, layer_1_2[4735:4728]};
      mid_2[1] = {1'b0,layer_2_2[4743:4736]} - {1'b0, layer_1_2[4743:4736]};
      mid_2[2] = {1'b0,layer_2_2[4751:4744]} - {1'b0, layer_1_2[4751:4744]};
      btm_0[0] = {1'b0,layer_3_0[4735:4728]} - {1'b0, layer_2_0[4735:4728]};
      btm_0[1] = {1'b0,layer_3_0[4743:4736]} - {1'b0, layer_2_0[4743:4736]};
      btm_0[2] = {1'b0,layer_3_0[4751:4744]} - {1'b0, layer_2_0[4751:4744]};
      btm_1[0] = {1'b0,layer_3_1[4735:4728]} - {1'b0, layer_2_1[4735:4728]};
      btm_1[1] = {1'b0,layer_3_1[4743:4736]} - {1'b0, layer_2_1[4743:4736]};
      btm_1[2] = {1'b0,layer_3_1[4751:4744]} - {1'b0, layer_2_1[4751:4744]};
      btm_2[0] = {1'b0,layer_3_2[4735:4728]} - {1'b0, layer_2_2[4735:4728]};
      btm_2[1] = {1'b0,layer_3_2[4743:4736]} - {1'b0, layer_2_2[4743:4736]};
      btm_2[2] = {1'b0,layer_3_2[4751:4744]} - {1'b0, layer_2_2[4751:4744]};
    end
    'd593: begin
      top_0[0] = {1'b0,layer_1_0[4743:4736]} - {1'b0, layer_0_0[4743:4736]};
      top_0[1] = {1'b0,layer_1_0[4751:4744]} - {1'b0, layer_0_0[4751:4744]};
      top_0[2] = {1'b0,layer_1_0[4759:4752]} - {1'b0, layer_0_0[4759:4752]};
      top_1[0] = {1'b0,layer_1_1[4743:4736]} - {1'b0, layer_0_1[4743:4736]};
      top_1[1] = {1'b0,layer_1_1[4751:4744]} - {1'b0, layer_0_1[4751:4744]};
      top_1[2] = {1'b0,layer_1_1[4759:4752]} - {1'b0, layer_0_1[4759:4752]};
      top_2[0] = {1'b0,layer_1_2[4743:4736]} - {1'b0, layer_0_2[4743:4736]};
      top_2[1] = {1'b0,layer_1_2[4751:4744]} - {1'b0, layer_0_2[4751:4744]};
      top_2[2] = {1'b0,layer_1_2[4759:4752]} - {1'b0, layer_0_2[4759:4752]};
      mid_0[0] = {1'b0,layer_2_0[4743:4736]} - {1'b0, layer_1_0[4743:4736]};
      mid_0[1] = {1'b0,layer_2_0[4751:4744]} - {1'b0, layer_1_0[4751:4744]};
      mid_0[2] = {1'b0,layer_2_0[4759:4752]} - {1'b0, layer_1_0[4759:4752]};
      mid_1[0] = {1'b0,layer_2_1[4743:4736]} - {1'b0, layer_1_1[4743:4736]};
      mid_1[1] = {1'b0,layer_2_1[4751:4744]} - {1'b0, layer_1_1[4751:4744]};
      mid_1[2] = {1'b0,layer_2_1[4759:4752]} - {1'b0, layer_1_1[4759:4752]};
      mid_2[0] = {1'b0,layer_2_2[4743:4736]} - {1'b0, layer_1_2[4743:4736]};
      mid_2[1] = {1'b0,layer_2_2[4751:4744]} - {1'b0, layer_1_2[4751:4744]};
      mid_2[2] = {1'b0,layer_2_2[4759:4752]} - {1'b0, layer_1_2[4759:4752]};
      btm_0[0] = {1'b0,layer_3_0[4743:4736]} - {1'b0, layer_2_0[4743:4736]};
      btm_0[1] = {1'b0,layer_3_0[4751:4744]} - {1'b0, layer_2_0[4751:4744]};
      btm_0[2] = {1'b0,layer_3_0[4759:4752]} - {1'b0, layer_2_0[4759:4752]};
      btm_1[0] = {1'b0,layer_3_1[4743:4736]} - {1'b0, layer_2_1[4743:4736]};
      btm_1[1] = {1'b0,layer_3_1[4751:4744]} - {1'b0, layer_2_1[4751:4744]};
      btm_1[2] = {1'b0,layer_3_1[4759:4752]} - {1'b0, layer_2_1[4759:4752]};
      btm_2[0] = {1'b0,layer_3_2[4743:4736]} - {1'b0, layer_2_2[4743:4736]};
      btm_2[1] = {1'b0,layer_3_2[4751:4744]} - {1'b0, layer_2_2[4751:4744]};
      btm_2[2] = {1'b0,layer_3_2[4759:4752]} - {1'b0, layer_2_2[4759:4752]};
    end
    'd594: begin
      top_0[0] = {1'b0,layer_1_0[4751:4744]} - {1'b0, layer_0_0[4751:4744]};
      top_0[1] = {1'b0,layer_1_0[4759:4752]} - {1'b0, layer_0_0[4759:4752]};
      top_0[2] = {1'b0,layer_1_0[4767:4760]} - {1'b0, layer_0_0[4767:4760]};
      top_1[0] = {1'b0,layer_1_1[4751:4744]} - {1'b0, layer_0_1[4751:4744]};
      top_1[1] = {1'b0,layer_1_1[4759:4752]} - {1'b0, layer_0_1[4759:4752]};
      top_1[2] = {1'b0,layer_1_1[4767:4760]} - {1'b0, layer_0_1[4767:4760]};
      top_2[0] = {1'b0,layer_1_2[4751:4744]} - {1'b0, layer_0_2[4751:4744]};
      top_2[1] = {1'b0,layer_1_2[4759:4752]} - {1'b0, layer_0_2[4759:4752]};
      top_2[2] = {1'b0,layer_1_2[4767:4760]} - {1'b0, layer_0_2[4767:4760]};
      mid_0[0] = {1'b0,layer_2_0[4751:4744]} - {1'b0, layer_1_0[4751:4744]};
      mid_0[1] = {1'b0,layer_2_0[4759:4752]} - {1'b0, layer_1_0[4759:4752]};
      mid_0[2] = {1'b0,layer_2_0[4767:4760]} - {1'b0, layer_1_0[4767:4760]};
      mid_1[0] = {1'b0,layer_2_1[4751:4744]} - {1'b0, layer_1_1[4751:4744]};
      mid_1[1] = {1'b0,layer_2_1[4759:4752]} - {1'b0, layer_1_1[4759:4752]};
      mid_1[2] = {1'b0,layer_2_1[4767:4760]} - {1'b0, layer_1_1[4767:4760]};
      mid_2[0] = {1'b0,layer_2_2[4751:4744]} - {1'b0, layer_1_2[4751:4744]};
      mid_2[1] = {1'b0,layer_2_2[4759:4752]} - {1'b0, layer_1_2[4759:4752]};
      mid_2[2] = {1'b0,layer_2_2[4767:4760]} - {1'b0, layer_1_2[4767:4760]};
      btm_0[0] = {1'b0,layer_3_0[4751:4744]} - {1'b0, layer_2_0[4751:4744]};
      btm_0[1] = {1'b0,layer_3_0[4759:4752]} - {1'b0, layer_2_0[4759:4752]};
      btm_0[2] = {1'b0,layer_3_0[4767:4760]} - {1'b0, layer_2_0[4767:4760]};
      btm_1[0] = {1'b0,layer_3_1[4751:4744]} - {1'b0, layer_2_1[4751:4744]};
      btm_1[1] = {1'b0,layer_3_1[4759:4752]} - {1'b0, layer_2_1[4759:4752]};
      btm_1[2] = {1'b0,layer_3_1[4767:4760]} - {1'b0, layer_2_1[4767:4760]};
      btm_2[0] = {1'b0,layer_3_2[4751:4744]} - {1'b0, layer_2_2[4751:4744]};
      btm_2[1] = {1'b0,layer_3_2[4759:4752]} - {1'b0, layer_2_2[4759:4752]};
      btm_2[2] = {1'b0,layer_3_2[4767:4760]} - {1'b0, layer_2_2[4767:4760]};
    end
    'd595: begin
      top_0[0] = {1'b0,layer_1_0[4759:4752]} - {1'b0, layer_0_0[4759:4752]};
      top_0[1] = {1'b0,layer_1_0[4767:4760]} - {1'b0, layer_0_0[4767:4760]};
      top_0[2] = {1'b0,layer_1_0[4775:4768]} - {1'b0, layer_0_0[4775:4768]};
      top_1[0] = {1'b0,layer_1_1[4759:4752]} - {1'b0, layer_0_1[4759:4752]};
      top_1[1] = {1'b0,layer_1_1[4767:4760]} - {1'b0, layer_0_1[4767:4760]};
      top_1[2] = {1'b0,layer_1_1[4775:4768]} - {1'b0, layer_0_1[4775:4768]};
      top_2[0] = {1'b0,layer_1_2[4759:4752]} - {1'b0, layer_0_2[4759:4752]};
      top_2[1] = {1'b0,layer_1_2[4767:4760]} - {1'b0, layer_0_2[4767:4760]};
      top_2[2] = {1'b0,layer_1_2[4775:4768]} - {1'b0, layer_0_2[4775:4768]};
      mid_0[0] = {1'b0,layer_2_0[4759:4752]} - {1'b0, layer_1_0[4759:4752]};
      mid_0[1] = {1'b0,layer_2_0[4767:4760]} - {1'b0, layer_1_0[4767:4760]};
      mid_0[2] = {1'b0,layer_2_0[4775:4768]} - {1'b0, layer_1_0[4775:4768]};
      mid_1[0] = {1'b0,layer_2_1[4759:4752]} - {1'b0, layer_1_1[4759:4752]};
      mid_1[1] = {1'b0,layer_2_1[4767:4760]} - {1'b0, layer_1_1[4767:4760]};
      mid_1[2] = {1'b0,layer_2_1[4775:4768]} - {1'b0, layer_1_1[4775:4768]};
      mid_2[0] = {1'b0,layer_2_2[4759:4752]} - {1'b0, layer_1_2[4759:4752]};
      mid_2[1] = {1'b0,layer_2_2[4767:4760]} - {1'b0, layer_1_2[4767:4760]};
      mid_2[2] = {1'b0,layer_2_2[4775:4768]} - {1'b0, layer_1_2[4775:4768]};
      btm_0[0] = {1'b0,layer_3_0[4759:4752]} - {1'b0, layer_2_0[4759:4752]};
      btm_0[1] = {1'b0,layer_3_0[4767:4760]} - {1'b0, layer_2_0[4767:4760]};
      btm_0[2] = {1'b0,layer_3_0[4775:4768]} - {1'b0, layer_2_0[4775:4768]};
      btm_1[0] = {1'b0,layer_3_1[4759:4752]} - {1'b0, layer_2_1[4759:4752]};
      btm_1[1] = {1'b0,layer_3_1[4767:4760]} - {1'b0, layer_2_1[4767:4760]};
      btm_1[2] = {1'b0,layer_3_1[4775:4768]} - {1'b0, layer_2_1[4775:4768]};
      btm_2[0] = {1'b0,layer_3_2[4759:4752]} - {1'b0, layer_2_2[4759:4752]};
      btm_2[1] = {1'b0,layer_3_2[4767:4760]} - {1'b0, layer_2_2[4767:4760]};
      btm_2[2] = {1'b0,layer_3_2[4775:4768]} - {1'b0, layer_2_2[4775:4768]};
    end
    'd596: begin
      top_0[0] = {1'b0,layer_1_0[4767:4760]} - {1'b0, layer_0_0[4767:4760]};
      top_0[1] = {1'b0,layer_1_0[4775:4768]} - {1'b0, layer_0_0[4775:4768]};
      top_0[2] = {1'b0,layer_1_0[4783:4776]} - {1'b0, layer_0_0[4783:4776]};
      top_1[0] = {1'b0,layer_1_1[4767:4760]} - {1'b0, layer_0_1[4767:4760]};
      top_1[1] = {1'b0,layer_1_1[4775:4768]} - {1'b0, layer_0_1[4775:4768]};
      top_1[2] = {1'b0,layer_1_1[4783:4776]} - {1'b0, layer_0_1[4783:4776]};
      top_2[0] = {1'b0,layer_1_2[4767:4760]} - {1'b0, layer_0_2[4767:4760]};
      top_2[1] = {1'b0,layer_1_2[4775:4768]} - {1'b0, layer_0_2[4775:4768]};
      top_2[2] = {1'b0,layer_1_2[4783:4776]} - {1'b0, layer_0_2[4783:4776]};
      mid_0[0] = {1'b0,layer_2_0[4767:4760]} - {1'b0, layer_1_0[4767:4760]};
      mid_0[1] = {1'b0,layer_2_0[4775:4768]} - {1'b0, layer_1_0[4775:4768]};
      mid_0[2] = {1'b0,layer_2_0[4783:4776]} - {1'b0, layer_1_0[4783:4776]};
      mid_1[0] = {1'b0,layer_2_1[4767:4760]} - {1'b0, layer_1_1[4767:4760]};
      mid_1[1] = {1'b0,layer_2_1[4775:4768]} - {1'b0, layer_1_1[4775:4768]};
      mid_1[2] = {1'b0,layer_2_1[4783:4776]} - {1'b0, layer_1_1[4783:4776]};
      mid_2[0] = {1'b0,layer_2_2[4767:4760]} - {1'b0, layer_1_2[4767:4760]};
      mid_2[1] = {1'b0,layer_2_2[4775:4768]} - {1'b0, layer_1_2[4775:4768]};
      mid_2[2] = {1'b0,layer_2_2[4783:4776]} - {1'b0, layer_1_2[4783:4776]};
      btm_0[0] = {1'b0,layer_3_0[4767:4760]} - {1'b0, layer_2_0[4767:4760]};
      btm_0[1] = {1'b0,layer_3_0[4775:4768]} - {1'b0, layer_2_0[4775:4768]};
      btm_0[2] = {1'b0,layer_3_0[4783:4776]} - {1'b0, layer_2_0[4783:4776]};
      btm_1[0] = {1'b0,layer_3_1[4767:4760]} - {1'b0, layer_2_1[4767:4760]};
      btm_1[1] = {1'b0,layer_3_1[4775:4768]} - {1'b0, layer_2_1[4775:4768]};
      btm_1[2] = {1'b0,layer_3_1[4783:4776]} - {1'b0, layer_2_1[4783:4776]};
      btm_2[0] = {1'b0,layer_3_2[4767:4760]} - {1'b0, layer_2_2[4767:4760]};
      btm_2[1] = {1'b0,layer_3_2[4775:4768]} - {1'b0, layer_2_2[4775:4768]};
      btm_2[2] = {1'b0,layer_3_2[4783:4776]} - {1'b0, layer_2_2[4783:4776]};
    end
    'd597: begin
      top_0[0] = {1'b0,layer_1_0[4775:4768]} - {1'b0, layer_0_0[4775:4768]};
      top_0[1] = {1'b0,layer_1_0[4783:4776]} - {1'b0, layer_0_0[4783:4776]};
      top_0[2] = {1'b0,layer_1_0[4791:4784]} - {1'b0, layer_0_0[4791:4784]};
      top_1[0] = {1'b0,layer_1_1[4775:4768]} - {1'b0, layer_0_1[4775:4768]};
      top_1[1] = {1'b0,layer_1_1[4783:4776]} - {1'b0, layer_0_1[4783:4776]};
      top_1[2] = {1'b0,layer_1_1[4791:4784]} - {1'b0, layer_0_1[4791:4784]};
      top_2[0] = {1'b0,layer_1_2[4775:4768]} - {1'b0, layer_0_2[4775:4768]};
      top_2[1] = {1'b0,layer_1_2[4783:4776]} - {1'b0, layer_0_2[4783:4776]};
      top_2[2] = {1'b0,layer_1_2[4791:4784]} - {1'b0, layer_0_2[4791:4784]};
      mid_0[0] = {1'b0,layer_2_0[4775:4768]} - {1'b0, layer_1_0[4775:4768]};
      mid_0[1] = {1'b0,layer_2_0[4783:4776]} - {1'b0, layer_1_0[4783:4776]};
      mid_0[2] = {1'b0,layer_2_0[4791:4784]} - {1'b0, layer_1_0[4791:4784]};
      mid_1[0] = {1'b0,layer_2_1[4775:4768]} - {1'b0, layer_1_1[4775:4768]};
      mid_1[1] = {1'b0,layer_2_1[4783:4776]} - {1'b0, layer_1_1[4783:4776]};
      mid_1[2] = {1'b0,layer_2_1[4791:4784]} - {1'b0, layer_1_1[4791:4784]};
      mid_2[0] = {1'b0,layer_2_2[4775:4768]} - {1'b0, layer_1_2[4775:4768]};
      mid_2[1] = {1'b0,layer_2_2[4783:4776]} - {1'b0, layer_1_2[4783:4776]};
      mid_2[2] = {1'b0,layer_2_2[4791:4784]} - {1'b0, layer_1_2[4791:4784]};
      btm_0[0] = {1'b0,layer_3_0[4775:4768]} - {1'b0, layer_2_0[4775:4768]};
      btm_0[1] = {1'b0,layer_3_0[4783:4776]} - {1'b0, layer_2_0[4783:4776]};
      btm_0[2] = {1'b0,layer_3_0[4791:4784]} - {1'b0, layer_2_0[4791:4784]};
      btm_1[0] = {1'b0,layer_3_1[4775:4768]} - {1'b0, layer_2_1[4775:4768]};
      btm_1[1] = {1'b0,layer_3_1[4783:4776]} - {1'b0, layer_2_1[4783:4776]};
      btm_1[2] = {1'b0,layer_3_1[4791:4784]} - {1'b0, layer_2_1[4791:4784]};
      btm_2[0] = {1'b0,layer_3_2[4775:4768]} - {1'b0, layer_2_2[4775:4768]};
      btm_2[1] = {1'b0,layer_3_2[4783:4776]} - {1'b0, layer_2_2[4783:4776]};
      btm_2[2] = {1'b0,layer_3_2[4791:4784]} - {1'b0, layer_2_2[4791:4784]};
    end
    'd598: begin
      top_0[0] = {1'b0,layer_1_0[4783:4776]} - {1'b0, layer_0_0[4783:4776]};
      top_0[1] = {1'b0,layer_1_0[4791:4784]} - {1'b0, layer_0_0[4791:4784]};
      top_0[2] = {1'b0,layer_1_0[4799:4792]} - {1'b0, layer_0_0[4799:4792]};
      top_1[0] = {1'b0,layer_1_1[4783:4776]} - {1'b0, layer_0_1[4783:4776]};
      top_1[1] = {1'b0,layer_1_1[4791:4784]} - {1'b0, layer_0_1[4791:4784]};
      top_1[2] = {1'b0,layer_1_1[4799:4792]} - {1'b0, layer_0_1[4799:4792]};
      top_2[0] = {1'b0,layer_1_2[4783:4776]} - {1'b0, layer_0_2[4783:4776]};
      top_2[1] = {1'b0,layer_1_2[4791:4784]} - {1'b0, layer_0_2[4791:4784]};
      top_2[2] = {1'b0,layer_1_2[4799:4792]} - {1'b0, layer_0_2[4799:4792]};
      mid_0[0] = {1'b0,layer_2_0[4783:4776]} - {1'b0, layer_1_0[4783:4776]};
      mid_0[1] = {1'b0,layer_2_0[4791:4784]} - {1'b0, layer_1_0[4791:4784]};
      mid_0[2] = {1'b0,layer_2_0[4799:4792]} - {1'b0, layer_1_0[4799:4792]};
      mid_1[0] = {1'b0,layer_2_1[4783:4776]} - {1'b0, layer_1_1[4783:4776]};
      mid_1[1] = {1'b0,layer_2_1[4791:4784]} - {1'b0, layer_1_1[4791:4784]};
      mid_1[2] = {1'b0,layer_2_1[4799:4792]} - {1'b0, layer_1_1[4799:4792]};
      mid_2[0] = {1'b0,layer_2_2[4783:4776]} - {1'b0, layer_1_2[4783:4776]};
      mid_2[1] = {1'b0,layer_2_2[4791:4784]} - {1'b0, layer_1_2[4791:4784]};
      mid_2[2] = {1'b0,layer_2_2[4799:4792]} - {1'b0, layer_1_2[4799:4792]};
      btm_0[0] = {1'b0,layer_3_0[4783:4776]} - {1'b0, layer_2_0[4783:4776]};
      btm_0[1] = {1'b0,layer_3_0[4791:4784]} - {1'b0, layer_2_0[4791:4784]};
      btm_0[2] = {1'b0,layer_3_0[4799:4792]} - {1'b0, layer_2_0[4799:4792]};
      btm_1[0] = {1'b0,layer_3_1[4783:4776]} - {1'b0, layer_2_1[4783:4776]};
      btm_1[1] = {1'b0,layer_3_1[4791:4784]} - {1'b0, layer_2_1[4791:4784]};
      btm_1[2] = {1'b0,layer_3_1[4799:4792]} - {1'b0, layer_2_1[4799:4792]};
      btm_2[0] = {1'b0,layer_3_2[4783:4776]} - {1'b0, layer_2_2[4783:4776]};
      btm_2[1] = {1'b0,layer_3_2[4791:4784]} - {1'b0, layer_2_2[4791:4784]};
      btm_2[2] = {1'b0,layer_3_2[4799:4792]} - {1'b0, layer_2_2[4799:4792]};
    end
    'd599: begin
      top_0[0] = {1'b0,layer_1_0[4791:4784]} - {1'b0, layer_0_0[4791:4784]};
      top_0[1] = {1'b0,layer_1_0[4799:4792]} - {1'b0, layer_0_0[4799:4792]};
      top_0[2] = {1'b0,layer_1_0[4807:4800]} - {1'b0, layer_0_0[4807:4800]};
      top_1[0] = {1'b0,layer_1_1[4791:4784]} - {1'b0, layer_0_1[4791:4784]};
      top_1[1] = {1'b0,layer_1_1[4799:4792]} - {1'b0, layer_0_1[4799:4792]};
      top_1[2] = {1'b0,layer_1_1[4807:4800]} - {1'b0, layer_0_1[4807:4800]};
      top_2[0] = {1'b0,layer_1_2[4791:4784]} - {1'b0, layer_0_2[4791:4784]};
      top_2[1] = {1'b0,layer_1_2[4799:4792]} - {1'b0, layer_0_2[4799:4792]};
      top_2[2] = {1'b0,layer_1_2[4807:4800]} - {1'b0, layer_0_2[4807:4800]};
      mid_0[0] = {1'b0,layer_2_0[4791:4784]} - {1'b0, layer_1_0[4791:4784]};
      mid_0[1] = {1'b0,layer_2_0[4799:4792]} - {1'b0, layer_1_0[4799:4792]};
      mid_0[2] = {1'b0,layer_2_0[4807:4800]} - {1'b0, layer_1_0[4807:4800]};
      mid_1[0] = {1'b0,layer_2_1[4791:4784]} - {1'b0, layer_1_1[4791:4784]};
      mid_1[1] = {1'b0,layer_2_1[4799:4792]} - {1'b0, layer_1_1[4799:4792]};
      mid_1[2] = {1'b0,layer_2_1[4807:4800]} - {1'b0, layer_1_1[4807:4800]};
      mid_2[0] = {1'b0,layer_2_2[4791:4784]} - {1'b0, layer_1_2[4791:4784]};
      mid_2[1] = {1'b0,layer_2_2[4799:4792]} - {1'b0, layer_1_2[4799:4792]};
      mid_2[2] = {1'b0,layer_2_2[4807:4800]} - {1'b0, layer_1_2[4807:4800]};
      btm_0[0] = {1'b0,layer_3_0[4791:4784]} - {1'b0, layer_2_0[4791:4784]};
      btm_0[1] = {1'b0,layer_3_0[4799:4792]} - {1'b0, layer_2_0[4799:4792]};
      btm_0[2] = {1'b0,layer_3_0[4807:4800]} - {1'b0, layer_2_0[4807:4800]};
      btm_1[0] = {1'b0,layer_3_1[4791:4784]} - {1'b0, layer_2_1[4791:4784]};
      btm_1[1] = {1'b0,layer_3_1[4799:4792]} - {1'b0, layer_2_1[4799:4792]};
      btm_1[2] = {1'b0,layer_3_1[4807:4800]} - {1'b0, layer_2_1[4807:4800]};
      btm_2[0] = {1'b0,layer_3_2[4791:4784]} - {1'b0, layer_2_2[4791:4784]};
      btm_2[1] = {1'b0,layer_3_2[4799:4792]} - {1'b0, layer_2_2[4799:4792]};
      btm_2[2] = {1'b0,layer_3_2[4807:4800]} - {1'b0, layer_2_2[4807:4800]};
    end
    'd600: begin
      top_0[0] = {1'b0,layer_1_0[4799:4792]} - {1'b0, layer_0_0[4799:4792]};
      top_0[1] = {1'b0,layer_1_0[4807:4800]} - {1'b0, layer_0_0[4807:4800]};
      top_0[2] = {1'b0,layer_1_0[4815:4808]} - {1'b0, layer_0_0[4815:4808]};
      top_1[0] = {1'b0,layer_1_1[4799:4792]} - {1'b0, layer_0_1[4799:4792]};
      top_1[1] = {1'b0,layer_1_1[4807:4800]} - {1'b0, layer_0_1[4807:4800]};
      top_1[2] = {1'b0,layer_1_1[4815:4808]} - {1'b0, layer_0_1[4815:4808]};
      top_2[0] = {1'b0,layer_1_2[4799:4792]} - {1'b0, layer_0_2[4799:4792]};
      top_2[1] = {1'b0,layer_1_2[4807:4800]} - {1'b0, layer_0_2[4807:4800]};
      top_2[2] = {1'b0,layer_1_2[4815:4808]} - {1'b0, layer_0_2[4815:4808]};
      mid_0[0] = {1'b0,layer_2_0[4799:4792]} - {1'b0, layer_1_0[4799:4792]};
      mid_0[1] = {1'b0,layer_2_0[4807:4800]} - {1'b0, layer_1_0[4807:4800]};
      mid_0[2] = {1'b0,layer_2_0[4815:4808]} - {1'b0, layer_1_0[4815:4808]};
      mid_1[0] = {1'b0,layer_2_1[4799:4792]} - {1'b0, layer_1_1[4799:4792]};
      mid_1[1] = {1'b0,layer_2_1[4807:4800]} - {1'b0, layer_1_1[4807:4800]};
      mid_1[2] = {1'b0,layer_2_1[4815:4808]} - {1'b0, layer_1_1[4815:4808]};
      mid_2[0] = {1'b0,layer_2_2[4799:4792]} - {1'b0, layer_1_2[4799:4792]};
      mid_2[1] = {1'b0,layer_2_2[4807:4800]} - {1'b0, layer_1_2[4807:4800]};
      mid_2[2] = {1'b0,layer_2_2[4815:4808]} - {1'b0, layer_1_2[4815:4808]};
      btm_0[0] = {1'b0,layer_3_0[4799:4792]} - {1'b0, layer_2_0[4799:4792]};
      btm_0[1] = {1'b0,layer_3_0[4807:4800]} - {1'b0, layer_2_0[4807:4800]};
      btm_0[2] = {1'b0,layer_3_0[4815:4808]} - {1'b0, layer_2_0[4815:4808]};
      btm_1[0] = {1'b0,layer_3_1[4799:4792]} - {1'b0, layer_2_1[4799:4792]};
      btm_1[1] = {1'b0,layer_3_1[4807:4800]} - {1'b0, layer_2_1[4807:4800]};
      btm_1[2] = {1'b0,layer_3_1[4815:4808]} - {1'b0, layer_2_1[4815:4808]};
      btm_2[0] = {1'b0,layer_3_2[4799:4792]} - {1'b0, layer_2_2[4799:4792]};
      btm_2[1] = {1'b0,layer_3_2[4807:4800]} - {1'b0, layer_2_2[4807:4800]};
      btm_2[2] = {1'b0,layer_3_2[4815:4808]} - {1'b0, layer_2_2[4815:4808]};
    end
    'd601: begin
      top_0[0] = {1'b0,layer_1_0[4807:4800]} - {1'b0, layer_0_0[4807:4800]};
      top_0[1] = {1'b0,layer_1_0[4815:4808]} - {1'b0, layer_0_0[4815:4808]};
      top_0[2] = {1'b0,layer_1_0[4823:4816]} - {1'b0, layer_0_0[4823:4816]};
      top_1[0] = {1'b0,layer_1_1[4807:4800]} - {1'b0, layer_0_1[4807:4800]};
      top_1[1] = {1'b0,layer_1_1[4815:4808]} - {1'b0, layer_0_1[4815:4808]};
      top_1[2] = {1'b0,layer_1_1[4823:4816]} - {1'b0, layer_0_1[4823:4816]};
      top_2[0] = {1'b0,layer_1_2[4807:4800]} - {1'b0, layer_0_2[4807:4800]};
      top_2[1] = {1'b0,layer_1_2[4815:4808]} - {1'b0, layer_0_2[4815:4808]};
      top_2[2] = {1'b0,layer_1_2[4823:4816]} - {1'b0, layer_0_2[4823:4816]};
      mid_0[0] = {1'b0,layer_2_0[4807:4800]} - {1'b0, layer_1_0[4807:4800]};
      mid_0[1] = {1'b0,layer_2_0[4815:4808]} - {1'b0, layer_1_0[4815:4808]};
      mid_0[2] = {1'b0,layer_2_0[4823:4816]} - {1'b0, layer_1_0[4823:4816]};
      mid_1[0] = {1'b0,layer_2_1[4807:4800]} - {1'b0, layer_1_1[4807:4800]};
      mid_1[1] = {1'b0,layer_2_1[4815:4808]} - {1'b0, layer_1_1[4815:4808]};
      mid_1[2] = {1'b0,layer_2_1[4823:4816]} - {1'b0, layer_1_1[4823:4816]};
      mid_2[0] = {1'b0,layer_2_2[4807:4800]} - {1'b0, layer_1_2[4807:4800]};
      mid_2[1] = {1'b0,layer_2_2[4815:4808]} - {1'b0, layer_1_2[4815:4808]};
      mid_2[2] = {1'b0,layer_2_2[4823:4816]} - {1'b0, layer_1_2[4823:4816]};
      btm_0[0] = {1'b0,layer_3_0[4807:4800]} - {1'b0, layer_2_0[4807:4800]};
      btm_0[1] = {1'b0,layer_3_0[4815:4808]} - {1'b0, layer_2_0[4815:4808]};
      btm_0[2] = {1'b0,layer_3_0[4823:4816]} - {1'b0, layer_2_0[4823:4816]};
      btm_1[0] = {1'b0,layer_3_1[4807:4800]} - {1'b0, layer_2_1[4807:4800]};
      btm_1[1] = {1'b0,layer_3_1[4815:4808]} - {1'b0, layer_2_1[4815:4808]};
      btm_1[2] = {1'b0,layer_3_1[4823:4816]} - {1'b0, layer_2_1[4823:4816]};
      btm_2[0] = {1'b0,layer_3_2[4807:4800]} - {1'b0, layer_2_2[4807:4800]};
      btm_2[1] = {1'b0,layer_3_2[4815:4808]} - {1'b0, layer_2_2[4815:4808]};
      btm_2[2] = {1'b0,layer_3_2[4823:4816]} - {1'b0, layer_2_2[4823:4816]};
    end
    'd602: begin
      top_0[0] = {1'b0,layer_1_0[4815:4808]} - {1'b0, layer_0_0[4815:4808]};
      top_0[1] = {1'b0,layer_1_0[4823:4816]} - {1'b0, layer_0_0[4823:4816]};
      top_0[2] = {1'b0,layer_1_0[4831:4824]} - {1'b0, layer_0_0[4831:4824]};
      top_1[0] = {1'b0,layer_1_1[4815:4808]} - {1'b0, layer_0_1[4815:4808]};
      top_1[1] = {1'b0,layer_1_1[4823:4816]} - {1'b0, layer_0_1[4823:4816]};
      top_1[2] = {1'b0,layer_1_1[4831:4824]} - {1'b0, layer_0_1[4831:4824]};
      top_2[0] = {1'b0,layer_1_2[4815:4808]} - {1'b0, layer_0_2[4815:4808]};
      top_2[1] = {1'b0,layer_1_2[4823:4816]} - {1'b0, layer_0_2[4823:4816]};
      top_2[2] = {1'b0,layer_1_2[4831:4824]} - {1'b0, layer_0_2[4831:4824]};
      mid_0[0] = {1'b0,layer_2_0[4815:4808]} - {1'b0, layer_1_0[4815:4808]};
      mid_0[1] = {1'b0,layer_2_0[4823:4816]} - {1'b0, layer_1_0[4823:4816]};
      mid_0[2] = {1'b0,layer_2_0[4831:4824]} - {1'b0, layer_1_0[4831:4824]};
      mid_1[0] = {1'b0,layer_2_1[4815:4808]} - {1'b0, layer_1_1[4815:4808]};
      mid_1[1] = {1'b0,layer_2_1[4823:4816]} - {1'b0, layer_1_1[4823:4816]};
      mid_1[2] = {1'b0,layer_2_1[4831:4824]} - {1'b0, layer_1_1[4831:4824]};
      mid_2[0] = {1'b0,layer_2_2[4815:4808]} - {1'b0, layer_1_2[4815:4808]};
      mid_2[1] = {1'b0,layer_2_2[4823:4816]} - {1'b0, layer_1_2[4823:4816]};
      mid_2[2] = {1'b0,layer_2_2[4831:4824]} - {1'b0, layer_1_2[4831:4824]};
      btm_0[0] = {1'b0,layer_3_0[4815:4808]} - {1'b0, layer_2_0[4815:4808]};
      btm_0[1] = {1'b0,layer_3_0[4823:4816]} - {1'b0, layer_2_0[4823:4816]};
      btm_0[2] = {1'b0,layer_3_0[4831:4824]} - {1'b0, layer_2_0[4831:4824]};
      btm_1[0] = {1'b0,layer_3_1[4815:4808]} - {1'b0, layer_2_1[4815:4808]};
      btm_1[1] = {1'b0,layer_3_1[4823:4816]} - {1'b0, layer_2_1[4823:4816]};
      btm_1[2] = {1'b0,layer_3_1[4831:4824]} - {1'b0, layer_2_1[4831:4824]};
      btm_2[0] = {1'b0,layer_3_2[4815:4808]} - {1'b0, layer_2_2[4815:4808]};
      btm_2[1] = {1'b0,layer_3_2[4823:4816]} - {1'b0, layer_2_2[4823:4816]};
      btm_2[2] = {1'b0,layer_3_2[4831:4824]} - {1'b0, layer_2_2[4831:4824]};
    end
    'd603: begin
      top_0[0] = {1'b0,layer_1_0[4823:4816]} - {1'b0, layer_0_0[4823:4816]};
      top_0[1] = {1'b0,layer_1_0[4831:4824]} - {1'b0, layer_0_0[4831:4824]};
      top_0[2] = {1'b0,layer_1_0[4839:4832]} - {1'b0, layer_0_0[4839:4832]};
      top_1[0] = {1'b0,layer_1_1[4823:4816]} - {1'b0, layer_0_1[4823:4816]};
      top_1[1] = {1'b0,layer_1_1[4831:4824]} - {1'b0, layer_0_1[4831:4824]};
      top_1[2] = {1'b0,layer_1_1[4839:4832]} - {1'b0, layer_0_1[4839:4832]};
      top_2[0] = {1'b0,layer_1_2[4823:4816]} - {1'b0, layer_0_2[4823:4816]};
      top_2[1] = {1'b0,layer_1_2[4831:4824]} - {1'b0, layer_0_2[4831:4824]};
      top_2[2] = {1'b0,layer_1_2[4839:4832]} - {1'b0, layer_0_2[4839:4832]};
      mid_0[0] = {1'b0,layer_2_0[4823:4816]} - {1'b0, layer_1_0[4823:4816]};
      mid_0[1] = {1'b0,layer_2_0[4831:4824]} - {1'b0, layer_1_0[4831:4824]};
      mid_0[2] = {1'b0,layer_2_0[4839:4832]} - {1'b0, layer_1_0[4839:4832]};
      mid_1[0] = {1'b0,layer_2_1[4823:4816]} - {1'b0, layer_1_1[4823:4816]};
      mid_1[1] = {1'b0,layer_2_1[4831:4824]} - {1'b0, layer_1_1[4831:4824]};
      mid_1[2] = {1'b0,layer_2_1[4839:4832]} - {1'b0, layer_1_1[4839:4832]};
      mid_2[0] = {1'b0,layer_2_2[4823:4816]} - {1'b0, layer_1_2[4823:4816]};
      mid_2[1] = {1'b0,layer_2_2[4831:4824]} - {1'b0, layer_1_2[4831:4824]};
      mid_2[2] = {1'b0,layer_2_2[4839:4832]} - {1'b0, layer_1_2[4839:4832]};
      btm_0[0] = {1'b0,layer_3_0[4823:4816]} - {1'b0, layer_2_0[4823:4816]};
      btm_0[1] = {1'b0,layer_3_0[4831:4824]} - {1'b0, layer_2_0[4831:4824]};
      btm_0[2] = {1'b0,layer_3_0[4839:4832]} - {1'b0, layer_2_0[4839:4832]};
      btm_1[0] = {1'b0,layer_3_1[4823:4816]} - {1'b0, layer_2_1[4823:4816]};
      btm_1[1] = {1'b0,layer_3_1[4831:4824]} - {1'b0, layer_2_1[4831:4824]};
      btm_1[2] = {1'b0,layer_3_1[4839:4832]} - {1'b0, layer_2_1[4839:4832]};
      btm_2[0] = {1'b0,layer_3_2[4823:4816]} - {1'b0, layer_2_2[4823:4816]};
      btm_2[1] = {1'b0,layer_3_2[4831:4824]} - {1'b0, layer_2_2[4831:4824]};
      btm_2[2] = {1'b0,layer_3_2[4839:4832]} - {1'b0, layer_2_2[4839:4832]};
    end
    'd604: begin
      top_0[0] = {1'b0,layer_1_0[4831:4824]} - {1'b0, layer_0_0[4831:4824]};
      top_0[1] = {1'b0,layer_1_0[4839:4832]} - {1'b0, layer_0_0[4839:4832]};
      top_0[2] = {1'b0,layer_1_0[4847:4840]} - {1'b0, layer_0_0[4847:4840]};
      top_1[0] = {1'b0,layer_1_1[4831:4824]} - {1'b0, layer_0_1[4831:4824]};
      top_1[1] = {1'b0,layer_1_1[4839:4832]} - {1'b0, layer_0_1[4839:4832]};
      top_1[2] = {1'b0,layer_1_1[4847:4840]} - {1'b0, layer_0_1[4847:4840]};
      top_2[0] = {1'b0,layer_1_2[4831:4824]} - {1'b0, layer_0_2[4831:4824]};
      top_2[1] = {1'b0,layer_1_2[4839:4832]} - {1'b0, layer_0_2[4839:4832]};
      top_2[2] = {1'b0,layer_1_2[4847:4840]} - {1'b0, layer_0_2[4847:4840]};
      mid_0[0] = {1'b0,layer_2_0[4831:4824]} - {1'b0, layer_1_0[4831:4824]};
      mid_0[1] = {1'b0,layer_2_0[4839:4832]} - {1'b0, layer_1_0[4839:4832]};
      mid_0[2] = {1'b0,layer_2_0[4847:4840]} - {1'b0, layer_1_0[4847:4840]};
      mid_1[0] = {1'b0,layer_2_1[4831:4824]} - {1'b0, layer_1_1[4831:4824]};
      mid_1[1] = {1'b0,layer_2_1[4839:4832]} - {1'b0, layer_1_1[4839:4832]};
      mid_1[2] = {1'b0,layer_2_1[4847:4840]} - {1'b0, layer_1_1[4847:4840]};
      mid_2[0] = {1'b0,layer_2_2[4831:4824]} - {1'b0, layer_1_2[4831:4824]};
      mid_2[1] = {1'b0,layer_2_2[4839:4832]} - {1'b0, layer_1_2[4839:4832]};
      mid_2[2] = {1'b0,layer_2_2[4847:4840]} - {1'b0, layer_1_2[4847:4840]};
      btm_0[0] = {1'b0,layer_3_0[4831:4824]} - {1'b0, layer_2_0[4831:4824]};
      btm_0[1] = {1'b0,layer_3_0[4839:4832]} - {1'b0, layer_2_0[4839:4832]};
      btm_0[2] = {1'b0,layer_3_0[4847:4840]} - {1'b0, layer_2_0[4847:4840]};
      btm_1[0] = {1'b0,layer_3_1[4831:4824]} - {1'b0, layer_2_1[4831:4824]};
      btm_1[1] = {1'b0,layer_3_1[4839:4832]} - {1'b0, layer_2_1[4839:4832]};
      btm_1[2] = {1'b0,layer_3_1[4847:4840]} - {1'b0, layer_2_1[4847:4840]};
      btm_2[0] = {1'b0,layer_3_2[4831:4824]} - {1'b0, layer_2_2[4831:4824]};
      btm_2[1] = {1'b0,layer_3_2[4839:4832]} - {1'b0, layer_2_2[4839:4832]};
      btm_2[2] = {1'b0,layer_3_2[4847:4840]} - {1'b0, layer_2_2[4847:4840]};
    end
    'd605: begin
      top_0[0] = {1'b0,layer_1_0[4839:4832]} - {1'b0, layer_0_0[4839:4832]};
      top_0[1] = {1'b0,layer_1_0[4847:4840]} - {1'b0, layer_0_0[4847:4840]};
      top_0[2] = {1'b0,layer_1_0[4855:4848]} - {1'b0, layer_0_0[4855:4848]};
      top_1[0] = {1'b0,layer_1_1[4839:4832]} - {1'b0, layer_0_1[4839:4832]};
      top_1[1] = {1'b0,layer_1_1[4847:4840]} - {1'b0, layer_0_1[4847:4840]};
      top_1[2] = {1'b0,layer_1_1[4855:4848]} - {1'b0, layer_0_1[4855:4848]};
      top_2[0] = {1'b0,layer_1_2[4839:4832]} - {1'b0, layer_0_2[4839:4832]};
      top_2[1] = {1'b0,layer_1_2[4847:4840]} - {1'b0, layer_0_2[4847:4840]};
      top_2[2] = {1'b0,layer_1_2[4855:4848]} - {1'b0, layer_0_2[4855:4848]};
      mid_0[0] = {1'b0,layer_2_0[4839:4832]} - {1'b0, layer_1_0[4839:4832]};
      mid_0[1] = {1'b0,layer_2_0[4847:4840]} - {1'b0, layer_1_0[4847:4840]};
      mid_0[2] = {1'b0,layer_2_0[4855:4848]} - {1'b0, layer_1_0[4855:4848]};
      mid_1[0] = {1'b0,layer_2_1[4839:4832]} - {1'b0, layer_1_1[4839:4832]};
      mid_1[1] = {1'b0,layer_2_1[4847:4840]} - {1'b0, layer_1_1[4847:4840]};
      mid_1[2] = {1'b0,layer_2_1[4855:4848]} - {1'b0, layer_1_1[4855:4848]};
      mid_2[0] = {1'b0,layer_2_2[4839:4832]} - {1'b0, layer_1_2[4839:4832]};
      mid_2[1] = {1'b0,layer_2_2[4847:4840]} - {1'b0, layer_1_2[4847:4840]};
      mid_2[2] = {1'b0,layer_2_2[4855:4848]} - {1'b0, layer_1_2[4855:4848]};
      btm_0[0] = {1'b0,layer_3_0[4839:4832]} - {1'b0, layer_2_0[4839:4832]};
      btm_0[1] = {1'b0,layer_3_0[4847:4840]} - {1'b0, layer_2_0[4847:4840]};
      btm_0[2] = {1'b0,layer_3_0[4855:4848]} - {1'b0, layer_2_0[4855:4848]};
      btm_1[0] = {1'b0,layer_3_1[4839:4832]} - {1'b0, layer_2_1[4839:4832]};
      btm_1[1] = {1'b0,layer_3_1[4847:4840]} - {1'b0, layer_2_1[4847:4840]};
      btm_1[2] = {1'b0,layer_3_1[4855:4848]} - {1'b0, layer_2_1[4855:4848]};
      btm_2[0] = {1'b0,layer_3_2[4839:4832]} - {1'b0, layer_2_2[4839:4832]};
      btm_2[1] = {1'b0,layer_3_2[4847:4840]} - {1'b0, layer_2_2[4847:4840]};
      btm_2[2] = {1'b0,layer_3_2[4855:4848]} - {1'b0, layer_2_2[4855:4848]};
    end
    'd606: begin
      top_0[0] = {1'b0,layer_1_0[4847:4840]} - {1'b0, layer_0_0[4847:4840]};
      top_0[1] = {1'b0,layer_1_0[4855:4848]} - {1'b0, layer_0_0[4855:4848]};
      top_0[2] = {1'b0,layer_1_0[4863:4856]} - {1'b0, layer_0_0[4863:4856]};
      top_1[0] = {1'b0,layer_1_1[4847:4840]} - {1'b0, layer_0_1[4847:4840]};
      top_1[1] = {1'b0,layer_1_1[4855:4848]} - {1'b0, layer_0_1[4855:4848]};
      top_1[2] = {1'b0,layer_1_1[4863:4856]} - {1'b0, layer_0_1[4863:4856]};
      top_2[0] = {1'b0,layer_1_2[4847:4840]} - {1'b0, layer_0_2[4847:4840]};
      top_2[1] = {1'b0,layer_1_2[4855:4848]} - {1'b0, layer_0_2[4855:4848]};
      top_2[2] = {1'b0,layer_1_2[4863:4856]} - {1'b0, layer_0_2[4863:4856]};
      mid_0[0] = {1'b0,layer_2_0[4847:4840]} - {1'b0, layer_1_0[4847:4840]};
      mid_0[1] = {1'b0,layer_2_0[4855:4848]} - {1'b0, layer_1_0[4855:4848]};
      mid_0[2] = {1'b0,layer_2_0[4863:4856]} - {1'b0, layer_1_0[4863:4856]};
      mid_1[0] = {1'b0,layer_2_1[4847:4840]} - {1'b0, layer_1_1[4847:4840]};
      mid_1[1] = {1'b0,layer_2_1[4855:4848]} - {1'b0, layer_1_1[4855:4848]};
      mid_1[2] = {1'b0,layer_2_1[4863:4856]} - {1'b0, layer_1_1[4863:4856]};
      mid_2[0] = {1'b0,layer_2_2[4847:4840]} - {1'b0, layer_1_2[4847:4840]};
      mid_2[1] = {1'b0,layer_2_2[4855:4848]} - {1'b0, layer_1_2[4855:4848]};
      mid_2[2] = {1'b0,layer_2_2[4863:4856]} - {1'b0, layer_1_2[4863:4856]};
      btm_0[0] = {1'b0,layer_3_0[4847:4840]} - {1'b0, layer_2_0[4847:4840]};
      btm_0[1] = {1'b0,layer_3_0[4855:4848]} - {1'b0, layer_2_0[4855:4848]};
      btm_0[2] = {1'b0,layer_3_0[4863:4856]} - {1'b0, layer_2_0[4863:4856]};
      btm_1[0] = {1'b0,layer_3_1[4847:4840]} - {1'b0, layer_2_1[4847:4840]};
      btm_1[1] = {1'b0,layer_3_1[4855:4848]} - {1'b0, layer_2_1[4855:4848]};
      btm_1[2] = {1'b0,layer_3_1[4863:4856]} - {1'b0, layer_2_1[4863:4856]};
      btm_2[0] = {1'b0,layer_3_2[4847:4840]} - {1'b0, layer_2_2[4847:4840]};
      btm_2[1] = {1'b0,layer_3_2[4855:4848]} - {1'b0, layer_2_2[4855:4848]};
      btm_2[2] = {1'b0,layer_3_2[4863:4856]} - {1'b0, layer_2_2[4863:4856]};
    end
    'd607: begin
      top_0[0] = {1'b0,layer_1_0[4855:4848]} - {1'b0, layer_0_0[4855:4848]};
      top_0[1] = {1'b0,layer_1_0[4863:4856]} - {1'b0, layer_0_0[4863:4856]};
      top_0[2] = {1'b0,layer_1_0[4871:4864]} - {1'b0, layer_0_0[4871:4864]};
      top_1[0] = {1'b0,layer_1_1[4855:4848]} - {1'b0, layer_0_1[4855:4848]};
      top_1[1] = {1'b0,layer_1_1[4863:4856]} - {1'b0, layer_0_1[4863:4856]};
      top_1[2] = {1'b0,layer_1_1[4871:4864]} - {1'b0, layer_0_1[4871:4864]};
      top_2[0] = {1'b0,layer_1_2[4855:4848]} - {1'b0, layer_0_2[4855:4848]};
      top_2[1] = {1'b0,layer_1_2[4863:4856]} - {1'b0, layer_0_2[4863:4856]};
      top_2[2] = {1'b0,layer_1_2[4871:4864]} - {1'b0, layer_0_2[4871:4864]};
      mid_0[0] = {1'b0,layer_2_0[4855:4848]} - {1'b0, layer_1_0[4855:4848]};
      mid_0[1] = {1'b0,layer_2_0[4863:4856]} - {1'b0, layer_1_0[4863:4856]};
      mid_0[2] = {1'b0,layer_2_0[4871:4864]} - {1'b0, layer_1_0[4871:4864]};
      mid_1[0] = {1'b0,layer_2_1[4855:4848]} - {1'b0, layer_1_1[4855:4848]};
      mid_1[1] = {1'b0,layer_2_1[4863:4856]} - {1'b0, layer_1_1[4863:4856]};
      mid_1[2] = {1'b0,layer_2_1[4871:4864]} - {1'b0, layer_1_1[4871:4864]};
      mid_2[0] = {1'b0,layer_2_2[4855:4848]} - {1'b0, layer_1_2[4855:4848]};
      mid_2[1] = {1'b0,layer_2_2[4863:4856]} - {1'b0, layer_1_2[4863:4856]};
      mid_2[2] = {1'b0,layer_2_2[4871:4864]} - {1'b0, layer_1_2[4871:4864]};
      btm_0[0] = {1'b0,layer_3_0[4855:4848]} - {1'b0, layer_2_0[4855:4848]};
      btm_0[1] = {1'b0,layer_3_0[4863:4856]} - {1'b0, layer_2_0[4863:4856]};
      btm_0[2] = {1'b0,layer_3_0[4871:4864]} - {1'b0, layer_2_0[4871:4864]};
      btm_1[0] = {1'b0,layer_3_1[4855:4848]} - {1'b0, layer_2_1[4855:4848]};
      btm_1[1] = {1'b0,layer_3_1[4863:4856]} - {1'b0, layer_2_1[4863:4856]};
      btm_1[2] = {1'b0,layer_3_1[4871:4864]} - {1'b0, layer_2_1[4871:4864]};
      btm_2[0] = {1'b0,layer_3_2[4855:4848]} - {1'b0, layer_2_2[4855:4848]};
      btm_2[1] = {1'b0,layer_3_2[4863:4856]} - {1'b0, layer_2_2[4863:4856]};
      btm_2[2] = {1'b0,layer_3_2[4871:4864]} - {1'b0, layer_2_2[4871:4864]};
    end
    'd608: begin
      top_0[0] = {1'b0,layer_1_0[4863:4856]} - {1'b0, layer_0_0[4863:4856]};
      top_0[1] = {1'b0,layer_1_0[4871:4864]} - {1'b0, layer_0_0[4871:4864]};
      top_0[2] = {1'b0,layer_1_0[4879:4872]} - {1'b0, layer_0_0[4879:4872]};
      top_1[0] = {1'b0,layer_1_1[4863:4856]} - {1'b0, layer_0_1[4863:4856]};
      top_1[1] = {1'b0,layer_1_1[4871:4864]} - {1'b0, layer_0_1[4871:4864]};
      top_1[2] = {1'b0,layer_1_1[4879:4872]} - {1'b0, layer_0_1[4879:4872]};
      top_2[0] = {1'b0,layer_1_2[4863:4856]} - {1'b0, layer_0_2[4863:4856]};
      top_2[1] = {1'b0,layer_1_2[4871:4864]} - {1'b0, layer_0_2[4871:4864]};
      top_2[2] = {1'b0,layer_1_2[4879:4872]} - {1'b0, layer_0_2[4879:4872]};
      mid_0[0] = {1'b0,layer_2_0[4863:4856]} - {1'b0, layer_1_0[4863:4856]};
      mid_0[1] = {1'b0,layer_2_0[4871:4864]} - {1'b0, layer_1_0[4871:4864]};
      mid_0[2] = {1'b0,layer_2_0[4879:4872]} - {1'b0, layer_1_0[4879:4872]};
      mid_1[0] = {1'b0,layer_2_1[4863:4856]} - {1'b0, layer_1_1[4863:4856]};
      mid_1[1] = {1'b0,layer_2_1[4871:4864]} - {1'b0, layer_1_1[4871:4864]};
      mid_1[2] = {1'b0,layer_2_1[4879:4872]} - {1'b0, layer_1_1[4879:4872]};
      mid_2[0] = {1'b0,layer_2_2[4863:4856]} - {1'b0, layer_1_2[4863:4856]};
      mid_2[1] = {1'b0,layer_2_2[4871:4864]} - {1'b0, layer_1_2[4871:4864]};
      mid_2[2] = {1'b0,layer_2_2[4879:4872]} - {1'b0, layer_1_2[4879:4872]};
      btm_0[0] = {1'b0,layer_3_0[4863:4856]} - {1'b0, layer_2_0[4863:4856]};
      btm_0[1] = {1'b0,layer_3_0[4871:4864]} - {1'b0, layer_2_0[4871:4864]};
      btm_0[2] = {1'b0,layer_3_0[4879:4872]} - {1'b0, layer_2_0[4879:4872]};
      btm_1[0] = {1'b0,layer_3_1[4863:4856]} - {1'b0, layer_2_1[4863:4856]};
      btm_1[1] = {1'b0,layer_3_1[4871:4864]} - {1'b0, layer_2_1[4871:4864]};
      btm_1[2] = {1'b0,layer_3_1[4879:4872]} - {1'b0, layer_2_1[4879:4872]};
      btm_2[0] = {1'b0,layer_3_2[4863:4856]} - {1'b0, layer_2_2[4863:4856]};
      btm_2[1] = {1'b0,layer_3_2[4871:4864]} - {1'b0, layer_2_2[4871:4864]};
      btm_2[2] = {1'b0,layer_3_2[4879:4872]} - {1'b0, layer_2_2[4879:4872]};
    end
    'd609: begin
      top_0[0] = {1'b0,layer_1_0[4871:4864]} - {1'b0, layer_0_0[4871:4864]};
      top_0[1] = {1'b0,layer_1_0[4879:4872]} - {1'b0, layer_0_0[4879:4872]};
      top_0[2] = {1'b0,layer_1_0[4887:4880]} - {1'b0, layer_0_0[4887:4880]};
      top_1[0] = {1'b0,layer_1_1[4871:4864]} - {1'b0, layer_0_1[4871:4864]};
      top_1[1] = {1'b0,layer_1_1[4879:4872]} - {1'b0, layer_0_1[4879:4872]};
      top_1[2] = {1'b0,layer_1_1[4887:4880]} - {1'b0, layer_0_1[4887:4880]};
      top_2[0] = {1'b0,layer_1_2[4871:4864]} - {1'b0, layer_0_2[4871:4864]};
      top_2[1] = {1'b0,layer_1_2[4879:4872]} - {1'b0, layer_0_2[4879:4872]};
      top_2[2] = {1'b0,layer_1_2[4887:4880]} - {1'b0, layer_0_2[4887:4880]};
      mid_0[0] = {1'b0,layer_2_0[4871:4864]} - {1'b0, layer_1_0[4871:4864]};
      mid_0[1] = {1'b0,layer_2_0[4879:4872]} - {1'b0, layer_1_0[4879:4872]};
      mid_0[2] = {1'b0,layer_2_0[4887:4880]} - {1'b0, layer_1_0[4887:4880]};
      mid_1[0] = {1'b0,layer_2_1[4871:4864]} - {1'b0, layer_1_1[4871:4864]};
      mid_1[1] = {1'b0,layer_2_1[4879:4872]} - {1'b0, layer_1_1[4879:4872]};
      mid_1[2] = {1'b0,layer_2_1[4887:4880]} - {1'b0, layer_1_1[4887:4880]};
      mid_2[0] = {1'b0,layer_2_2[4871:4864]} - {1'b0, layer_1_2[4871:4864]};
      mid_2[1] = {1'b0,layer_2_2[4879:4872]} - {1'b0, layer_1_2[4879:4872]};
      mid_2[2] = {1'b0,layer_2_2[4887:4880]} - {1'b0, layer_1_2[4887:4880]};
      btm_0[0] = {1'b0,layer_3_0[4871:4864]} - {1'b0, layer_2_0[4871:4864]};
      btm_0[1] = {1'b0,layer_3_0[4879:4872]} - {1'b0, layer_2_0[4879:4872]};
      btm_0[2] = {1'b0,layer_3_0[4887:4880]} - {1'b0, layer_2_0[4887:4880]};
      btm_1[0] = {1'b0,layer_3_1[4871:4864]} - {1'b0, layer_2_1[4871:4864]};
      btm_1[1] = {1'b0,layer_3_1[4879:4872]} - {1'b0, layer_2_1[4879:4872]};
      btm_1[2] = {1'b0,layer_3_1[4887:4880]} - {1'b0, layer_2_1[4887:4880]};
      btm_2[0] = {1'b0,layer_3_2[4871:4864]} - {1'b0, layer_2_2[4871:4864]};
      btm_2[1] = {1'b0,layer_3_2[4879:4872]} - {1'b0, layer_2_2[4879:4872]};
      btm_2[2] = {1'b0,layer_3_2[4887:4880]} - {1'b0, layer_2_2[4887:4880]};
    end
    'd610: begin
      top_0[0] = {1'b0,layer_1_0[4879:4872]} - {1'b0, layer_0_0[4879:4872]};
      top_0[1] = {1'b0,layer_1_0[4887:4880]} - {1'b0, layer_0_0[4887:4880]};
      top_0[2] = {1'b0,layer_1_0[4895:4888]} - {1'b0, layer_0_0[4895:4888]};
      top_1[0] = {1'b0,layer_1_1[4879:4872]} - {1'b0, layer_0_1[4879:4872]};
      top_1[1] = {1'b0,layer_1_1[4887:4880]} - {1'b0, layer_0_1[4887:4880]};
      top_1[2] = {1'b0,layer_1_1[4895:4888]} - {1'b0, layer_0_1[4895:4888]};
      top_2[0] = {1'b0,layer_1_2[4879:4872]} - {1'b0, layer_0_2[4879:4872]};
      top_2[1] = {1'b0,layer_1_2[4887:4880]} - {1'b0, layer_0_2[4887:4880]};
      top_2[2] = {1'b0,layer_1_2[4895:4888]} - {1'b0, layer_0_2[4895:4888]};
      mid_0[0] = {1'b0,layer_2_0[4879:4872]} - {1'b0, layer_1_0[4879:4872]};
      mid_0[1] = {1'b0,layer_2_0[4887:4880]} - {1'b0, layer_1_0[4887:4880]};
      mid_0[2] = {1'b0,layer_2_0[4895:4888]} - {1'b0, layer_1_0[4895:4888]};
      mid_1[0] = {1'b0,layer_2_1[4879:4872]} - {1'b0, layer_1_1[4879:4872]};
      mid_1[1] = {1'b0,layer_2_1[4887:4880]} - {1'b0, layer_1_1[4887:4880]};
      mid_1[2] = {1'b0,layer_2_1[4895:4888]} - {1'b0, layer_1_1[4895:4888]};
      mid_2[0] = {1'b0,layer_2_2[4879:4872]} - {1'b0, layer_1_2[4879:4872]};
      mid_2[1] = {1'b0,layer_2_2[4887:4880]} - {1'b0, layer_1_2[4887:4880]};
      mid_2[2] = {1'b0,layer_2_2[4895:4888]} - {1'b0, layer_1_2[4895:4888]};
      btm_0[0] = {1'b0,layer_3_0[4879:4872]} - {1'b0, layer_2_0[4879:4872]};
      btm_0[1] = {1'b0,layer_3_0[4887:4880]} - {1'b0, layer_2_0[4887:4880]};
      btm_0[2] = {1'b0,layer_3_0[4895:4888]} - {1'b0, layer_2_0[4895:4888]};
      btm_1[0] = {1'b0,layer_3_1[4879:4872]} - {1'b0, layer_2_1[4879:4872]};
      btm_1[1] = {1'b0,layer_3_1[4887:4880]} - {1'b0, layer_2_1[4887:4880]};
      btm_1[2] = {1'b0,layer_3_1[4895:4888]} - {1'b0, layer_2_1[4895:4888]};
      btm_2[0] = {1'b0,layer_3_2[4879:4872]} - {1'b0, layer_2_2[4879:4872]};
      btm_2[1] = {1'b0,layer_3_2[4887:4880]} - {1'b0, layer_2_2[4887:4880]};
      btm_2[2] = {1'b0,layer_3_2[4895:4888]} - {1'b0, layer_2_2[4895:4888]};
    end
    'd611: begin
      top_0[0] = {1'b0,layer_1_0[4887:4880]} - {1'b0, layer_0_0[4887:4880]};
      top_0[1] = {1'b0,layer_1_0[4895:4888]} - {1'b0, layer_0_0[4895:4888]};
      top_0[2] = {1'b0,layer_1_0[4903:4896]} - {1'b0, layer_0_0[4903:4896]};
      top_1[0] = {1'b0,layer_1_1[4887:4880]} - {1'b0, layer_0_1[4887:4880]};
      top_1[1] = {1'b0,layer_1_1[4895:4888]} - {1'b0, layer_0_1[4895:4888]};
      top_1[2] = {1'b0,layer_1_1[4903:4896]} - {1'b0, layer_0_1[4903:4896]};
      top_2[0] = {1'b0,layer_1_2[4887:4880]} - {1'b0, layer_0_2[4887:4880]};
      top_2[1] = {1'b0,layer_1_2[4895:4888]} - {1'b0, layer_0_2[4895:4888]};
      top_2[2] = {1'b0,layer_1_2[4903:4896]} - {1'b0, layer_0_2[4903:4896]};
      mid_0[0] = {1'b0,layer_2_0[4887:4880]} - {1'b0, layer_1_0[4887:4880]};
      mid_0[1] = {1'b0,layer_2_0[4895:4888]} - {1'b0, layer_1_0[4895:4888]};
      mid_0[2] = {1'b0,layer_2_0[4903:4896]} - {1'b0, layer_1_0[4903:4896]};
      mid_1[0] = {1'b0,layer_2_1[4887:4880]} - {1'b0, layer_1_1[4887:4880]};
      mid_1[1] = {1'b0,layer_2_1[4895:4888]} - {1'b0, layer_1_1[4895:4888]};
      mid_1[2] = {1'b0,layer_2_1[4903:4896]} - {1'b0, layer_1_1[4903:4896]};
      mid_2[0] = {1'b0,layer_2_2[4887:4880]} - {1'b0, layer_1_2[4887:4880]};
      mid_2[1] = {1'b0,layer_2_2[4895:4888]} - {1'b0, layer_1_2[4895:4888]};
      mid_2[2] = {1'b0,layer_2_2[4903:4896]} - {1'b0, layer_1_2[4903:4896]};
      btm_0[0] = {1'b0,layer_3_0[4887:4880]} - {1'b0, layer_2_0[4887:4880]};
      btm_0[1] = {1'b0,layer_3_0[4895:4888]} - {1'b0, layer_2_0[4895:4888]};
      btm_0[2] = {1'b0,layer_3_0[4903:4896]} - {1'b0, layer_2_0[4903:4896]};
      btm_1[0] = {1'b0,layer_3_1[4887:4880]} - {1'b0, layer_2_1[4887:4880]};
      btm_1[1] = {1'b0,layer_3_1[4895:4888]} - {1'b0, layer_2_1[4895:4888]};
      btm_1[2] = {1'b0,layer_3_1[4903:4896]} - {1'b0, layer_2_1[4903:4896]};
      btm_2[0] = {1'b0,layer_3_2[4887:4880]} - {1'b0, layer_2_2[4887:4880]};
      btm_2[1] = {1'b0,layer_3_2[4895:4888]} - {1'b0, layer_2_2[4895:4888]};
      btm_2[2] = {1'b0,layer_3_2[4903:4896]} - {1'b0, layer_2_2[4903:4896]};
    end
    'd612: begin
      top_0[0] = {1'b0,layer_1_0[4895:4888]} - {1'b0, layer_0_0[4895:4888]};
      top_0[1] = {1'b0,layer_1_0[4903:4896]} - {1'b0, layer_0_0[4903:4896]};
      top_0[2] = {1'b0,layer_1_0[4911:4904]} - {1'b0, layer_0_0[4911:4904]};
      top_1[0] = {1'b0,layer_1_1[4895:4888]} - {1'b0, layer_0_1[4895:4888]};
      top_1[1] = {1'b0,layer_1_1[4903:4896]} - {1'b0, layer_0_1[4903:4896]};
      top_1[2] = {1'b0,layer_1_1[4911:4904]} - {1'b0, layer_0_1[4911:4904]};
      top_2[0] = {1'b0,layer_1_2[4895:4888]} - {1'b0, layer_0_2[4895:4888]};
      top_2[1] = {1'b0,layer_1_2[4903:4896]} - {1'b0, layer_0_2[4903:4896]};
      top_2[2] = {1'b0,layer_1_2[4911:4904]} - {1'b0, layer_0_2[4911:4904]};
      mid_0[0] = {1'b0,layer_2_0[4895:4888]} - {1'b0, layer_1_0[4895:4888]};
      mid_0[1] = {1'b0,layer_2_0[4903:4896]} - {1'b0, layer_1_0[4903:4896]};
      mid_0[2] = {1'b0,layer_2_0[4911:4904]} - {1'b0, layer_1_0[4911:4904]};
      mid_1[0] = {1'b0,layer_2_1[4895:4888]} - {1'b0, layer_1_1[4895:4888]};
      mid_1[1] = {1'b0,layer_2_1[4903:4896]} - {1'b0, layer_1_1[4903:4896]};
      mid_1[2] = {1'b0,layer_2_1[4911:4904]} - {1'b0, layer_1_1[4911:4904]};
      mid_2[0] = {1'b0,layer_2_2[4895:4888]} - {1'b0, layer_1_2[4895:4888]};
      mid_2[1] = {1'b0,layer_2_2[4903:4896]} - {1'b0, layer_1_2[4903:4896]};
      mid_2[2] = {1'b0,layer_2_2[4911:4904]} - {1'b0, layer_1_2[4911:4904]};
      btm_0[0] = {1'b0,layer_3_0[4895:4888]} - {1'b0, layer_2_0[4895:4888]};
      btm_0[1] = {1'b0,layer_3_0[4903:4896]} - {1'b0, layer_2_0[4903:4896]};
      btm_0[2] = {1'b0,layer_3_0[4911:4904]} - {1'b0, layer_2_0[4911:4904]};
      btm_1[0] = {1'b0,layer_3_1[4895:4888]} - {1'b0, layer_2_1[4895:4888]};
      btm_1[1] = {1'b0,layer_3_1[4903:4896]} - {1'b0, layer_2_1[4903:4896]};
      btm_1[2] = {1'b0,layer_3_1[4911:4904]} - {1'b0, layer_2_1[4911:4904]};
      btm_2[0] = {1'b0,layer_3_2[4895:4888]} - {1'b0, layer_2_2[4895:4888]};
      btm_2[1] = {1'b0,layer_3_2[4903:4896]} - {1'b0, layer_2_2[4903:4896]};
      btm_2[2] = {1'b0,layer_3_2[4911:4904]} - {1'b0, layer_2_2[4911:4904]};
    end
    'd613: begin
      top_0[0] = {1'b0,layer_1_0[4903:4896]} - {1'b0, layer_0_0[4903:4896]};
      top_0[1] = {1'b0,layer_1_0[4911:4904]} - {1'b0, layer_0_0[4911:4904]};
      top_0[2] = {1'b0,layer_1_0[4919:4912]} - {1'b0, layer_0_0[4919:4912]};
      top_1[0] = {1'b0,layer_1_1[4903:4896]} - {1'b0, layer_0_1[4903:4896]};
      top_1[1] = {1'b0,layer_1_1[4911:4904]} - {1'b0, layer_0_1[4911:4904]};
      top_1[2] = {1'b0,layer_1_1[4919:4912]} - {1'b0, layer_0_1[4919:4912]};
      top_2[0] = {1'b0,layer_1_2[4903:4896]} - {1'b0, layer_0_2[4903:4896]};
      top_2[1] = {1'b0,layer_1_2[4911:4904]} - {1'b0, layer_0_2[4911:4904]};
      top_2[2] = {1'b0,layer_1_2[4919:4912]} - {1'b0, layer_0_2[4919:4912]};
      mid_0[0] = {1'b0,layer_2_0[4903:4896]} - {1'b0, layer_1_0[4903:4896]};
      mid_0[1] = {1'b0,layer_2_0[4911:4904]} - {1'b0, layer_1_0[4911:4904]};
      mid_0[2] = {1'b0,layer_2_0[4919:4912]} - {1'b0, layer_1_0[4919:4912]};
      mid_1[0] = {1'b0,layer_2_1[4903:4896]} - {1'b0, layer_1_1[4903:4896]};
      mid_1[1] = {1'b0,layer_2_1[4911:4904]} - {1'b0, layer_1_1[4911:4904]};
      mid_1[2] = {1'b0,layer_2_1[4919:4912]} - {1'b0, layer_1_1[4919:4912]};
      mid_2[0] = {1'b0,layer_2_2[4903:4896]} - {1'b0, layer_1_2[4903:4896]};
      mid_2[1] = {1'b0,layer_2_2[4911:4904]} - {1'b0, layer_1_2[4911:4904]};
      mid_2[2] = {1'b0,layer_2_2[4919:4912]} - {1'b0, layer_1_2[4919:4912]};
      btm_0[0] = {1'b0,layer_3_0[4903:4896]} - {1'b0, layer_2_0[4903:4896]};
      btm_0[1] = {1'b0,layer_3_0[4911:4904]} - {1'b0, layer_2_0[4911:4904]};
      btm_0[2] = {1'b0,layer_3_0[4919:4912]} - {1'b0, layer_2_0[4919:4912]};
      btm_1[0] = {1'b0,layer_3_1[4903:4896]} - {1'b0, layer_2_1[4903:4896]};
      btm_1[1] = {1'b0,layer_3_1[4911:4904]} - {1'b0, layer_2_1[4911:4904]};
      btm_1[2] = {1'b0,layer_3_1[4919:4912]} - {1'b0, layer_2_1[4919:4912]};
      btm_2[0] = {1'b0,layer_3_2[4903:4896]} - {1'b0, layer_2_2[4903:4896]};
      btm_2[1] = {1'b0,layer_3_2[4911:4904]} - {1'b0, layer_2_2[4911:4904]};
      btm_2[2] = {1'b0,layer_3_2[4919:4912]} - {1'b0, layer_2_2[4919:4912]};
    end
    'd614: begin
      top_0[0] = {1'b0,layer_1_0[4911:4904]} - {1'b0, layer_0_0[4911:4904]};
      top_0[1] = {1'b0,layer_1_0[4919:4912]} - {1'b0, layer_0_0[4919:4912]};
      top_0[2] = {1'b0,layer_1_0[4927:4920]} - {1'b0, layer_0_0[4927:4920]};
      top_1[0] = {1'b0,layer_1_1[4911:4904]} - {1'b0, layer_0_1[4911:4904]};
      top_1[1] = {1'b0,layer_1_1[4919:4912]} - {1'b0, layer_0_1[4919:4912]};
      top_1[2] = {1'b0,layer_1_1[4927:4920]} - {1'b0, layer_0_1[4927:4920]};
      top_2[0] = {1'b0,layer_1_2[4911:4904]} - {1'b0, layer_0_2[4911:4904]};
      top_2[1] = {1'b0,layer_1_2[4919:4912]} - {1'b0, layer_0_2[4919:4912]};
      top_2[2] = {1'b0,layer_1_2[4927:4920]} - {1'b0, layer_0_2[4927:4920]};
      mid_0[0] = {1'b0,layer_2_0[4911:4904]} - {1'b0, layer_1_0[4911:4904]};
      mid_0[1] = {1'b0,layer_2_0[4919:4912]} - {1'b0, layer_1_0[4919:4912]};
      mid_0[2] = {1'b0,layer_2_0[4927:4920]} - {1'b0, layer_1_0[4927:4920]};
      mid_1[0] = {1'b0,layer_2_1[4911:4904]} - {1'b0, layer_1_1[4911:4904]};
      mid_1[1] = {1'b0,layer_2_1[4919:4912]} - {1'b0, layer_1_1[4919:4912]};
      mid_1[2] = {1'b0,layer_2_1[4927:4920]} - {1'b0, layer_1_1[4927:4920]};
      mid_2[0] = {1'b0,layer_2_2[4911:4904]} - {1'b0, layer_1_2[4911:4904]};
      mid_2[1] = {1'b0,layer_2_2[4919:4912]} - {1'b0, layer_1_2[4919:4912]};
      mid_2[2] = {1'b0,layer_2_2[4927:4920]} - {1'b0, layer_1_2[4927:4920]};
      btm_0[0] = {1'b0,layer_3_0[4911:4904]} - {1'b0, layer_2_0[4911:4904]};
      btm_0[1] = {1'b0,layer_3_0[4919:4912]} - {1'b0, layer_2_0[4919:4912]};
      btm_0[2] = {1'b0,layer_3_0[4927:4920]} - {1'b0, layer_2_0[4927:4920]};
      btm_1[0] = {1'b0,layer_3_1[4911:4904]} - {1'b0, layer_2_1[4911:4904]};
      btm_1[1] = {1'b0,layer_3_1[4919:4912]} - {1'b0, layer_2_1[4919:4912]};
      btm_1[2] = {1'b0,layer_3_1[4927:4920]} - {1'b0, layer_2_1[4927:4920]};
      btm_2[0] = {1'b0,layer_3_2[4911:4904]} - {1'b0, layer_2_2[4911:4904]};
      btm_2[1] = {1'b0,layer_3_2[4919:4912]} - {1'b0, layer_2_2[4919:4912]};
      btm_2[2] = {1'b0,layer_3_2[4927:4920]} - {1'b0, layer_2_2[4927:4920]};
    end
    'd615: begin
      top_0[0] = {1'b0,layer_1_0[4919:4912]} - {1'b0, layer_0_0[4919:4912]};
      top_0[1] = {1'b0,layer_1_0[4927:4920]} - {1'b0, layer_0_0[4927:4920]};
      top_0[2] = {1'b0,layer_1_0[4935:4928]} - {1'b0, layer_0_0[4935:4928]};
      top_1[0] = {1'b0,layer_1_1[4919:4912]} - {1'b0, layer_0_1[4919:4912]};
      top_1[1] = {1'b0,layer_1_1[4927:4920]} - {1'b0, layer_0_1[4927:4920]};
      top_1[2] = {1'b0,layer_1_1[4935:4928]} - {1'b0, layer_0_1[4935:4928]};
      top_2[0] = {1'b0,layer_1_2[4919:4912]} - {1'b0, layer_0_2[4919:4912]};
      top_2[1] = {1'b0,layer_1_2[4927:4920]} - {1'b0, layer_0_2[4927:4920]};
      top_2[2] = {1'b0,layer_1_2[4935:4928]} - {1'b0, layer_0_2[4935:4928]};
      mid_0[0] = {1'b0,layer_2_0[4919:4912]} - {1'b0, layer_1_0[4919:4912]};
      mid_0[1] = {1'b0,layer_2_0[4927:4920]} - {1'b0, layer_1_0[4927:4920]};
      mid_0[2] = {1'b0,layer_2_0[4935:4928]} - {1'b0, layer_1_0[4935:4928]};
      mid_1[0] = {1'b0,layer_2_1[4919:4912]} - {1'b0, layer_1_1[4919:4912]};
      mid_1[1] = {1'b0,layer_2_1[4927:4920]} - {1'b0, layer_1_1[4927:4920]};
      mid_1[2] = {1'b0,layer_2_1[4935:4928]} - {1'b0, layer_1_1[4935:4928]};
      mid_2[0] = {1'b0,layer_2_2[4919:4912]} - {1'b0, layer_1_2[4919:4912]};
      mid_2[1] = {1'b0,layer_2_2[4927:4920]} - {1'b0, layer_1_2[4927:4920]};
      mid_2[2] = {1'b0,layer_2_2[4935:4928]} - {1'b0, layer_1_2[4935:4928]};
      btm_0[0] = {1'b0,layer_3_0[4919:4912]} - {1'b0, layer_2_0[4919:4912]};
      btm_0[1] = {1'b0,layer_3_0[4927:4920]} - {1'b0, layer_2_0[4927:4920]};
      btm_0[2] = {1'b0,layer_3_0[4935:4928]} - {1'b0, layer_2_0[4935:4928]};
      btm_1[0] = {1'b0,layer_3_1[4919:4912]} - {1'b0, layer_2_1[4919:4912]};
      btm_1[1] = {1'b0,layer_3_1[4927:4920]} - {1'b0, layer_2_1[4927:4920]};
      btm_1[2] = {1'b0,layer_3_1[4935:4928]} - {1'b0, layer_2_1[4935:4928]};
      btm_2[0] = {1'b0,layer_3_2[4919:4912]} - {1'b0, layer_2_2[4919:4912]};
      btm_2[1] = {1'b0,layer_3_2[4927:4920]} - {1'b0, layer_2_2[4927:4920]};
      btm_2[2] = {1'b0,layer_3_2[4935:4928]} - {1'b0, layer_2_2[4935:4928]};
    end
    'd616: begin
      top_0[0] = {1'b0,layer_1_0[4927:4920]} - {1'b0, layer_0_0[4927:4920]};
      top_0[1] = {1'b0,layer_1_0[4935:4928]} - {1'b0, layer_0_0[4935:4928]};
      top_0[2] = {1'b0,layer_1_0[4943:4936]} - {1'b0, layer_0_0[4943:4936]};
      top_1[0] = {1'b0,layer_1_1[4927:4920]} - {1'b0, layer_0_1[4927:4920]};
      top_1[1] = {1'b0,layer_1_1[4935:4928]} - {1'b0, layer_0_1[4935:4928]};
      top_1[2] = {1'b0,layer_1_1[4943:4936]} - {1'b0, layer_0_1[4943:4936]};
      top_2[0] = {1'b0,layer_1_2[4927:4920]} - {1'b0, layer_0_2[4927:4920]};
      top_2[1] = {1'b0,layer_1_2[4935:4928]} - {1'b0, layer_0_2[4935:4928]};
      top_2[2] = {1'b0,layer_1_2[4943:4936]} - {1'b0, layer_0_2[4943:4936]};
      mid_0[0] = {1'b0,layer_2_0[4927:4920]} - {1'b0, layer_1_0[4927:4920]};
      mid_0[1] = {1'b0,layer_2_0[4935:4928]} - {1'b0, layer_1_0[4935:4928]};
      mid_0[2] = {1'b0,layer_2_0[4943:4936]} - {1'b0, layer_1_0[4943:4936]};
      mid_1[0] = {1'b0,layer_2_1[4927:4920]} - {1'b0, layer_1_1[4927:4920]};
      mid_1[1] = {1'b0,layer_2_1[4935:4928]} - {1'b0, layer_1_1[4935:4928]};
      mid_1[2] = {1'b0,layer_2_1[4943:4936]} - {1'b0, layer_1_1[4943:4936]};
      mid_2[0] = {1'b0,layer_2_2[4927:4920]} - {1'b0, layer_1_2[4927:4920]};
      mid_2[1] = {1'b0,layer_2_2[4935:4928]} - {1'b0, layer_1_2[4935:4928]};
      mid_2[2] = {1'b0,layer_2_2[4943:4936]} - {1'b0, layer_1_2[4943:4936]};
      btm_0[0] = {1'b0,layer_3_0[4927:4920]} - {1'b0, layer_2_0[4927:4920]};
      btm_0[1] = {1'b0,layer_3_0[4935:4928]} - {1'b0, layer_2_0[4935:4928]};
      btm_0[2] = {1'b0,layer_3_0[4943:4936]} - {1'b0, layer_2_0[4943:4936]};
      btm_1[0] = {1'b0,layer_3_1[4927:4920]} - {1'b0, layer_2_1[4927:4920]};
      btm_1[1] = {1'b0,layer_3_1[4935:4928]} - {1'b0, layer_2_1[4935:4928]};
      btm_1[2] = {1'b0,layer_3_1[4943:4936]} - {1'b0, layer_2_1[4943:4936]};
      btm_2[0] = {1'b0,layer_3_2[4927:4920]} - {1'b0, layer_2_2[4927:4920]};
      btm_2[1] = {1'b0,layer_3_2[4935:4928]} - {1'b0, layer_2_2[4935:4928]};
      btm_2[2] = {1'b0,layer_3_2[4943:4936]} - {1'b0, layer_2_2[4943:4936]};
    end
    'd617: begin
      top_0[0] = {1'b0,layer_1_0[4935:4928]} - {1'b0, layer_0_0[4935:4928]};
      top_0[1] = {1'b0,layer_1_0[4943:4936]} - {1'b0, layer_0_0[4943:4936]};
      top_0[2] = {1'b0,layer_1_0[4951:4944]} - {1'b0, layer_0_0[4951:4944]};
      top_1[0] = {1'b0,layer_1_1[4935:4928]} - {1'b0, layer_0_1[4935:4928]};
      top_1[1] = {1'b0,layer_1_1[4943:4936]} - {1'b0, layer_0_1[4943:4936]};
      top_1[2] = {1'b0,layer_1_1[4951:4944]} - {1'b0, layer_0_1[4951:4944]};
      top_2[0] = {1'b0,layer_1_2[4935:4928]} - {1'b0, layer_0_2[4935:4928]};
      top_2[1] = {1'b0,layer_1_2[4943:4936]} - {1'b0, layer_0_2[4943:4936]};
      top_2[2] = {1'b0,layer_1_2[4951:4944]} - {1'b0, layer_0_2[4951:4944]};
      mid_0[0] = {1'b0,layer_2_0[4935:4928]} - {1'b0, layer_1_0[4935:4928]};
      mid_0[1] = {1'b0,layer_2_0[4943:4936]} - {1'b0, layer_1_0[4943:4936]};
      mid_0[2] = {1'b0,layer_2_0[4951:4944]} - {1'b0, layer_1_0[4951:4944]};
      mid_1[0] = {1'b0,layer_2_1[4935:4928]} - {1'b0, layer_1_1[4935:4928]};
      mid_1[1] = {1'b0,layer_2_1[4943:4936]} - {1'b0, layer_1_1[4943:4936]};
      mid_1[2] = {1'b0,layer_2_1[4951:4944]} - {1'b0, layer_1_1[4951:4944]};
      mid_2[0] = {1'b0,layer_2_2[4935:4928]} - {1'b0, layer_1_2[4935:4928]};
      mid_2[1] = {1'b0,layer_2_2[4943:4936]} - {1'b0, layer_1_2[4943:4936]};
      mid_2[2] = {1'b0,layer_2_2[4951:4944]} - {1'b0, layer_1_2[4951:4944]};
      btm_0[0] = {1'b0,layer_3_0[4935:4928]} - {1'b0, layer_2_0[4935:4928]};
      btm_0[1] = {1'b0,layer_3_0[4943:4936]} - {1'b0, layer_2_0[4943:4936]};
      btm_0[2] = {1'b0,layer_3_0[4951:4944]} - {1'b0, layer_2_0[4951:4944]};
      btm_1[0] = {1'b0,layer_3_1[4935:4928]} - {1'b0, layer_2_1[4935:4928]};
      btm_1[1] = {1'b0,layer_3_1[4943:4936]} - {1'b0, layer_2_1[4943:4936]};
      btm_1[2] = {1'b0,layer_3_1[4951:4944]} - {1'b0, layer_2_1[4951:4944]};
      btm_2[0] = {1'b0,layer_3_2[4935:4928]} - {1'b0, layer_2_2[4935:4928]};
      btm_2[1] = {1'b0,layer_3_2[4943:4936]} - {1'b0, layer_2_2[4943:4936]};
      btm_2[2] = {1'b0,layer_3_2[4951:4944]} - {1'b0, layer_2_2[4951:4944]};
    end
    'd618: begin
      top_0[0] = {1'b0,layer_1_0[4943:4936]} - {1'b0, layer_0_0[4943:4936]};
      top_0[1] = {1'b0,layer_1_0[4951:4944]} - {1'b0, layer_0_0[4951:4944]};
      top_0[2] = {1'b0,layer_1_0[4959:4952]} - {1'b0, layer_0_0[4959:4952]};
      top_1[0] = {1'b0,layer_1_1[4943:4936]} - {1'b0, layer_0_1[4943:4936]};
      top_1[1] = {1'b0,layer_1_1[4951:4944]} - {1'b0, layer_0_1[4951:4944]};
      top_1[2] = {1'b0,layer_1_1[4959:4952]} - {1'b0, layer_0_1[4959:4952]};
      top_2[0] = {1'b0,layer_1_2[4943:4936]} - {1'b0, layer_0_2[4943:4936]};
      top_2[1] = {1'b0,layer_1_2[4951:4944]} - {1'b0, layer_0_2[4951:4944]};
      top_2[2] = {1'b0,layer_1_2[4959:4952]} - {1'b0, layer_0_2[4959:4952]};
      mid_0[0] = {1'b0,layer_2_0[4943:4936]} - {1'b0, layer_1_0[4943:4936]};
      mid_0[1] = {1'b0,layer_2_0[4951:4944]} - {1'b0, layer_1_0[4951:4944]};
      mid_0[2] = {1'b0,layer_2_0[4959:4952]} - {1'b0, layer_1_0[4959:4952]};
      mid_1[0] = {1'b0,layer_2_1[4943:4936]} - {1'b0, layer_1_1[4943:4936]};
      mid_1[1] = {1'b0,layer_2_1[4951:4944]} - {1'b0, layer_1_1[4951:4944]};
      mid_1[2] = {1'b0,layer_2_1[4959:4952]} - {1'b0, layer_1_1[4959:4952]};
      mid_2[0] = {1'b0,layer_2_2[4943:4936]} - {1'b0, layer_1_2[4943:4936]};
      mid_2[1] = {1'b0,layer_2_2[4951:4944]} - {1'b0, layer_1_2[4951:4944]};
      mid_2[2] = {1'b0,layer_2_2[4959:4952]} - {1'b0, layer_1_2[4959:4952]};
      btm_0[0] = {1'b0,layer_3_0[4943:4936]} - {1'b0, layer_2_0[4943:4936]};
      btm_0[1] = {1'b0,layer_3_0[4951:4944]} - {1'b0, layer_2_0[4951:4944]};
      btm_0[2] = {1'b0,layer_3_0[4959:4952]} - {1'b0, layer_2_0[4959:4952]};
      btm_1[0] = {1'b0,layer_3_1[4943:4936]} - {1'b0, layer_2_1[4943:4936]};
      btm_1[1] = {1'b0,layer_3_1[4951:4944]} - {1'b0, layer_2_1[4951:4944]};
      btm_1[2] = {1'b0,layer_3_1[4959:4952]} - {1'b0, layer_2_1[4959:4952]};
      btm_2[0] = {1'b0,layer_3_2[4943:4936]} - {1'b0, layer_2_2[4943:4936]};
      btm_2[1] = {1'b0,layer_3_2[4951:4944]} - {1'b0, layer_2_2[4951:4944]};
      btm_2[2] = {1'b0,layer_3_2[4959:4952]} - {1'b0, layer_2_2[4959:4952]};
    end
    'd619: begin
      top_0[0] = {1'b0,layer_1_0[4951:4944]} - {1'b0, layer_0_0[4951:4944]};
      top_0[1] = {1'b0,layer_1_0[4959:4952]} - {1'b0, layer_0_0[4959:4952]};
      top_0[2] = {1'b0,layer_1_0[4967:4960]} - {1'b0, layer_0_0[4967:4960]};
      top_1[0] = {1'b0,layer_1_1[4951:4944]} - {1'b0, layer_0_1[4951:4944]};
      top_1[1] = {1'b0,layer_1_1[4959:4952]} - {1'b0, layer_0_1[4959:4952]};
      top_1[2] = {1'b0,layer_1_1[4967:4960]} - {1'b0, layer_0_1[4967:4960]};
      top_2[0] = {1'b0,layer_1_2[4951:4944]} - {1'b0, layer_0_2[4951:4944]};
      top_2[1] = {1'b0,layer_1_2[4959:4952]} - {1'b0, layer_0_2[4959:4952]};
      top_2[2] = {1'b0,layer_1_2[4967:4960]} - {1'b0, layer_0_2[4967:4960]};
      mid_0[0] = {1'b0,layer_2_0[4951:4944]} - {1'b0, layer_1_0[4951:4944]};
      mid_0[1] = {1'b0,layer_2_0[4959:4952]} - {1'b0, layer_1_0[4959:4952]};
      mid_0[2] = {1'b0,layer_2_0[4967:4960]} - {1'b0, layer_1_0[4967:4960]};
      mid_1[0] = {1'b0,layer_2_1[4951:4944]} - {1'b0, layer_1_1[4951:4944]};
      mid_1[1] = {1'b0,layer_2_1[4959:4952]} - {1'b0, layer_1_1[4959:4952]};
      mid_1[2] = {1'b0,layer_2_1[4967:4960]} - {1'b0, layer_1_1[4967:4960]};
      mid_2[0] = {1'b0,layer_2_2[4951:4944]} - {1'b0, layer_1_2[4951:4944]};
      mid_2[1] = {1'b0,layer_2_2[4959:4952]} - {1'b0, layer_1_2[4959:4952]};
      mid_2[2] = {1'b0,layer_2_2[4967:4960]} - {1'b0, layer_1_2[4967:4960]};
      btm_0[0] = {1'b0,layer_3_0[4951:4944]} - {1'b0, layer_2_0[4951:4944]};
      btm_0[1] = {1'b0,layer_3_0[4959:4952]} - {1'b0, layer_2_0[4959:4952]};
      btm_0[2] = {1'b0,layer_3_0[4967:4960]} - {1'b0, layer_2_0[4967:4960]};
      btm_1[0] = {1'b0,layer_3_1[4951:4944]} - {1'b0, layer_2_1[4951:4944]};
      btm_1[1] = {1'b0,layer_3_1[4959:4952]} - {1'b0, layer_2_1[4959:4952]};
      btm_1[2] = {1'b0,layer_3_1[4967:4960]} - {1'b0, layer_2_1[4967:4960]};
      btm_2[0] = {1'b0,layer_3_2[4951:4944]} - {1'b0, layer_2_2[4951:4944]};
      btm_2[1] = {1'b0,layer_3_2[4959:4952]} - {1'b0, layer_2_2[4959:4952]};
      btm_2[2] = {1'b0,layer_3_2[4967:4960]} - {1'b0, layer_2_2[4967:4960]};
    end
    'd620: begin
      top_0[0] = {1'b0,layer_1_0[4959:4952]} - {1'b0, layer_0_0[4959:4952]};
      top_0[1] = {1'b0,layer_1_0[4967:4960]} - {1'b0, layer_0_0[4967:4960]};
      top_0[2] = {1'b0,layer_1_0[4975:4968]} - {1'b0, layer_0_0[4975:4968]};
      top_1[0] = {1'b0,layer_1_1[4959:4952]} - {1'b0, layer_0_1[4959:4952]};
      top_1[1] = {1'b0,layer_1_1[4967:4960]} - {1'b0, layer_0_1[4967:4960]};
      top_1[2] = {1'b0,layer_1_1[4975:4968]} - {1'b0, layer_0_1[4975:4968]};
      top_2[0] = {1'b0,layer_1_2[4959:4952]} - {1'b0, layer_0_2[4959:4952]};
      top_2[1] = {1'b0,layer_1_2[4967:4960]} - {1'b0, layer_0_2[4967:4960]};
      top_2[2] = {1'b0,layer_1_2[4975:4968]} - {1'b0, layer_0_2[4975:4968]};
      mid_0[0] = {1'b0,layer_2_0[4959:4952]} - {1'b0, layer_1_0[4959:4952]};
      mid_0[1] = {1'b0,layer_2_0[4967:4960]} - {1'b0, layer_1_0[4967:4960]};
      mid_0[2] = {1'b0,layer_2_0[4975:4968]} - {1'b0, layer_1_0[4975:4968]};
      mid_1[0] = {1'b0,layer_2_1[4959:4952]} - {1'b0, layer_1_1[4959:4952]};
      mid_1[1] = {1'b0,layer_2_1[4967:4960]} - {1'b0, layer_1_1[4967:4960]};
      mid_1[2] = {1'b0,layer_2_1[4975:4968]} - {1'b0, layer_1_1[4975:4968]};
      mid_2[0] = {1'b0,layer_2_2[4959:4952]} - {1'b0, layer_1_2[4959:4952]};
      mid_2[1] = {1'b0,layer_2_2[4967:4960]} - {1'b0, layer_1_2[4967:4960]};
      mid_2[2] = {1'b0,layer_2_2[4975:4968]} - {1'b0, layer_1_2[4975:4968]};
      btm_0[0] = {1'b0,layer_3_0[4959:4952]} - {1'b0, layer_2_0[4959:4952]};
      btm_0[1] = {1'b0,layer_3_0[4967:4960]} - {1'b0, layer_2_0[4967:4960]};
      btm_0[2] = {1'b0,layer_3_0[4975:4968]} - {1'b0, layer_2_0[4975:4968]};
      btm_1[0] = {1'b0,layer_3_1[4959:4952]} - {1'b0, layer_2_1[4959:4952]};
      btm_1[1] = {1'b0,layer_3_1[4967:4960]} - {1'b0, layer_2_1[4967:4960]};
      btm_1[2] = {1'b0,layer_3_1[4975:4968]} - {1'b0, layer_2_1[4975:4968]};
      btm_2[0] = {1'b0,layer_3_2[4959:4952]} - {1'b0, layer_2_2[4959:4952]};
      btm_2[1] = {1'b0,layer_3_2[4967:4960]} - {1'b0, layer_2_2[4967:4960]};
      btm_2[2] = {1'b0,layer_3_2[4975:4968]} - {1'b0, layer_2_2[4975:4968]};
    end
    'd621: begin
      top_0[0] = {1'b0,layer_1_0[4967:4960]} - {1'b0, layer_0_0[4967:4960]};
      top_0[1] = {1'b0,layer_1_0[4975:4968]} - {1'b0, layer_0_0[4975:4968]};
      top_0[2] = {1'b0,layer_1_0[4983:4976]} - {1'b0, layer_0_0[4983:4976]};
      top_1[0] = {1'b0,layer_1_1[4967:4960]} - {1'b0, layer_0_1[4967:4960]};
      top_1[1] = {1'b0,layer_1_1[4975:4968]} - {1'b0, layer_0_1[4975:4968]};
      top_1[2] = {1'b0,layer_1_1[4983:4976]} - {1'b0, layer_0_1[4983:4976]};
      top_2[0] = {1'b0,layer_1_2[4967:4960]} - {1'b0, layer_0_2[4967:4960]};
      top_2[1] = {1'b0,layer_1_2[4975:4968]} - {1'b0, layer_0_2[4975:4968]};
      top_2[2] = {1'b0,layer_1_2[4983:4976]} - {1'b0, layer_0_2[4983:4976]};
      mid_0[0] = {1'b0,layer_2_0[4967:4960]} - {1'b0, layer_1_0[4967:4960]};
      mid_0[1] = {1'b0,layer_2_0[4975:4968]} - {1'b0, layer_1_0[4975:4968]};
      mid_0[2] = {1'b0,layer_2_0[4983:4976]} - {1'b0, layer_1_0[4983:4976]};
      mid_1[0] = {1'b0,layer_2_1[4967:4960]} - {1'b0, layer_1_1[4967:4960]};
      mid_1[1] = {1'b0,layer_2_1[4975:4968]} - {1'b0, layer_1_1[4975:4968]};
      mid_1[2] = {1'b0,layer_2_1[4983:4976]} - {1'b0, layer_1_1[4983:4976]};
      mid_2[0] = {1'b0,layer_2_2[4967:4960]} - {1'b0, layer_1_2[4967:4960]};
      mid_2[1] = {1'b0,layer_2_2[4975:4968]} - {1'b0, layer_1_2[4975:4968]};
      mid_2[2] = {1'b0,layer_2_2[4983:4976]} - {1'b0, layer_1_2[4983:4976]};
      btm_0[0] = {1'b0,layer_3_0[4967:4960]} - {1'b0, layer_2_0[4967:4960]};
      btm_0[1] = {1'b0,layer_3_0[4975:4968]} - {1'b0, layer_2_0[4975:4968]};
      btm_0[2] = {1'b0,layer_3_0[4983:4976]} - {1'b0, layer_2_0[4983:4976]};
      btm_1[0] = {1'b0,layer_3_1[4967:4960]} - {1'b0, layer_2_1[4967:4960]};
      btm_1[1] = {1'b0,layer_3_1[4975:4968]} - {1'b0, layer_2_1[4975:4968]};
      btm_1[2] = {1'b0,layer_3_1[4983:4976]} - {1'b0, layer_2_1[4983:4976]};
      btm_2[0] = {1'b0,layer_3_2[4967:4960]} - {1'b0, layer_2_2[4967:4960]};
      btm_2[1] = {1'b0,layer_3_2[4975:4968]} - {1'b0, layer_2_2[4975:4968]};
      btm_2[2] = {1'b0,layer_3_2[4983:4976]} - {1'b0, layer_2_2[4983:4976]};
    end
    'd622: begin
      top_0[0] = {1'b0,layer_1_0[4975:4968]} - {1'b0, layer_0_0[4975:4968]};
      top_0[1] = {1'b0,layer_1_0[4983:4976]} - {1'b0, layer_0_0[4983:4976]};
      top_0[2] = {1'b0,layer_1_0[4991:4984]} - {1'b0, layer_0_0[4991:4984]};
      top_1[0] = {1'b0,layer_1_1[4975:4968]} - {1'b0, layer_0_1[4975:4968]};
      top_1[1] = {1'b0,layer_1_1[4983:4976]} - {1'b0, layer_0_1[4983:4976]};
      top_1[2] = {1'b0,layer_1_1[4991:4984]} - {1'b0, layer_0_1[4991:4984]};
      top_2[0] = {1'b0,layer_1_2[4975:4968]} - {1'b0, layer_0_2[4975:4968]};
      top_2[1] = {1'b0,layer_1_2[4983:4976]} - {1'b0, layer_0_2[4983:4976]};
      top_2[2] = {1'b0,layer_1_2[4991:4984]} - {1'b0, layer_0_2[4991:4984]};
      mid_0[0] = {1'b0,layer_2_0[4975:4968]} - {1'b0, layer_1_0[4975:4968]};
      mid_0[1] = {1'b0,layer_2_0[4983:4976]} - {1'b0, layer_1_0[4983:4976]};
      mid_0[2] = {1'b0,layer_2_0[4991:4984]} - {1'b0, layer_1_0[4991:4984]};
      mid_1[0] = {1'b0,layer_2_1[4975:4968]} - {1'b0, layer_1_1[4975:4968]};
      mid_1[1] = {1'b0,layer_2_1[4983:4976]} - {1'b0, layer_1_1[4983:4976]};
      mid_1[2] = {1'b0,layer_2_1[4991:4984]} - {1'b0, layer_1_1[4991:4984]};
      mid_2[0] = {1'b0,layer_2_2[4975:4968]} - {1'b0, layer_1_2[4975:4968]};
      mid_2[1] = {1'b0,layer_2_2[4983:4976]} - {1'b0, layer_1_2[4983:4976]};
      mid_2[2] = {1'b0,layer_2_2[4991:4984]} - {1'b0, layer_1_2[4991:4984]};
      btm_0[0] = {1'b0,layer_3_0[4975:4968]} - {1'b0, layer_2_0[4975:4968]};
      btm_0[1] = {1'b0,layer_3_0[4983:4976]} - {1'b0, layer_2_0[4983:4976]};
      btm_0[2] = {1'b0,layer_3_0[4991:4984]} - {1'b0, layer_2_0[4991:4984]};
      btm_1[0] = {1'b0,layer_3_1[4975:4968]} - {1'b0, layer_2_1[4975:4968]};
      btm_1[1] = {1'b0,layer_3_1[4983:4976]} - {1'b0, layer_2_1[4983:4976]};
      btm_1[2] = {1'b0,layer_3_1[4991:4984]} - {1'b0, layer_2_1[4991:4984]};
      btm_2[0] = {1'b0,layer_3_2[4975:4968]} - {1'b0, layer_2_2[4975:4968]};
      btm_2[1] = {1'b0,layer_3_2[4983:4976]} - {1'b0, layer_2_2[4983:4976]};
      btm_2[2] = {1'b0,layer_3_2[4991:4984]} - {1'b0, layer_2_2[4991:4984]};
    end
    'd623: begin
      top_0[0] = {1'b0,layer_1_0[4983:4976]} - {1'b0, layer_0_0[4983:4976]};
      top_0[1] = {1'b0,layer_1_0[4991:4984]} - {1'b0, layer_0_0[4991:4984]};
      top_0[2] = {1'b0,layer_1_0[4999:4992]} - {1'b0, layer_0_0[4999:4992]};
      top_1[0] = {1'b0,layer_1_1[4983:4976]} - {1'b0, layer_0_1[4983:4976]};
      top_1[1] = {1'b0,layer_1_1[4991:4984]} - {1'b0, layer_0_1[4991:4984]};
      top_1[2] = {1'b0,layer_1_1[4999:4992]} - {1'b0, layer_0_1[4999:4992]};
      top_2[0] = {1'b0,layer_1_2[4983:4976]} - {1'b0, layer_0_2[4983:4976]};
      top_2[1] = {1'b0,layer_1_2[4991:4984]} - {1'b0, layer_0_2[4991:4984]};
      top_2[2] = {1'b0,layer_1_2[4999:4992]} - {1'b0, layer_0_2[4999:4992]};
      mid_0[0] = {1'b0,layer_2_0[4983:4976]} - {1'b0, layer_1_0[4983:4976]};
      mid_0[1] = {1'b0,layer_2_0[4991:4984]} - {1'b0, layer_1_0[4991:4984]};
      mid_0[2] = {1'b0,layer_2_0[4999:4992]} - {1'b0, layer_1_0[4999:4992]};
      mid_1[0] = {1'b0,layer_2_1[4983:4976]} - {1'b0, layer_1_1[4983:4976]};
      mid_1[1] = {1'b0,layer_2_1[4991:4984]} - {1'b0, layer_1_1[4991:4984]};
      mid_1[2] = {1'b0,layer_2_1[4999:4992]} - {1'b0, layer_1_1[4999:4992]};
      mid_2[0] = {1'b0,layer_2_2[4983:4976]} - {1'b0, layer_1_2[4983:4976]};
      mid_2[1] = {1'b0,layer_2_2[4991:4984]} - {1'b0, layer_1_2[4991:4984]};
      mid_2[2] = {1'b0,layer_2_2[4999:4992]} - {1'b0, layer_1_2[4999:4992]};
      btm_0[0] = {1'b0,layer_3_0[4983:4976]} - {1'b0, layer_2_0[4983:4976]};
      btm_0[1] = {1'b0,layer_3_0[4991:4984]} - {1'b0, layer_2_0[4991:4984]};
      btm_0[2] = {1'b0,layer_3_0[4999:4992]} - {1'b0, layer_2_0[4999:4992]};
      btm_1[0] = {1'b0,layer_3_1[4983:4976]} - {1'b0, layer_2_1[4983:4976]};
      btm_1[1] = {1'b0,layer_3_1[4991:4984]} - {1'b0, layer_2_1[4991:4984]};
      btm_1[2] = {1'b0,layer_3_1[4999:4992]} - {1'b0, layer_2_1[4999:4992]};
      btm_2[0] = {1'b0,layer_3_2[4983:4976]} - {1'b0, layer_2_2[4983:4976]};
      btm_2[1] = {1'b0,layer_3_2[4991:4984]} - {1'b0, layer_2_2[4991:4984]};
      btm_2[2] = {1'b0,layer_3_2[4999:4992]} - {1'b0, layer_2_2[4999:4992]};
    end
    'd624: begin
      top_0[0] = {1'b0,layer_1_0[4991:4984]} - {1'b0, layer_0_0[4991:4984]};
      top_0[1] = {1'b0,layer_1_0[4999:4992]} - {1'b0, layer_0_0[4999:4992]};
      top_0[2] = {1'b0,layer_1_0[5007:5000]} - {1'b0, layer_0_0[5007:5000]};
      top_1[0] = {1'b0,layer_1_1[4991:4984]} - {1'b0, layer_0_1[4991:4984]};
      top_1[1] = {1'b0,layer_1_1[4999:4992]} - {1'b0, layer_0_1[4999:4992]};
      top_1[2] = {1'b0,layer_1_1[5007:5000]} - {1'b0, layer_0_1[5007:5000]};
      top_2[0] = {1'b0,layer_1_2[4991:4984]} - {1'b0, layer_0_2[4991:4984]};
      top_2[1] = {1'b0,layer_1_2[4999:4992]} - {1'b0, layer_0_2[4999:4992]};
      top_2[2] = {1'b0,layer_1_2[5007:5000]} - {1'b0, layer_0_2[5007:5000]};
      mid_0[0] = {1'b0,layer_2_0[4991:4984]} - {1'b0, layer_1_0[4991:4984]};
      mid_0[1] = {1'b0,layer_2_0[4999:4992]} - {1'b0, layer_1_0[4999:4992]};
      mid_0[2] = {1'b0,layer_2_0[5007:5000]} - {1'b0, layer_1_0[5007:5000]};
      mid_1[0] = {1'b0,layer_2_1[4991:4984]} - {1'b0, layer_1_1[4991:4984]};
      mid_1[1] = {1'b0,layer_2_1[4999:4992]} - {1'b0, layer_1_1[4999:4992]};
      mid_1[2] = {1'b0,layer_2_1[5007:5000]} - {1'b0, layer_1_1[5007:5000]};
      mid_2[0] = {1'b0,layer_2_2[4991:4984]} - {1'b0, layer_1_2[4991:4984]};
      mid_2[1] = {1'b0,layer_2_2[4999:4992]} - {1'b0, layer_1_2[4999:4992]};
      mid_2[2] = {1'b0,layer_2_2[5007:5000]} - {1'b0, layer_1_2[5007:5000]};
      btm_0[0] = {1'b0,layer_3_0[4991:4984]} - {1'b0, layer_2_0[4991:4984]};
      btm_0[1] = {1'b0,layer_3_0[4999:4992]} - {1'b0, layer_2_0[4999:4992]};
      btm_0[2] = {1'b0,layer_3_0[5007:5000]} - {1'b0, layer_2_0[5007:5000]};
      btm_1[0] = {1'b0,layer_3_1[4991:4984]} - {1'b0, layer_2_1[4991:4984]};
      btm_1[1] = {1'b0,layer_3_1[4999:4992]} - {1'b0, layer_2_1[4999:4992]};
      btm_1[2] = {1'b0,layer_3_1[5007:5000]} - {1'b0, layer_2_1[5007:5000]};
      btm_2[0] = {1'b0,layer_3_2[4991:4984]} - {1'b0, layer_2_2[4991:4984]};
      btm_2[1] = {1'b0,layer_3_2[4999:4992]} - {1'b0, layer_2_2[4999:4992]};
      btm_2[2] = {1'b0,layer_3_2[5007:5000]} - {1'b0, layer_2_2[5007:5000]};
    end
    'd625: begin
      top_0[0] = {1'b0,layer_1_0[4999:4992]} - {1'b0, layer_0_0[4999:4992]};
      top_0[1] = {1'b0,layer_1_0[5007:5000]} - {1'b0, layer_0_0[5007:5000]};
      top_0[2] = {1'b0,layer_1_0[5015:5008]} - {1'b0, layer_0_0[5015:5008]};
      top_1[0] = {1'b0,layer_1_1[4999:4992]} - {1'b0, layer_0_1[4999:4992]};
      top_1[1] = {1'b0,layer_1_1[5007:5000]} - {1'b0, layer_0_1[5007:5000]};
      top_1[2] = {1'b0,layer_1_1[5015:5008]} - {1'b0, layer_0_1[5015:5008]};
      top_2[0] = {1'b0,layer_1_2[4999:4992]} - {1'b0, layer_0_2[4999:4992]};
      top_2[1] = {1'b0,layer_1_2[5007:5000]} - {1'b0, layer_0_2[5007:5000]};
      top_2[2] = {1'b0,layer_1_2[5015:5008]} - {1'b0, layer_0_2[5015:5008]};
      mid_0[0] = {1'b0,layer_2_0[4999:4992]} - {1'b0, layer_1_0[4999:4992]};
      mid_0[1] = {1'b0,layer_2_0[5007:5000]} - {1'b0, layer_1_0[5007:5000]};
      mid_0[2] = {1'b0,layer_2_0[5015:5008]} - {1'b0, layer_1_0[5015:5008]};
      mid_1[0] = {1'b0,layer_2_1[4999:4992]} - {1'b0, layer_1_1[4999:4992]};
      mid_1[1] = {1'b0,layer_2_1[5007:5000]} - {1'b0, layer_1_1[5007:5000]};
      mid_1[2] = {1'b0,layer_2_1[5015:5008]} - {1'b0, layer_1_1[5015:5008]};
      mid_2[0] = {1'b0,layer_2_2[4999:4992]} - {1'b0, layer_1_2[4999:4992]};
      mid_2[1] = {1'b0,layer_2_2[5007:5000]} - {1'b0, layer_1_2[5007:5000]};
      mid_2[2] = {1'b0,layer_2_2[5015:5008]} - {1'b0, layer_1_2[5015:5008]};
      btm_0[0] = {1'b0,layer_3_0[4999:4992]} - {1'b0, layer_2_0[4999:4992]};
      btm_0[1] = {1'b0,layer_3_0[5007:5000]} - {1'b0, layer_2_0[5007:5000]};
      btm_0[2] = {1'b0,layer_3_0[5015:5008]} - {1'b0, layer_2_0[5015:5008]};
      btm_1[0] = {1'b0,layer_3_1[4999:4992]} - {1'b0, layer_2_1[4999:4992]};
      btm_1[1] = {1'b0,layer_3_1[5007:5000]} - {1'b0, layer_2_1[5007:5000]};
      btm_1[2] = {1'b0,layer_3_1[5015:5008]} - {1'b0, layer_2_1[5015:5008]};
      btm_2[0] = {1'b0,layer_3_2[4999:4992]} - {1'b0, layer_2_2[4999:4992]};
      btm_2[1] = {1'b0,layer_3_2[5007:5000]} - {1'b0, layer_2_2[5007:5000]};
      btm_2[2] = {1'b0,layer_3_2[5015:5008]} - {1'b0, layer_2_2[5015:5008]};
    end
    'd626: begin
      top_0[0] = {1'b0,layer_1_0[5007:5000]} - {1'b0, layer_0_0[5007:5000]};
      top_0[1] = {1'b0,layer_1_0[5015:5008]} - {1'b0, layer_0_0[5015:5008]};
      top_0[2] = {1'b0,layer_1_0[5023:5016]} - {1'b0, layer_0_0[5023:5016]};
      top_1[0] = {1'b0,layer_1_1[5007:5000]} - {1'b0, layer_0_1[5007:5000]};
      top_1[1] = {1'b0,layer_1_1[5015:5008]} - {1'b0, layer_0_1[5015:5008]};
      top_1[2] = {1'b0,layer_1_1[5023:5016]} - {1'b0, layer_0_1[5023:5016]};
      top_2[0] = {1'b0,layer_1_2[5007:5000]} - {1'b0, layer_0_2[5007:5000]};
      top_2[1] = {1'b0,layer_1_2[5015:5008]} - {1'b0, layer_0_2[5015:5008]};
      top_2[2] = {1'b0,layer_1_2[5023:5016]} - {1'b0, layer_0_2[5023:5016]};
      mid_0[0] = {1'b0,layer_2_0[5007:5000]} - {1'b0, layer_1_0[5007:5000]};
      mid_0[1] = {1'b0,layer_2_0[5015:5008]} - {1'b0, layer_1_0[5015:5008]};
      mid_0[2] = {1'b0,layer_2_0[5023:5016]} - {1'b0, layer_1_0[5023:5016]};
      mid_1[0] = {1'b0,layer_2_1[5007:5000]} - {1'b0, layer_1_1[5007:5000]};
      mid_1[1] = {1'b0,layer_2_1[5015:5008]} - {1'b0, layer_1_1[5015:5008]};
      mid_1[2] = {1'b0,layer_2_1[5023:5016]} - {1'b0, layer_1_1[5023:5016]};
      mid_2[0] = {1'b0,layer_2_2[5007:5000]} - {1'b0, layer_1_2[5007:5000]};
      mid_2[1] = {1'b0,layer_2_2[5015:5008]} - {1'b0, layer_1_2[5015:5008]};
      mid_2[2] = {1'b0,layer_2_2[5023:5016]} - {1'b0, layer_1_2[5023:5016]};
      btm_0[0] = {1'b0,layer_3_0[5007:5000]} - {1'b0, layer_2_0[5007:5000]};
      btm_0[1] = {1'b0,layer_3_0[5015:5008]} - {1'b0, layer_2_0[5015:5008]};
      btm_0[2] = {1'b0,layer_3_0[5023:5016]} - {1'b0, layer_2_0[5023:5016]};
      btm_1[0] = {1'b0,layer_3_1[5007:5000]} - {1'b0, layer_2_1[5007:5000]};
      btm_1[1] = {1'b0,layer_3_1[5015:5008]} - {1'b0, layer_2_1[5015:5008]};
      btm_1[2] = {1'b0,layer_3_1[5023:5016]} - {1'b0, layer_2_1[5023:5016]};
      btm_2[0] = {1'b0,layer_3_2[5007:5000]} - {1'b0, layer_2_2[5007:5000]};
      btm_2[1] = {1'b0,layer_3_2[5015:5008]} - {1'b0, layer_2_2[5015:5008]};
      btm_2[2] = {1'b0,layer_3_2[5023:5016]} - {1'b0, layer_2_2[5023:5016]};
    end
    'd627: begin
      top_0[0] = {1'b0,layer_1_0[5015:5008]} - {1'b0, layer_0_0[5015:5008]};
      top_0[1] = {1'b0,layer_1_0[5023:5016]} - {1'b0, layer_0_0[5023:5016]};
      top_0[2] = {1'b0,layer_1_0[5031:5024]} - {1'b0, layer_0_0[5031:5024]};
      top_1[0] = {1'b0,layer_1_1[5015:5008]} - {1'b0, layer_0_1[5015:5008]};
      top_1[1] = {1'b0,layer_1_1[5023:5016]} - {1'b0, layer_0_1[5023:5016]};
      top_1[2] = {1'b0,layer_1_1[5031:5024]} - {1'b0, layer_0_1[5031:5024]};
      top_2[0] = {1'b0,layer_1_2[5015:5008]} - {1'b0, layer_0_2[5015:5008]};
      top_2[1] = {1'b0,layer_1_2[5023:5016]} - {1'b0, layer_0_2[5023:5016]};
      top_2[2] = {1'b0,layer_1_2[5031:5024]} - {1'b0, layer_0_2[5031:5024]};
      mid_0[0] = {1'b0,layer_2_0[5015:5008]} - {1'b0, layer_1_0[5015:5008]};
      mid_0[1] = {1'b0,layer_2_0[5023:5016]} - {1'b0, layer_1_0[5023:5016]};
      mid_0[2] = {1'b0,layer_2_0[5031:5024]} - {1'b0, layer_1_0[5031:5024]};
      mid_1[0] = {1'b0,layer_2_1[5015:5008]} - {1'b0, layer_1_1[5015:5008]};
      mid_1[1] = {1'b0,layer_2_1[5023:5016]} - {1'b0, layer_1_1[5023:5016]};
      mid_1[2] = {1'b0,layer_2_1[5031:5024]} - {1'b0, layer_1_1[5031:5024]};
      mid_2[0] = {1'b0,layer_2_2[5015:5008]} - {1'b0, layer_1_2[5015:5008]};
      mid_2[1] = {1'b0,layer_2_2[5023:5016]} - {1'b0, layer_1_2[5023:5016]};
      mid_2[2] = {1'b0,layer_2_2[5031:5024]} - {1'b0, layer_1_2[5031:5024]};
      btm_0[0] = {1'b0,layer_3_0[5015:5008]} - {1'b0, layer_2_0[5015:5008]};
      btm_0[1] = {1'b0,layer_3_0[5023:5016]} - {1'b0, layer_2_0[5023:5016]};
      btm_0[2] = {1'b0,layer_3_0[5031:5024]} - {1'b0, layer_2_0[5031:5024]};
      btm_1[0] = {1'b0,layer_3_1[5015:5008]} - {1'b0, layer_2_1[5015:5008]};
      btm_1[1] = {1'b0,layer_3_1[5023:5016]} - {1'b0, layer_2_1[5023:5016]};
      btm_1[2] = {1'b0,layer_3_1[5031:5024]} - {1'b0, layer_2_1[5031:5024]};
      btm_2[0] = {1'b0,layer_3_2[5015:5008]} - {1'b0, layer_2_2[5015:5008]};
      btm_2[1] = {1'b0,layer_3_2[5023:5016]} - {1'b0, layer_2_2[5023:5016]};
      btm_2[2] = {1'b0,layer_3_2[5031:5024]} - {1'b0, layer_2_2[5031:5024]};
    end
    'd628: begin
      top_0[0] = {1'b0,layer_1_0[5023:5016]} - {1'b0, layer_0_0[5023:5016]};
      top_0[1] = {1'b0,layer_1_0[5031:5024]} - {1'b0, layer_0_0[5031:5024]};
      top_0[2] = {1'b0,layer_1_0[5039:5032]} - {1'b0, layer_0_0[5039:5032]};
      top_1[0] = {1'b0,layer_1_1[5023:5016]} - {1'b0, layer_0_1[5023:5016]};
      top_1[1] = {1'b0,layer_1_1[5031:5024]} - {1'b0, layer_0_1[5031:5024]};
      top_1[2] = {1'b0,layer_1_1[5039:5032]} - {1'b0, layer_0_1[5039:5032]};
      top_2[0] = {1'b0,layer_1_2[5023:5016]} - {1'b0, layer_0_2[5023:5016]};
      top_2[1] = {1'b0,layer_1_2[5031:5024]} - {1'b0, layer_0_2[5031:5024]};
      top_2[2] = {1'b0,layer_1_2[5039:5032]} - {1'b0, layer_0_2[5039:5032]};
      mid_0[0] = {1'b0,layer_2_0[5023:5016]} - {1'b0, layer_1_0[5023:5016]};
      mid_0[1] = {1'b0,layer_2_0[5031:5024]} - {1'b0, layer_1_0[5031:5024]};
      mid_0[2] = {1'b0,layer_2_0[5039:5032]} - {1'b0, layer_1_0[5039:5032]};
      mid_1[0] = {1'b0,layer_2_1[5023:5016]} - {1'b0, layer_1_1[5023:5016]};
      mid_1[1] = {1'b0,layer_2_1[5031:5024]} - {1'b0, layer_1_1[5031:5024]};
      mid_1[2] = {1'b0,layer_2_1[5039:5032]} - {1'b0, layer_1_1[5039:5032]};
      mid_2[0] = {1'b0,layer_2_2[5023:5016]} - {1'b0, layer_1_2[5023:5016]};
      mid_2[1] = {1'b0,layer_2_2[5031:5024]} - {1'b0, layer_1_2[5031:5024]};
      mid_2[2] = {1'b0,layer_2_2[5039:5032]} - {1'b0, layer_1_2[5039:5032]};
      btm_0[0] = {1'b0,layer_3_0[5023:5016]} - {1'b0, layer_2_0[5023:5016]};
      btm_0[1] = {1'b0,layer_3_0[5031:5024]} - {1'b0, layer_2_0[5031:5024]};
      btm_0[2] = {1'b0,layer_3_0[5039:5032]} - {1'b0, layer_2_0[5039:5032]};
      btm_1[0] = {1'b0,layer_3_1[5023:5016]} - {1'b0, layer_2_1[5023:5016]};
      btm_1[1] = {1'b0,layer_3_1[5031:5024]} - {1'b0, layer_2_1[5031:5024]};
      btm_1[2] = {1'b0,layer_3_1[5039:5032]} - {1'b0, layer_2_1[5039:5032]};
      btm_2[0] = {1'b0,layer_3_2[5023:5016]} - {1'b0, layer_2_2[5023:5016]};
      btm_2[1] = {1'b0,layer_3_2[5031:5024]} - {1'b0, layer_2_2[5031:5024]};
      btm_2[2] = {1'b0,layer_3_2[5039:5032]} - {1'b0, layer_2_2[5039:5032]};
    end
    'd629: begin
      top_0[0] = {1'b0,layer_1_0[5031:5024]} - {1'b0, layer_0_0[5031:5024]};
      top_0[1] = {1'b0,layer_1_0[5039:5032]} - {1'b0, layer_0_0[5039:5032]};
      top_0[2] = {1'b0,layer_1_0[5047:5040]} - {1'b0, layer_0_0[5047:5040]};
      top_1[0] = {1'b0,layer_1_1[5031:5024]} - {1'b0, layer_0_1[5031:5024]};
      top_1[1] = {1'b0,layer_1_1[5039:5032]} - {1'b0, layer_0_1[5039:5032]};
      top_1[2] = {1'b0,layer_1_1[5047:5040]} - {1'b0, layer_0_1[5047:5040]};
      top_2[0] = {1'b0,layer_1_2[5031:5024]} - {1'b0, layer_0_2[5031:5024]};
      top_2[1] = {1'b0,layer_1_2[5039:5032]} - {1'b0, layer_0_2[5039:5032]};
      top_2[2] = {1'b0,layer_1_2[5047:5040]} - {1'b0, layer_0_2[5047:5040]};
      mid_0[0] = {1'b0,layer_2_0[5031:5024]} - {1'b0, layer_1_0[5031:5024]};
      mid_0[1] = {1'b0,layer_2_0[5039:5032]} - {1'b0, layer_1_0[5039:5032]};
      mid_0[2] = {1'b0,layer_2_0[5047:5040]} - {1'b0, layer_1_0[5047:5040]};
      mid_1[0] = {1'b0,layer_2_1[5031:5024]} - {1'b0, layer_1_1[5031:5024]};
      mid_1[1] = {1'b0,layer_2_1[5039:5032]} - {1'b0, layer_1_1[5039:5032]};
      mid_1[2] = {1'b0,layer_2_1[5047:5040]} - {1'b0, layer_1_1[5047:5040]};
      mid_2[0] = {1'b0,layer_2_2[5031:5024]} - {1'b0, layer_1_2[5031:5024]};
      mid_2[1] = {1'b0,layer_2_2[5039:5032]} - {1'b0, layer_1_2[5039:5032]};
      mid_2[2] = {1'b0,layer_2_2[5047:5040]} - {1'b0, layer_1_2[5047:5040]};
      btm_0[0] = {1'b0,layer_3_0[5031:5024]} - {1'b0, layer_2_0[5031:5024]};
      btm_0[1] = {1'b0,layer_3_0[5039:5032]} - {1'b0, layer_2_0[5039:5032]};
      btm_0[2] = {1'b0,layer_3_0[5047:5040]} - {1'b0, layer_2_0[5047:5040]};
      btm_1[0] = {1'b0,layer_3_1[5031:5024]} - {1'b0, layer_2_1[5031:5024]};
      btm_1[1] = {1'b0,layer_3_1[5039:5032]} - {1'b0, layer_2_1[5039:5032]};
      btm_1[2] = {1'b0,layer_3_1[5047:5040]} - {1'b0, layer_2_1[5047:5040]};
      btm_2[0] = {1'b0,layer_3_2[5031:5024]} - {1'b0, layer_2_2[5031:5024]};
      btm_2[1] = {1'b0,layer_3_2[5039:5032]} - {1'b0, layer_2_2[5039:5032]};
      btm_2[2] = {1'b0,layer_3_2[5047:5040]} - {1'b0, layer_2_2[5047:5040]};
    end
    'd630: begin
      top_0[0] = {1'b0,layer_1_0[5039:5032]} - {1'b0, layer_0_0[5039:5032]};
      top_0[1] = {1'b0,layer_1_0[5047:5040]} - {1'b0, layer_0_0[5047:5040]};
      top_0[2] = {1'b0,layer_1_0[5055:5048]} - {1'b0, layer_0_0[5055:5048]};
      top_1[0] = {1'b0,layer_1_1[5039:5032]} - {1'b0, layer_0_1[5039:5032]};
      top_1[1] = {1'b0,layer_1_1[5047:5040]} - {1'b0, layer_0_1[5047:5040]};
      top_1[2] = {1'b0,layer_1_1[5055:5048]} - {1'b0, layer_0_1[5055:5048]};
      top_2[0] = {1'b0,layer_1_2[5039:5032]} - {1'b0, layer_0_2[5039:5032]};
      top_2[1] = {1'b0,layer_1_2[5047:5040]} - {1'b0, layer_0_2[5047:5040]};
      top_2[2] = {1'b0,layer_1_2[5055:5048]} - {1'b0, layer_0_2[5055:5048]};
      mid_0[0] = {1'b0,layer_2_0[5039:5032]} - {1'b0, layer_1_0[5039:5032]};
      mid_0[1] = {1'b0,layer_2_0[5047:5040]} - {1'b0, layer_1_0[5047:5040]};
      mid_0[2] = {1'b0,layer_2_0[5055:5048]} - {1'b0, layer_1_0[5055:5048]};
      mid_1[0] = {1'b0,layer_2_1[5039:5032]} - {1'b0, layer_1_1[5039:5032]};
      mid_1[1] = {1'b0,layer_2_1[5047:5040]} - {1'b0, layer_1_1[5047:5040]};
      mid_1[2] = {1'b0,layer_2_1[5055:5048]} - {1'b0, layer_1_1[5055:5048]};
      mid_2[0] = {1'b0,layer_2_2[5039:5032]} - {1'b0, layer_1_2[5039:5032]};
      mid_2[1] = {1'b0,layer_2_2[5047:5040]} - {1'b0, layer_1_2[5047:5040]};
      mid_2[2] = {1'b0,layer_2_2[5055:5048]} - {1'b0, layer_1_2[5055:5048]};
      btm_0[0] = {1'b0,layer_3_0[5039:5032]} - {1'b0, layer_2_0[5039:5032]};
      btm_0[1] = {1'b0,layer_3_0[5047:5040]} - {1'b0, layer_2_0[5047:5040]};
      btm_0[2] = {1'b0,layer_3_0[5055:5048]} - {1'b0, layer_2_0[5055:5048]};
      btm_1[0] = {1'b0,layer_3_1[5039:5032]} - {1'b0, layer_2_1[5039:5032]};
      btm_1[1] = {1'b0,layer_3_1[5047:5040]} - {1'b0, layer_2_1[5047:5040]};
      btm_1[2] = {1'b0,layer_3_1[5055:5048]} - {1'b0, layer_2_1[5055:5048]};
      btm_2[0] = {1'b0,layer_3_2[5039:5032]} - {1'b0, layer_2_2[5039:5032]};
      btm_2[1] = {1'b0,layer_3_2[5047:5040]} - {1'b0, layer_2_2[5047:5040]};
      btm_2[2] = {1'b0,layer_3_2[5055:5048]} - {1'b0, layer_2_2[5055:5048]};
    end
    default: begin
      top_0[0] = 'd0;
      top_0[1] = 'd0;
      top_0[2] = 'd0;
      top_1[0] = 'd0;
      top_1[1] = 'd0;
      top_1[2] = 'd0;
      top_2[0] = 'd0;
      top_2[1] = 'd0;
      top_2[2] = 'd0;
      mid_0[0] = 'd0;
      mid_0[1] = 'd0;
      mid_0[2] = 'd0;
      mid_1[0] = 'd0;
      mid_1[1] = 'd0;
      mid_1[2] = 'd0;
      mid_2[0] = 'd0;
      mid_2[1] = 'd0;
      mid_2[2] = 'd0;
      btm_0[0] = 'd0;
      btm_0[1] = 'd0;
      btm_0[2] = 'd0;
      btm_1[0] = 'd0;
      btm_1[1] = 'd0;
      btm_1[2] = 'd0;
      btm_2[0] = 'd0;
      btm_2[1] = 'd0;
      btm_2[2] = 'd0;
    end
  endcase
end

reg    [11:0]      detect_max; //wire
always@(*) begin
  if(mid_1[1] > top_0[1])
    detect_max[0] = 1;
  else
    detect_max[0] = 0;
  if(mid_1[1] > top_1[0])
    detect_max[1] = 1;
  else
    detect_max[1] = 0;
  if(mid_1[1] > top_1[2])
    detect_max[2] = 1;
  else
    detect_max[2] = 0;
  if(mid_1[1] > top_2[1])
    detect_max[3] = 1;
  else
    detect_max[3] = 0;
  if(mid_1[1] > mid_0[0])
    detect_max[4] = 1;
  else
    detect_max[4] = 0;
  if(mid_1[1] > mid_0[2])
    detect_max[5] = 1;
  else
    detect_max[5] = 0;
  if(mid_1[1] > mid_2[0])
    detect_max[6] = 1;
  else
    detect_max[6] = 0;
  if(mid_1[1] > mid_2[2])
    detect_max[7] = 1;
  else
    detect_max[7] = 0;
  if(mid_1[1] > btm_0[1])
    detect_max[8] = 1;
  else
    detect_max[8] = 0;
  if(mid_1[1] > btm_1[0])
    detect_max[9] = 1;
  else
    detect_max[9] = 0;
  if(mid_1[1] > btm_1[2])
    detect_max[10] = 1;
  else
    detect_max[10] = 0;
  if(mid_1[1] > btm_2[1])
    detect_max[11] = 1;
  else
    detect_max[11] = 0;
end

reg    [11:0]      detect_min; //wire
always@(*) begin
  if(mid_1[1] < top_0[1])
    detect_min[0] = 1;
  else
    detect_min[0] = 0;
  if(mid_1[1] < top_1[0])
    detect_min[1] = 1;
  else
    detect_min[1] = 0;
  if(mid_1[1] < top_1[2])
    detect_min[2] = 1;
  else
    detect_min[2] = 0;
  if(mid_1[1] < top_2[1])
    detect_min[3] = 1;
  else
    detect_min[3] = 0;
  if(mid_1[1] < mid_0[0])
    detect_min[4] = 1;
  else
    detect_min[4] = 0;
  if(mid_1[1] < mid_0[2])
    detect_min[5] = 1;
  else
    detect_min[5] = 0;
  if(mid_1[1] < mid_2[0])
    detect_min[6] = 1;
  else
    detect_min[6] = 0;
  if(mid_1[1] < mid_2[2])
    detect_min[7] = 1;
  else
    detect_min[7] = 0;
  if(mid_1[1] < btm_0[1])
    detect_min[8] = 1;
  else
    detect_min[8] = 0;
  if(mid_1[1] < btm_1[0])
    detect_min[9] = 1;
  else
    detect_min[9] = 0;
  if(mid_1[1] < btm_1[2])
    detect_min[10] = 1;
  else
    detect_min[10] = 0;
  if(mid_1[1] < btm_2[1])
    detect_min[11] = 1;
  else
    detect_min[11] = 0;
end

wire is_max = (&detect_max) ? 1:0;
wire is_min = (&detect_min) ? 1:0;
assign is_keypoint = is_max | is_min;

endmodule