module Gaussian_Blur_7x7(
  clk,
  rst_n,
  buffer_data_0,
  buffer_data_1,
  buffer_data_2,
  buffer_data_3,
  buffer_data_4,
  buffer_data_5,
  buffer_data_6,
  current_col,
  blur_out,
  start,
  done
);

input                 clk;
input                 rst_n;
input                 start;
output                done;
input         [5:0]   current_col;
input       [175:0]   buffer_data_0;
input       [175:0]   buffer_data_1;
input       [175:0]   buffer_data_2;
input       [175:0]   buffer_data_3;
input       [175:0]   buffer_data_4;
input       [175:0]   buffer_data_5;
input       [175:0]   buffer_data_6;
output reg  [127:0]   blur_out; // wire

parameter  ST_MUX         = 0,
           ST_MUL         = 1,
           ST_ADD         = 2,
           ST_UPDATE      = 3;
reg     [2:0] current_state,
              next_state;
assign done = (current_state==ST_UPDATE) ? 1 : 0;

wire       [55:0] G_Kernel_7x7_0;
wire       [55:0] G_Kernel_7x7_1;
wire       [55:0] G_Kernel_7x7_2;
wire       [55:0] G_Kernel_7x7_3;
assign  G_Kernel_7x7_0[7:0]   = 8'h03; //C6EBCB; //18'b000000111100011011;//'d014754;
assign  G_Kernel_7x7_0[15:8]  = 8'h04; //6AA8A8; //18'b000001000110101010;//'d017252;
assign  G_Kernel_7x7_0[23:16] = 8'h04; //D9ED31; //18'b000001001101100111;//'d018950;
assign  G_Kernel_7x7_0[31:24] = 8'h05; //0165DE; //18'b000001010000000101;//'d019552;
assign  G_Kernel_7x7_0[39:32] = 8'h04; //D9ED31; //18'b000001001101100111;//'d018950;
assign  G_Kernel_7x7_0[47:40] = 8'h04; //6AA8A8; //18'b000001000110101010;//'d017252;
assign  G_Kernel_7x7_0[55:48] = 8'h03; //C6EBCB; //18'b000000111100011011;//'d014754;
assign  G_Kernel_7x7_1[7:0]   = 8'h04; //6AA8A8; //18'b000001000110101010;//'d017252;
assign  G_Kernel_7x7_1[15:8]  = 8'h05; //2A1FB1; //18'b000001010010101000;//'d020174;
assign  G_Kernel_7x7_1[23:16] = 8'h05; //AC3BC7; //18'b000001011010110000;//'d022159;
assign  G_Kernel_7x7_1[31:24] = 8'h05; //DA6392; //18'b000001011101101001;//'d022863;
assign  G_Kernel_7x7_1[39:32] = 8'h05; //AC3BC7; //18'b000001011010110000;//'d022159;
assign  G_Kernel_7x7_1[47:40] = 8'h05; //2A1FB1; //18'b000001010010101000;//'d020174;
assign  G_Kernel_7x7_1[55:48] = 8'h04; //6AA8A8; //18'b000001000110101010;//'d017252;
assign  G_Kernel_7x7_2[7:0]   = 8'h04; //D9ED31; //18'b000001001101100111;//'d018950;
assign  G_Kernel_7x7_2[15:8]  = 8'h05; //AC3BC7; //18'b000001011010110000;//'d022159;
assign  G_Kernel_7x7_2[23:16] = 8'h06; //3B25B2; //18'b000001100011101100;//'d024340;
assign  G_Kernel_7x7_2[31:24] = 8'h06; //6DD847; //18'b000001100110110111;//'d025113;
assign  G_Kernel_7x7_2[39:32] = 8'h06; //3B25B2; //18'b000001100011101100;//'d024340;
assign  G_Kernel_7x7_2[47:40] = 8'h05; //AC3BC7; //18'b000001011010110000;//'d022159;
assign  G_Kernel_7x7_2[55:48] = 8'h04; //D9ED31; //18'b000001001101100111;//'d018950;
assign  G_Kernel_7x7_3[7:0]   = 8'h05; //0165DE; //18'b000001010000000101;//'d019552;
assign  G_Kernel_7x7_3[15:8]  = 8'h05; //DA6392; //18'b000001011101101001;//'d022863;
assign  G_Kernel_7x7_3[23:16] = 8'h06; //6DD847; //18'b000001100110110111;//'d025113;
assign  G_Kernel_7x7_3[31:24] = 8'h06; //A2275A; //18'b000001101010001000;//'d025911;
assign  G_Kernel_7x7_3[39:32] = 8'h06; //6DD847; //18'b000001100110110111;//'d025113;
assign  G_Kernel_7x7_3[47:40] = 8'h05; //DA6392; //18'b000001011101101001;//'d022863;
assign  G_Kernel_7x7_3[55:48] = 8'h05; //0165DE; //18'b000001010000000101;//'d019552;

reg    [55:0]    layer0[0:15]; //wire
reg    [55:0]    layer1[0:15]; //wire
reg    [55:0]    layer2[0:15]; //wire
reg    [55:0]    layer3[0:15]; //wire
reg    [55:0]    layer4[0:15]; //wire
reg    [55:0]    layer5[0:15]; //wire
reg    [55:0]    layer6[0:15]; //wire
always @(posedge clk) begin
  if(!rst_n) begin
    layer0[0] <= 'd0;
    layer0[1] <= 'd0;
    layer0[2] <= 'd0;
    layer0[3] <= 'd0;
    layer0[4] <= 'd0;
    layer0[5] <= 'd0;
    layer0[6] <= 'd0;
    layer0[7] <= 'd0;
    layer0[8] <= 'd0;
    layer0[9] <= 'd0;
    layer0[10] <= 'd0;
    layer0[11] <= 'd0;
    layer0[12] <= 'd0;
    layer0[13] <= 'd0;
    layer0[14] <= 'd0;
    layer0[15] <= 'd0;
    layer1[0] <= 'd0;
    layer1[1] <= 'd0;
    layer1[2] <= 'd0;
    layer1[3] <= 'd0;
    layer1[4] <= 'd0;
    layer1[5] <= 'd0;
    layer1[6] <= 'd0;
    layer1[7] <= 'd0;
    layer1[8] <= 'd0;
    layer1[9] <= 'd0;
    layer1[10] <= 'd0;
    layer1[11] <= 'd0;
    layer1[12] <= 'd0;
    layer1[13] <= 'd0;
    layer1[14] <= 'd0;
    layer1[15] <= 'd0;
    layer2[0] <= 'd0;
    layer2[1] <= 'd0;
    layer2[2] <= 'd0;
    layer2[3] <= 'd0;
    layer2[4] <= 'd0;
    layer2[5] <= 'd0;
    layer2[6] <= 'd0;
    layer2[7] <= 'd0;
    layer2[8] <= 'd0;
    layer2[9] <= 'd0;
    layer2[10] <= 'd0;
    layer2[11] <= 'd0;
    layer2[12] <= 'd0;
    layer2[13] <= 'd0;
    layer2[14] <= 'd0;
    layer2[15] <= 'd0;
    layer3[0] <= 'd0;
    layer3[1] <= 'd0;
    layer3[2] <= 'd0;
    layer3[3] <= 'd0;
    layer3[4] <= 'd0;
    layer3[5] <= 'd0;
    layer3[6] <= 'd0;
    layer3[7] <= 'd0;
    layer3[8] <= 'd0;
    layer3[9] <= 'd0;
    layer3[10] <= 'd0;
    layer3[11] <= 'd0;
    layer3[12] <= 'd0;
    layer3[13] <= 'd0;
    layer3[14] <= 'd0;
    layer3[15] <= 'd0;
    layer4[0] <= 'd0;
    layer4[1] <= 'd0;
    layer4[2] <= 'd0;
    layer4[3] <= 'd0;
    layer4[4] <= 'd0;
    layer4[5] <= 'd0;
    layer4[6] <= 'd0;
    layer4[7] <= 'd0;
    layer4[8] <= 'd0;
    layer4[9] <= 'd0;
    layer4[10] <= 'd0;
    layer4[11] <= 'd0;
    layer4[12] <= 'd0;
    layer4[13] <= 'd0;
    layer4[14] <= 'd0;
    layer4[15] <= 'd0;
    layer5[0] <= 'd0;
    layer5[1] <= 'd0;
    layer5[2] <= 'd0;
    layer5[3] <= 'd0;
    layer5[4] <= 'd0;
    layer5[5] <= 'd0;
    layer5[6] <= 'd0;
    layer5[7] <= 'd0;
    layer5[8] <= 'd0;
    layer5[9] <= 'd0;
    layer5[10] <= 'd0;
    layer5[11] <= 'd0;
    layer5[12] <= 'd0;
    layer5[13] <= 'd0;
    layer5[14] <= 'd0;
    layer5[15] <= 'd0;
    layer6[0] <= 'd0;
    layer6[1] <= 'd0;
    layer6[2] <= 'd0;
    layer6[3] <= 'd0;
    layer6[4] <= 'd0;
    layer6[5] <= 'd0;
    layer6[6] <= 'd0;
    layer6[7] <= 'd0;
    layer6[8] <= 'd0;
    layer6[9] <= 'd0;
    layer6[10] <= 'd0;
    layer6[11] <= 'd0;
    layer6[12] <= 'd0;
    layer6[13] <= 'd0;
    layer6[14] <= 'd0;
    layer6[15] <= 'd0;
  end
  else if(current_state==ST_MUX) begin
    case(current_col)
      'd0: begin
        layer0[0][7:0] <= 0;
        layer0[0][15:8] <= 0;
        layer0[0][23:16] <= 0;
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= 0;
        layer1[0][15:8] <= 0;
        layer1[0][23:16] <= 0;
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= 0;
        layer2[0][15:8] <= 0;
        layer2[0][23:16] <= 0;
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= 0;
        layer3[0][15:8] <= 0;
        layer3[0][23:16] <= 0;
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= 0;
        layer4[0][15:8] <= 0;
        layer4[0][23:16] <= 0;
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= 0;
        layer5[0][15:8] <= 0;
        layer5[0][23:16] <= 0;
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= 0;
        layer6[0][15:8] <= 0;
        layer6[0][23:16] <= 0;
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= 0;
        layer0[1][15:8] <= 0;
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= 0;
        layer1[1][15:8] <= 0;
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= 0;
        layer2[1][15:8] <= 0;
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= 0;
        layer3[1][15:8] <= 0;
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= 0;
        layer4[1][15:8] <= 0;
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= 0;
        layer5[1][15:8] <= 0;
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= 0;
        layer6[1][15:8] <= 0;
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= 0;
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= 0;
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= 0;
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= 0;
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= 0;
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= 0;
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= 0;
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd1: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd2: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd3: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd4: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd5: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd6: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd7: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd8: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd9: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd10: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd11: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd12: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd13: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd14: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd15: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd16: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd17: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd18: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd19: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd20: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd21: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd22: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd23: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd24: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd25: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd26: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd27: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd28: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd29: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd30: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd31: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd32: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd33: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd34: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd35: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd36: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd37: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd38: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= buffer_data_6[159:152];
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= buffer_data_5[159:152];
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= buffer_data_4[159:152];
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= buffer_data_3[159:152];
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= buffer_data_2[159:152];
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= buffer_data_1[159:152];
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= buffer_data_0[159:152];
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= buffer_data_6[159:152];
        layer0[14][55:48] <= buffer_data_6[167:160];
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= buffer_data_5[159:152];
        layer1[14][55:48] <= buffer_data_5[167:160];
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= buffer_data_4[159:152];
        layer2[14][55:48] <= buffer_data_4[167:160];
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= buffer_data_3[159:152];
        layer3[14][55:48] <= buffer_data_3[167:160];
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= buffer_data_2[159:152];
        layer4[14][55:48] <= buffer_data_2[167:160];
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= buffer_data_1[159:152];
        layer5[14][55:48] <= buffer_data_1[167:160];
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= buffer_data_0[159:152];
        layer6[14][55:48] <= buffer_data_0[167:160];
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= buffer_data_6[159:152];
        layer0[15][47:40] <= buffer_data_6[167:160];
        layer0[15][55:48] <= buffer_data_6[175:168];
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= buffer_data_5[159:152];
        layer1[15][47:40] <= buffer_data_5[167:160];
        layer1[15][55:48] <= buffer_data_5[175:168];
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= buffer_data_4[159:152];
        layer2[15][47:40] <= buffer_data_4[167:160];
        layer2[15][55:48] <= buffer_data_4[175:168];
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= buffer_data_3[159:152];
        layer3[15][47:40] <= buffer_data_3[167:160];
        layer3[15][55:48] <= buffer_data_3[175:168];
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= buffer_data_2[159:152];
        layer4[15][47:40] <= buffer_data_2[167:160];
        layer4[15][55:48] <= buffer_data_2[175:168];
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= buffer_data_1[159:152];
        layer5[15][47:40] <= buffer_data_1[167:160];
        layer5[15][55:48] <= buffer_data_1[175:168];
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= buffer_data_0[159:152];
        layer6[15][47:40] <= buffer_data_0[167:160];
        layer6[15][55:48] <= buffer_data_0[175:168];
    end
      'd39: begin
        layer0[0][7:0] <= buffer_data_6[7:0];
        layer0[0][15:8] <= buffer_data_6[15:8];
        layer0[0][23:16] <= buffer_data_6[23:16];
        layer0[0][31:24] <= buffer_data_6[31:24];
        layer0[0][39:32] <= buffer_data_6[39:32];
        layer0[0][47:40] <= buffer_data_6[47:40];
        layer0[0][55:48] <= buffer_data_6[55:48];
        layer1[0][7:0] <= buffer_data_5[7:0];
        layer1[0][15:8] <= buffer_data_5[15:8];
        layer1[0][23:16] <= buffer_data_5[23:16];
        layer1[0][31:24] <= buffer_data_5[31:24];
        layer1[0][39:32] <= buffer_data_5[39:32];
        layer1[0][47:40] <= buffer_data_5[47:40];
        layer1[0][55:48] <= buffer_data_5[55:48];
        layer2[0][7:0] <= buffer_data_4[7:0];
        layer2[0][15:8] <= buffer_data_4[15:8];
        layer2[0][23:16] <= buffer_data_4[23:16];
        layer2[0][31:24] <= buffer_data_4[31:24];
        layer2[0][39:32] <= buffer_data_4[39:32];
        layer2[0][47:40] <= buffer_data_4[47:40];
        layer2[0][55:48] <= buffer_data_4[55:48];
        layer3[0][7:0] <= buffer_data_3[7:0];
        layer3[0][15:8] <= buffer_data_3[15:8];
        layer3[0][23:16] <= buffer_data_3[23:16];
        layer3[0][31:24] <= buffer_data_3[31:24];
        layer3[0][39:32] <= buffer_data_3[39:32];
        layer3[0][47:40] <= buffer_data_3[47:40];
        layer3[0][55:48] <= buffer_data_3[55:48];
        layer4[0][7:0] <= buffer_data_2[7:0];
        layer4[0][15:8] <= buffer_data_2[15:8];
        layer4[0][23:16] <= buffer_data_2[23:16];
        layer4[0][31:24] <= buffer_data_2[31:24];
        layer4[0][39:32] <= buffer_data_2[39:32];
        layer4[0][47:40] <= buffer_data_2[47:40];
        layer4[0][55:48] <= buffer_data_2[55:48];
        layer5[0][7:0] <= buffer_data_1[7:0];
        layer5[0][15:8] <= buffer_data_1[15:8];
        layer5[0][23:16] <= buffer_data_1[23:16];
        layer5[0][31:24] <= buffer_data_1[31:24];
        layer5[0][39:32] <= buffer_data_1[39:32];
        layer5[0][47:40] <= buffer_data_1[47:40];
        layer5[0][55:48] <= buffer_data_1[55:48];
        layer6[0][7:0] <= buffer_data_0[7:0];
        layer6[0][15:8] <= buffer_data_0[15:8];
        layer6[0][23:16] <= buffer_data_0[23:16];
        layer6[0][31:24] <= buffer_data_0[31:24];
        layer6[0][39:32] <= buffer_data_0[39:32];
        layer6[0][47:40] <= buffer_data_0[47:40];
        layer6[0][55:48] <= buffer_data_0[55:48];
        layer0[1][7:0] <= buffer_data_6[15:8];
        layer0[1][15:8] <= buffer_data_6[23:16];
        layer0[1][23:16] <= buffer_data_6[31:24];
        layer0[1][31:24] <= buffer_data_6[39:32];
        layer0[1][39:32] <= buffer_data_6[47:40];
        layer0[1][47:40] <= buffer_data_6[55:48];
        layer0[1][55:48] <= buffer_data_6[63:56];
        layer1[1][7:0] <= buffer_data_5[15:8];
        layer1[1][15:8] <= buffer_data_5[23:16];
        layer1[1][23:16] <= buffer_data_5[31:24];
        layer1[1][31:24] <= buffer_data_5[39:32];
        layer1[1][39:32] <= buffer_data_5[47:40];
        layer1[1][47:40] <= buffer_data_5[55:48];
        layer1[1][55:48] <= buffer_data_5[63:56];
        layer2[1][7:0] <= buffer_data_4[15:8];
        layer2[1][15:8] <= buffer_data_4[23:16];
        layer2[1][23:16] <= buffer_data_4[31:24];
        layer2[1][31:24] <= buffer_data_4[39:32];
        layer2[1][39:32] <= buffer_data_4[47:40];
        layer2[1][47:40] <= buffer_data_4[55:48];
        layer2[1][55:48] <= buffer_data_4[63:56];
        layer3[1][7:0] <= buffer_data_3[15:8];
        layer3[1][15:8] <= buffer_data_3[23:16];
        layer3[1][23:16] <= buffer_data_3[31:24];
        layer3[1][31:24] <= buffer_data_3[39:32];
        layer3[1][39:32] <= buffer_data_3[47:40];
        layer3[1][47:40] <= buffer_data_3[55:48];
        layer3[1][55:48] <= buffer_data_3[63:56];
        layer4[1][7:0] <= buffer_data_2[15:8];
        layer4[1][15:8] <= buffer_data_2[23:16];
        layer4[1][23:16] <= buffer_data_2[31:24];
        layer4[1][31:24] <= buffer_data_2[39:32];
        layer4[1][39:32] <= buffer_data_2[47:40];
        layer4[1][47:40] <= buffer_data_2[55:48];
        layer4[1][55:48] <= buffer_data_2[63:56];
        layer5[1][7:0] <= buffer_data_1[15:8];
        layer5[1][15:8] <= buffer_data_1[23:16];
        layer5[1][23:16] <= buffer_data_1[31:24];
        layer5[1][31:24] <= buffer_data_1[39:32];
        layer5[1][39:32] <= buffer_data_1[47:40];
        layer5[1][47:40] <= buffer_data_1[55:48];
        layer5[1][55:48] <= buffer_data_1[63:56];
        layer6[1][7:0] <= buffer_data_0[15:8];
        layer6[1][15:8] <= buffer_data_0[23:16];
        layer6[1][23:16] <= buffer_data_0[31:24];
        layer6[1][31:24] <= buffer_data_0[39:32];
        layer6[1][39:32] <= buffer_data_0[47:40];
        layer6[1][47:40] <= buffer_data_0[55:48];
        layer6[1][55:48] <= buffer_data_0[63:56];
        layer0[2][7:0] <= buffer_data_6[23:16];
        layer0[2][15:8] <= buffer_data_6[31:24];
        layer0[2][23:16] <= buffer_data_6[39:32];
        layer0[2][31:24] <= buffer_data_6[47:40];
        layer0[2][39:32] <= buffer_data_6[55:48];
        layer0[2][47:40] <= buffer_data_6[63:56];
        layer0[2][55:48] <= buffer_data_6[71:64];
        layer1[2][7:0] <= buffer_data_5[23:16];
        layer1[2][15:8] <= buffer_data_5[31:24];
        layer1[2][23:16] <= buffer_data_5[39:32];
        layer1[2][31:24] <= buffer_data_5[47:40];
        layer1[2][39:32] <= buffer_data_5[55:48];
        layer1[2][47:40] <= buffer_data_5[63:56];
        layer1[2][55:48] <= buffer_data_5[71:64];
        layer2[2][7:0] <= buffer_data_4[23:16];
        layer2[2][15:8] <= buffer_data_4[31:24];
        layer2[2][23:16] <= buffer_data_4[39:32];
        layer2[2][31:24] <= buffer_data_4[47:40];
        layer2[2][39:32] <= buffer_data_4[55:48];
        layer2[2][47:40] <= buffer_data_4[63:56];
        layer2[2][55:48] <= buffer_data_4[71:64];
        layer3[2][7:0] <= buffer_data_3[23:16];
        layer3[2][15:8] <= buffer_data_3[31:24];
        layer3[2][23:16] <= buffer_data_3[39:32];
        layer3[2][31:24] <= buffer_data_3[47:40];
        layer3[2][39:32] <= buffer_data_3[55:48];
        layer3[2][47:40] <= buffer_data_3[63:56];
        layer3[2][55:48] <= buffer_data_3[71:64];
        layer4[2][7:0] <= buffer_data_2[23:16];
        layer4[2][15:8] <= buffer_data_2[31:24];
        layer4[2][23:16] <= buffer_data_2[39:32];
        layer4[2][31:24] <= buffer_data_2[47:40];
        layer4[2][39:32] <= buffer_data_2[55:48];
        layer4[2][47:40] <= buffer_data_2[63:56];
        layer4[2][55:48] <= buffer_data_2[71:64];
        layer5[2][7:0] <= buffer_data_1[23:16];
        layer5[2][15:8] <= buffer_data_1[31:24];
        layer5[2][23:16] <= buffer_data_1[39:32];
        layer5[2][31:24] <= buffer_data_1[47:40];
        layer5[2][39:32] <= buffer_data_1[55:48];
        layer5[2][47:40] <= buffer_data_1[63:56];
        layer5[2][55:48] <= buffer_data_1[71:64];
        layer6[2][7:0] <= buffer_data_0[23:16];
        layer6[2][15:8] <= buffer_data_0[31:24];
        layer6[2][23:16] <= buffer_data_0[39:32];
        layer6[2][31:24] <= buffer_data_0[47:40];
        layer6[2][39:32] <= buffer_data_0[55:48];
        layer6[2][47:40] <= buffer_data_0[63:56];
        layer6[2][55:48] <= buffer_data_0[71:64];
        layer0[3][7:0] <= buffer_data_6[31:24];
        layer0[3][15:8] <= buffer_data_6[39:32];
        layer0[3][23:16] <= buffer_data_6[47:40];
        layer0[3][31:24] <= buffer_data_6[55:48];
        layer0[3][39:32] <= buffer_data_6[63:56];
        layer0[3][47:40] <= buffer_data_6[71:64];
        layer0[3][55:48] <= buffer_data_6[79:72];
        layer1[3][7:0] <= buffer_data_5[31:24];
        layer1[3][15:8] <= buffer_data_5[39:32];
        layer1[3][23:16] <= buffer_data_5[47:40];
        layer1[3][31:24] <= buffer_data_5[55:48];
        layer1[3][39:32] <= buffer_data_5[63:56];
        layer1[3][47:40] <= buffer_data_5[71:64];
        layer1[3][55:48] <= buffer_data_5[79:72];
        layer2[3][7:0] <= buffer_data_4[31:24];
        layer2[3][15:8] <= buffer_data_4[39:32];
        layer2[3][23:16] <= buffer_data_4[47:40];
        layer2[3][31:24] <= buffer_data_4[55:48];
        layer2[3][39:32] <= buffer_data_4[63:56];
        layer2[3][47:40] <= buffer_data_4[71:64];
        layer2[3][55:48] <= buffer_data_4[79:72];
        layer3[3][7:0] <= buffer_data_3[31:24];
        layer3[3][15:8] <= buffer_data_3[39:32];
        layer3[3][23:16] <= buffer_data_3[47:40];
        layer3[3][31:24] <= buffer_data_3[55:48];
        layer3[3][39:32] <= buffer_data_3[63:56];
        layer3[3][47:40] <= buffer_data_3[71:64];
        layer3[3][55:48] <= buffer_data_3[79:72];
        layer4[3][7:0] <= buffer_data_2[31:24];
        layer4[3][15:8] <= buffer_data_2[39:32];
        layer4[3][23:16] <= buffer_data_2[47:40];
        layer4[3][31:24] <= buffer_data_2[55:48];
        layer4[3][39:32] <= buffer_data_2[63:56];
        layer4[3][47:40] <= buffer_data_2[71:64];
        layer4[3][55:48] <= buffer_data_2[79:72];
        layer5[3][7:0] <= buffer_data_1[31:24];
        layer5[3][15:8] <= buffer_data_1[39:32];
        layer5[3][23:16] <= buffer_data_1[47:40];
        layer5[3][31:24] <= buffer_data_1[55:48];
        layer5[3][39:32] <= buffer_data_1[63:56];
        layer5[3][47:40] <= buffer_data_1[71:64];
        layer5[3][55:48] <= buffer_data_1[79:72];
        layer6[3][7:0] <= buffer_data_0[31:24];
        layer6[3][15:8] <= buffer_data_0[39:32];
        layer6[3][23:16] <= buffer_data_0[47:40];
        layer6[3][31:24] <= buffer_data_0[55:48];
        layer6[3][39:32] <= buffer_data_0[63:56];
        layer6[3][47:40] <= buffer_data_0[71:64];
        layer6[3][55:48] <= buffer_data_0[79:72];
        layer0[4][7:0] <= buffer_data_6[39:32];
        layer0[4][15:8] <= buffer_data_6[47:40];
        layer0[4][23:16] <= buffer_data_6[55:48];
        layer0[4][31:24] <= buffer_data_6[63:56];
        layer0[4][39:32] <= buffer_data_6[71:64];
        layer0[4][47:40] <= buffer_data_6[79:72];
        layer0[4][55:48] <= buffer_data_6[87:80];
        layer1[4][7:0] <= buffer_data_5[39:32];
        layer1[4][15:8] <= buffer_data_5[47:40];
        layer1[4][23:16] <= buffer_data_5[55:48];
        layer1[4][31:24] <= buffer_data_5[63:56];
        layer1[4][39:32] <= buffer_data_5[71:64];
        layer1[4][47:40] <= buffer_data_5[79:72];
        layer1[4][55:48] <= buffer_data_5[87:80];
        layer2[4][7:0] <= buffer_data_4[39:32];
        layer2[4][15:8] <= buffer_data_4[47:40];
        layer2[4][23:16] <= buffer_data_4[55:48];
        layer2[4][31:24] <= buffer_data_4[63:56];
        layer2[4][39:32] <= buffer_data_4[71:64];
        layer2[4][47:40] <= buffer_data_4[79:72];
        layer2[4][55:48] <= buffer_data_4[87:80];
        layer3[4][7:0] <= buffer_data_3[39:32];
        layer3[4][15:8] <= buffer_data_3[47:40];
        layer3[4][23:16] <= buffer_data_3[55:48];
        layer3[4][31:24] <= buffer_data_3[63:56];
        layer3[4][39:32] <= buffer_data_3[71:64];
        layer3[4][47:40] <= buffer_data_3[79:72];
        layer3[4][55:48] <= buffer_data_3[87:80];
        layer4[4][7:0] <= buffer_data_2[39:32];
        layer4[4][15:8] <= buffer_data_2[47:40];
        layer4[4][23:16] <= buffer_data_2[55:48];
        layer4[4][31:24] <= buffer_data_2[63:56];
        layer4[4][39:32] <= buffer_data_2[71:64];
        layer4[4][47:40] <= buffer_data_2[79:72];
        layer4[4][55:48] <= buffer_data_2[87:80];
        layer5[4][7:0] <= buffer_data_1[39:32];
        layer5[4][15:8] <= buffer_data_1[47:40];
        layer5[4][23:16] <= buffer_data_1[55:48];
        layer5[4][31:24] <= buffer_data_1[63:56];
        layer5[4][39:32] <= buffer_data_1[71:64];
        layer5[4][47:40] <= buffer_data_1[79:72];
        layer5[4][55:48] <= buffer_data_1[87:80];
        layer6[4][7:0] <= buffer_data_0[39:32];
        layer6[4][15:8] <= buffer_data_0[47:40];
        layer6[4][23:16] <= buffer_data_0[55:48];
        layer6[4][31:24] <= buffer_data_0[63:56];
        layer6[4][39:32] <= buffer_data_0[71:64];
        layer6[4][47:40] <= buffer_data_0[79:72];
        layer6[4][55:48] <= buffer_data_0[87:80];
        layer0[5][7:0] <= buffer_data_6[47:40];
        layer0[5][15:8] <= buffer_data_6[55:48];
        layer0[5][23:16] <= buffer_data_6[63:56];
        layer0[5][31:24] <= buffer_data_6[71:64];
        layer0[5][39:32] <= buffer_data_6[79:72];
        layer0[5][47:40] <= buffer_data_6[87:80];
        layer0[5][55:48] <= buffer_data_6[95:88];
        layer1[5][7:0] <= buffer_data_5[47:40];
        layer1[5][15:8] <= buffer_data_5[55:48];
        layer1[5][23:16] <= buffer_data_5[63:56];
        layer1[5][31:24] <= buffer_data_5[71:64];
        layer1[5][39:32] <= buffer_data_5[79:72];
        layer1[5][47:40] <= buffer_data_5[87:80];
        layer1[5][55:48] <= buffer_data_5[95:88];
        layer2[5][7:0] <= buffer_data_4[47:40];
        layer2[5][15:8] <= buffer_data_4[55:48];
        layer2[5][23:16] <= buffer_data_4[63:56];
        layer2[5][31:24] <= buffer_data_4[71:64];
        layer2[5][39:32] <= buffer_data_4[79:72];
        layer2[5][47:40] <= buffer_data_4[87:80];
        layer2[5][55:48] <= buffer_data_4[95:88];
        layer3[5][7:0] <= buffer_data_3[47:40];
        layer3[5][15:8] <= buffer_data_3[55:48];
        layer3[5][23:16] <= buffer_data_3[63:56];
        layer3[5][31:24] <= buffer_data_3[71:64];
        layer3[5][39:32] <= buffer_data_3[79:72];
        layer3[5][47:40] <= buffer_data_3[87:80];
        layer3[5][55:48] <= buffer_data_3[95:88];
        layer4[5][7:0] <= buffer_data_2[47:40];
        layer4[5][15:8] <= buffer_data_2[55:48];
        layer4[5][23:16] <= buffer_data_2[63:56];
        layer4[5][31:24] <= buffer_data_2[71:64];
        layer4[5][39:32] <= buffer_data_2[79:72];
        layer4[5][47:40] <= buffer_data_2[87:80];
        layer4[5][55:48] <= buffer_data_2[95:88];
        layer5[5][7:0] <= buffer_data_1[47:40];
        layer5[5][15:8] <= buffer_data_1[55:48];
        layer5[5][23:16] <= buffer_data_1[63:56];
        layer5[5][31:24] <= buffer_data_1[71:64];
        layer5[5][39:32] <= buffer_data_1[79:72];
        layer5[5][47:40] <= buffer_data_1[87:80];
        layer5[5][55:48] <= buffer_data_1[95:88];
        layer6[5][7:0] <= buffer_data_0[47:40];
        layer6[5][15:8] <= buffer_data_0[55:48];
        layer6[5][23:16] <= buffer_data_0[63:56];
        layer6[5][31:24] <= buffer_data_0[71:64];
        layer6[5][39:32] <= buffer_data_0[79:72];
        layer6[5][47:40] <= buffer_data_0[87:80];
        layer6[5][55:48] <= buffer_data_0[95:88];
        layer0[6][7:0] <= buffer_data_6[55:48];
        layer0[6][15:8] <= buffer_data_6[63:56];
        layer0[6][23:16] <= buffer_data_6[71:64];
        layer0[6][31:24] <= buffer_data_6[79:72];
        layer0[6][39:32] <= buffer_data_6[87:80];
        layer0[6][47:40] <= buffer_data_6[95:88];
        layer0[6][55:48] <= buffer_data_6[103:96];
        layer1[6][7:0] <= buffer_data_5[55:48];
        layer1[6][15:8] <= buffer_data_5[63:56];
        layer1[6][23:16] <= buffer_data_5[71:64];
        layer1[6][31:24] <= buffer_data_5[79:72];
        layer1[6][39:32] <= buffer_data_5[87:80];
        layer1[6][47:40] <= buffer_data_5[95:88];
        layer1[6][55:48] <= buffer_data_5[103:96];
        layer2[6][7:0] <= buffer_data_4[55:48];
        layer2[6][15:8] <= buffer_data_4[63:56];
        layer2[6][23:16] <= buffer_data_4[71:64];
        layer2[6][31:24] <= buffer_data_4[79:72];
        layer2[6][39:32] <= buffer_data_4[87:80];
        layer2[6][47:40] <= buffer_data_4[95:88];
        layer2[6][55:48] <= buffer_data_4[103:96];
        layer3[6][7:0] <= buffer_data_3[55:48];
        layer3[6][15:8] <= buffer_data_3[63:56];
        layer3[6][23:16] <= buffer_data_3[71:64];
        layer3[6][31:24] <= buffer_data_3[79:72];
        layer3[6][39:32] <= buffer_data_3[87:80];
        layer3[6][47:40] <= buffer_data_3[95:88];
        layer3[6][55:48] <= buffer_data_3[103:96];
        layer4[6][7:0] <= buffer_data_2[55:48];
        layer4[6][15:8] <= buffer_data_2[63:56];
        layer4[6][23:16] <= buffer_data_2[71:64];
        layer4[6][31:24] <= buffer_data_2[79:72];
        layer4[6][39:32] <= buffer_data_2[87:80];
        layer4[6][47:40] <= buffer_data_2[95:88];
        layer4[6][55:48] <= buffer_data_2[103:96];
        layer5[6][7:0] <= buffer_data_1[55:48];
        layer5[6][15:8] <= buffer_data_1[63:56];
        layer5[6][23:16] <= buffer_data_1[71:64];
        layer5[6][31:24] <= buffer_data_1[79:72];
        layer5[6][39:32] <= buffer_data_1[87:80];
        layer5[6][47:40] <= buffer_data_1[95:88];
        layer5[6][55:48] <= buffer_data_1[103:96];
        layer6[6][7:0] <= buffer_data_0[55:48];
        layer6[6][15:8] <= buffer_data_0[63:56];
        layer6[6][23:16] <= buffer_data_0[71:64];
        layer6[6][31:24] <= buffer_data_0[79:72];
        layer6[6][39:32] <= buffer_data_0[87:80];
        layer6[6][47:40] <= buffer_data_0[95:88];
        layer6[6][55:48] <= buffer_data_0[103:96];
        layer0[7][7:0] <= buffer_data_6[63:56];
        layer0[7][15:8] <= buffer_data_6[71:64];
        layer0[7][23:16] <= buffer_data_6[79:72];
        layer0[7][31:24] <= buffer_data_6[87:80];
        layer0[7][39:32] <= buffer_data_6[95:88];
        layer0[7][47:40] <= buffer_data_6[103:96];
        layer0[7][55:48] <= buffer_data_6[111:104];
        layer1[7][7:0] <= buffer_data_5[63:56];
        layer1[7][15:8] <= buffer_data_5[71:64];
        layer1[7][23:16] <= buffer_data_5[79:72];
        layer1[7][31:24] <= buffer_data_5[87:80];
        layer1[7][39:32] <= buffer_data_5[95:88];
        layer1[7][47:40] <= buffer_data_5[103:96];
        layer1[7][55:48] <= buffer_data_5[111:104];
        layer2[7][7:0] <= buffer_data_4[63:56];
        layer2[7][15:8] <= buffer_data_4[71:64];
        layer2[7][23:16] <= buffer_data_4[79:72];
        layer2[7][31:24] <= buffer_data_4[87:80];
        layer2[7][39:32] <= buffer_data_4[95:88];
        layer2[7][47:40] <= buffer_data_4[103:96];
        layer2[7][55:48] <= buffer_data_4[111:104];
        layer3[7][7:0] <= buffer_data_3[63:56];
        layer3[7][15:8] <= buffer_data_3[71:64];
        layer3[7][23:16] <= buffer_data_3[79:72];
        layer3[7][31:24] <= buffer_data_3[87:80];
        layer3[7][39:32] <= buffer_data_3[95:88];
        layer3[7][47:40] <= buffer_data_3[103:96];
        layer3[7][55:48] <= buffer_data_3[111:104];
        layer4[7][7:0] <= buffer_data_2[63:56];
        layer4[7][15:8] <= buffer_data_2[71:64];
        layer4[7][23:16] <= buffer_data_2[79:72];
        layer4[7][31:24] <= buffer_data_2[87:80];
        layer4[7][39:32] <= buffer_data_2[95:88];
        layer4[7][47:40] <= buffer_data_2[103:96];
        layer4[7][55:48] <= buffer_data_2[111:104];
        layer5[7][7:0] <= buffer_data_1[63:56];
        layer5[7][15:8] <= buffer_data_1[71:64];
        layer5[7][23:16] <= buffer_data_1[79:72];
        layer5[7][31:24] <= buffer_data_1[87:80];
        layer5[7][39:32] <= buffer_data_1[95:88];
        layer5[7][47:40] <= buffer_data_1[103:96];
        layer5[7][55:48] <= buffer_data_1[111:104];
        layer6[7][7:0] <= buffer_data_0[63:56];
        layer6[7][15:8] <= buffer_data_0[71:64];
        layer6[7][23:16] <= buffer_data_0[79:72];
        layer6[7][31:24] <= buffer_data_0[87:80];
        layer6[7][39:32] <= buffer_data_0[95:88];
        layer6[7][47:40] <= buffer_data_0[103:96];
        layer6[7][55:48] <= buffer_data_0[111:104];
        layer0[8][7:0] <= buffer_data_6[71:64];
        layer0[8][15:8] <= buffer_data_6[79:72];
        layer0[8][23:16] <= buffer_data_6[87:80];
        layer0[8][31:24] <= buffer_data_6[95:88];
        layer0[8][39:32] <= buffer_data_6[103:96];
        layer0[8][47:40] <= buffer_data_6[111:104];
        layer0[8][55:48] <= buffer_data_6[119:112];
        layer1[8][7:0] <= buffer_data_5[71:64];
        layer1[8][15:8] <= buffer_data_5[79:72];
        layer1[8][23:16] <= buffer_data_5[87:80];
        layer1[8][31:24] <= buffer_data_5[95:88];
        layer1[8][39:32] <= buffer_data_5[103:96];
        layer1[8][47:40] <= buffer_data_5[111:104];
        layer1[8][55:48] <= buffer_data_5[119:112];
        layer2[8][7:0] <= buffer_data_4[71:64];
        layer2[8][15:8] <= buffer_data_4[79:72];
        layer2[8][23:16] <= buffer_data_4[87:80];
        layer2[8][31:24] <= buffer_data_4[95:88];
        layer2[8][39:32] <= buffer_data_4[103:96];
        layer2[8][47:40] <= buffer_data_4[111:104];
        layer2[8][55:48] <= buffer_data_4[119:112];
        layer3[8][7:0] <= buffer_data_3[71:64];
        layer3[8][15:8] <= buffer_data_3[79:72];
        layer3[8][23:16] <= buffer_data_3[87:80];
        layer3[8][31:24] <= buffer_data_3[95:88];
        layer3[8][39:32] <= buffer_data_3[103:96];
        layer3[8][47:40] <= buffer_data_3[111:104];
        layer3[8][55:48] <= buffer_data_3[119:112];
        layer4[8][7:0] <= buffer_data_2[71:64];
        layer4[8][15:8] <= buffer_data_2[79:72];
        layer4[8][23:16] <= buffer_data_2[87:80];
        layer4[8][31:24] <= buffer_data_2[95:88];
        layer4[8][39:32] <= buffer_data_2[103:96];
        layer4[8][47:40] <= buffer_data_2[111:104];
        layer4[8][55:48] <= buffer_data_2[119:112];
        layer5[8][7:0] <= buffer_data_1[71:64];
        layer5[8][15:8] <= buffer_data_1[79:72];
        layer5[8][23:16] <= buffer_data_1[87:80];
        layer5[8][31:24] <= buffer_data_1[95:88];
        layer5[8][39:32] <= buffer_data_1[103:96];
        layer5[8][47:40] <= buffer_data_1[111:104];
        layer5[8][55:48] <= buffer_data_1[119:112];
        layer6[8][7:0] <= buffer_data_0[71:64];
        layer6[8][15:8] <= buffer_data_0[79:72];
        layer6[8][23:16] <= buffer_data_0[87:80];
        layer6[8][31:24] <= buffer_data_0[95:88];
        layer6[8][39:32] <= buffer_data_0[103:96];
        layer6[8][47:40] <= buffer_data_0[111:104];
        layer6[8][55:48] <= buffer_data_0[119:112];
        layer0[9][7:0] <= buffer_data_6[79:72];
        layer0[9][15:8] <= buffer_data_6[87:80];
        layer0[9][23:16] <= buffer_data_6[95:88];
        layer0[9][31:24] <= buffer_data_6[103:96];
        layer0[9][39:32] <= buffer_data_6[111:104];
        layer0[9][47:40] <= buffer_data_6[119:112];
        layer0[9][55:48] <= buffer_data_6[127:120];
        layer1[9][7:0] <= buffer_data_5[79:72];
        layer1[9][15:8] <= buffer_data_5[87:80];
        layer1[9][23:16] <= buffer_data_5[95:88];
        layer1[9][31:24] <= buffer_data_5[103:96];
        layer1[9][39:32] <= buffer_data_5[111:104];
        layer1[9][47:40] <= buffer_data_5[119:112];
        layer1[9][55:48] <= buffer_data_5[127:120];
        layer2[9][7:0] <= buffer_data_4[79:72];
        layer2[9][15:8] <= buffer_data_4[87:80];
        layer2[9][23:16] <= buffer_data_4[95:88];
        layer2[9][31:24] <= buffer_data_4[103:96];
        layer2[9][39:32] <= buffer_data_4[111:104];
        layer2[9][47:40] <= buffer_data_4[119:112];
        layer2[9][55:48] <= buffer_data_4[127:120];
        layer3[9][7:0] <= buffer_data_3[79:72];
        layer3[9][15:8] <= buffer_data_3[87:80];
        layer3[9][23:16] <= buffer_data_3[95:88];
        layer3[9][31:24] <= buffer_data_3[103:96];
        layer3[9][39:32] <= buffer_data_3[111:104];
        layer3[9][47:40] <= buffer_data_3[119:112];
        layer3[9][55:48] <= buffer_data_3[127:120];
        layer4[9][7:0] <= buffer_data_2[79:72];
        layer4[9][15:8] <= buffer_data_2[87:80];
        layer4[9][23:16] <= buffer_data_2[95:88];
        layer4[9][31:24] <= buffer_data_2[103:96];
        layer4[9][39:32] <= buffer_data_2[111:104];
        layer4[9][47:40] <= buffer_data_2[119:112];
        layer4[9][55:48] <= buffer_data_2[127:120];
        layer5[9][7:0] <= buffer_data_1[79:72];
        layer5[9][15:8] <= buffer_data_1[87:80];
        layer5[9][23:16] <= buffer_data_1[95:88];
        layer5[9][31:24] <= buffer_data_1[103:96];
        layer5[9][39:32] <= buffer_data_1[111:104];
        layer5[9][47:40] <= buffer_data_1[119:112];
        layer5[9][55:48] <= buffer_data_1[127:120];
        layer6[9][7:0] <= buffer_data_0[79:72];
        layer6[9][15:8] <= buffer_data_0[87:80];
        layer6[9][23:16] <= buffer_data_0[95:88];
        layer6[9][31:24] <= buffer_data_0[103:96];
        layer6[9][39:32] <= buffer_data_0[111:104];
        layer6[9][47:40] <= buffer_data_0[119:112];
        layer6[9][55:48] <= buffer_data_0[127:120];
        layer0[10][7:0] <= buffer_data_6[87:80];
        layer0[10][15:8] <= buffer_data_6[95:88];
        layer0[10][23:16] <= buffer_data_6[103:96];
        layer0[10][31:24] <= buffer_data_6[111:104];
        layer0[10][39:32] <= buffer_data_6[119:112];
        layer0[10][47:40] <= buffer_data_6[127:120];
        layer0[10][55:48] <= buffer_data_6[135:128];
        layer1[10][7:0] <= buffer_data_5[87:80];
        layer1[10][15:8] <= buffer_data_5[95:88];
        layer1[10][23:16] <= buffer_data_5[103:96];
        layer1[10][31:24] <= buffer_data_5[111:104];
        layer1[10][39:32] <= buffer_data_5[119:112];
        layer1[10][47:40] <= buffer_data_5[127:120];
        layer1[10][55:48] <= buffer_data_5[135:128];
        layer2[10][7:0] <= buffer_data_4[87:80];
        layer2[10][15:8] <= buffer_data_4[95:88];
        layer2[10][23:16] <= buffer_data_4[103:96];
        layer2[10][31:24] <= buffer_data_4[111:104];
        layer2[10][39:32] <= buffer_data_4[119:112];
        layer2[10][47:40] <= buffer_data_4[127:120];
        layer2[10][55:48] <= buffer_data_4[135:128];
        layer3[10][7:0] <= buffer_data_3[87:80];
        layer3[10][15:8] <= buffer_data_3[95:88];
        layer3[10][23:16] <= buffer_data_3[103:96];
        layer3[10][31:24] <= buffer_data_3[111:104];
        layer3[10][39:32] <= buffer_data_3[119:112];
        layer3[10][47:40] <= buffer_data_3[127:120];
        layer3[10][55:48] <= buffer_data_3[135:128];
        layer4[10][7:0] <= buffer_data_2[87:80];
        layer4[10][15:8] <= buffer_data_2[95:88];
        layer4[10][23:16] <= buffer_data_2[103:96];
        layer4[10][31:24] <= buffer_data_2[111:104];
        layer4[10][39:32] <= buffer_data_2[119:112];
        layer4[10][47:40] <= buffer_data_2[127:120];
        layer4[10][55:48] <= buffer_data_2[135:128];
        layer5[10][7:0] <= buffer_data_1[87:80];
        layer5[10][15:8] <= buffer_data_1[95:88];
        layer5[10][23:16] <= buffer_data_1[103:96];
        layer5[10][31:24] <= buffer_data_1[111:104];
        layer5[10][39:32] <= buffer_data_1[119:112];
        layer5[10][47:40] <= buffer_data_1[127:120];
        layer5[10][55:48] <= buffer_data_1[135:128];
        layer6[10][7:0] <= buffer_data_0[87:80];
        layer6[10][15:8] <= buffer_data_0[95:88];
        layer6[10][23:16] <= buffer_data_0[103:96];
        layer6[10][31:24] <= buffer_data_0[111:104];
        layer6[10][39:32] <= buffer_data_0[119:112];
        layer6[10][47:40] <= buffer_data_0[127:120];
        layer6[10][55:48] <= buffer_data_0[135:128];
        layer0[11][7:0] <= buffer_data_6[95:88];
        layer0[11][15:8] <= buffer_data_6[103:96];
        layer0[11][23:16] <= buffer_data_6[111:104];
        layer0[11][31:24] <= buffer_data_6[119:112];
        layer0[11][39:32] <= buffer_data_6[127:120];
        layer0[11][47:40] <= buffer_data_6[135:128];
        layer0[11][55:48] <= buffer_data_6[143:136];
        layer1[11][7:0] <= buffer_data_5[95:88];
        layer1[11][15:8] <= buffer_data_5[103:96];
        layer1[11][23:16] <= buffer_data_5[111:104];
        layer1[11][31:24] <= buffer_data_5[119:112];
        layer1[11][39:32] <= buffer_data_5[127:120];
        layer1[11][47:40] <= buffer_data_5[135:128];
        layer1[11][55:48] <= buffer_data_5[143:136];
        layer2[11][7:0] <= buffer_data_4[95:88];
        layer2[11][15:8] <= buffer_data_4[103:96];
        layer2[11][23:16] <= buffer_data_4[111:104];
        layer2[11][31:24] <= buffer_data_4[119:112];
        layer2[11][39:32] <= buffer_data_4[127:120];
        layer2[11][47:40] <= buffer_data_4[135:128];
        layer2[11][55:48] <= buffer_data_4[143:136];
        layer3[11][7:0] <= buffer_data_3[95:88];
        layer3[11][15:8] <= buffer_data_3[103:96];
        layer3[11][23:16] <= buffer_data_3[111:104];
        layer3[11][31:24] <= buffer_data_3[119:112];
        layer3[11][39:32] <= buffer_data_3[127:120];
        layer3[11][47:40] <= buffer_data_3[135:128];
        layer3[11][55:48] <= buffer_data_3[143:136];
        layer4[11][7:0] <= buffer_data_2[95:88];
        layer4[11][15:8] <= buffer_data_2[103:96];
        layer4[11][23:16] <= buffer_data_2[111:104];
        layer4[11][31:24] <= buffer_data_2[119:112];
        layer4[11][39:32] <= buffer_data_2[127:120];
        layer4[11][47:40] <= buffer_data_2[135:128];
        layer4[11][55:48] <= buffer_data_2[143:136];
        layer5[11][7:0] <= buffer_data_1[95:88];
        layer5[11][15:8] <= buffer_data_1[103:96];
        layer5[11][23:16] <= buffer_data_1[111:104];
        layer5[11][31:24] <= buffer_data_1[119:112];
        layer5[11][39:32] <= buffer_data_1[127:120];
        layer5[11][47:40] <= buffer_data_1[135:128];
        layer5[11][55:48] <= buffer_data_1[143:136];
        layer6[11][7:0] <= buffer_data_0[95:88];
        layer6[11][15:8] <= buffer_data_0[103:96];
        layer6[11][23:16] <= buffer_data_0[111:104];
        layer6[11][31:24] <= buffer_data_0[119:112];
        layer6[11][39:32] <= buffer_data_0[127:120];
        layer6[11][47:40] <= buffer_data_0[135:128];
        layer6[11][55:48] <= buffer_data_0[143:136];
        layer0[12][7:0] <= buffer_data_6[103:96];
        layer0[12][15:8] <= buffer_data_6[111:104];
        layer0[12][23:16] <= buffer_data_6[119:112];
        layer0[12][31:24] <= buffer_data_6[127:120];
        layer0[12][39:32] <= buffer_data_6[135:128];
        layer0[12][47:40] <= buffer_data_6[143:136];
        layer0[12][55:48] <= buffer_data_6[151:144];
        layer1[12][7:0] <= buffer_data_5[103:96];
        layer1[12][15:8] <= buffer_data_5[111:104];
        layer1[12][23:16] <= buffer_data_5[119:112];
        layer1[12][31:24] <= buffer_data_5[127:120];
        layer1[12][39:32] <= buffer_data_5[135:128];
        layer1[12][47:40] <= buffer_data_5[143:136];
        layer1[12][55:48] <= buffer_data_5[151:144];
        layer2[12][7:0] <= buffer_data_4[103:96];
        layer2[12][15:8] <= buffer_data_4[111:104];
        layer2[12][23:16] <= buffer_data_4[119:112];
        layer2[12][31:24] <= buffer_data_4[127:120];
        layer2[12][39:32] <= buffer_data_4[135:128];
        layer2[12][47:40] <= buffer_data_4[143:136];
        layer2[12][55:48] <= buffer_data_4[151:144];
        layer3[12][7:0] <= buffer_data_3[103:96];
        layer3[12][15:8] <= buffer_data_3[111:104];
        layer3[12][23:16] <= buffer_data_3[119:112];
        layer3[12][31:24] <= buffer_data_3[127:120];
        layer3[12][39:32] <= buffer_data_3[135:128];
        layer3[12][47:40] <= buffer_data_3[143:136];
        layer3[12][55:48] <= buffer_data_3[151:144];
        layer4[12][7:0] <= buffer_data_2[103:96];
        layer4[12][15:8] <= buffer_data_2[111:104];
        layer4[12][23:16] <= buffer_data_2[119:112];
        layer4[12][31:24] <= buffer_data_2[127:120];
        layer4[12][39:32] <= buffer_data_2[135:128];
        layer4[12][47:40] <= buffer_data_2[143:136];
        layer4[12][55:48] <= buffer_data_2[151:144];
        layer5[12][7:0] <= buffer_data_1[103:96];
        layer5[12][15:8] <= buffer_data_1[111:104];
        layer5[12][23:16] <= buffer_data_1[119:112];
        layer5[12][31:24] <= buffer_data_1[127:120];
        layer5[12][39:32] <= buffer_data_1[135:128];
        layer5[12][47:40] <= buffer_data_1[143:136];
        layer5[12][55:48] <= buffer_data_1[151:144];
        layer6[12][7:0] <= buffer_data_0[103:96];
        layer6[12][15:8] <= buffer_data_0[111:104];
        layer6[12][23:16] <= buffer_data_0[119:112];
        layer6[12][31:24] <= buffer_data_0[127:120];
        layer6[12][39:32] <= buffer_data_0[135:128];
        layer6[12][47:40] <= buffer_data_0[143:136];
        layer6[12][55:48] <= buffer_data_0[151:144];
        layer0[13][7:0] <= buffer_data_6[111:104];
        layer0[13][15:8] <= buffer_data_6[119:112];
        layer0[13][23:16] <= buffer_data_6[127:120];
        layer0[13][31:24] <= buffer_data_6[135:128];
        layer0[13][39:32] <= buffer_data_6[143:136];
        layer0[13][47:40] <= buffer_data_6[151:144];
        layer0[13][55:48] <= 0;
        layer1[13][7:0] <= buffer_data_5[111:104];
        layer1[13][15:8] <= buffer_data_5[119:112];
        layer1[13][23:16] <= buffer_data_5[127:120];
        layer1[13][31:24] <= buffer_data_5[135:128];
        layer1[13][39:32] <= buffer_data_5[143:136];
        layer1[13][47:40] <= buffer_data_5[151:144];
        layer1[13][55:48] <= 0;
        layer2[13][7:0] <= buffer_data_4[111:104];
        layer2[13][15:8] <= buffer_data_4[119:112];
        layer2[13][23:16] <= buffer_data_4[127:120];
        layer2[13][31:24] <= buffer_data_4[135:128];
        layer2[13][39:32] <= buffer_data_4[143:136];
        layer2[13][47:40] <= buffer_data_4[151:144];
        layer2[13][55:48] <= 0;
        layer3[13][7:0] <= buffer_data_3[111:104];
        layer3[13][15:8] <= buffer_data_3[119:112];
        layer3[13][23:16] <= buffer_data_3[127:120];
        layer3[13][31:24] <= buffer_data_3[135:128];
        layer3[13][39:32] <= buffer_data_3[143:136];
        layer3[13][47:40] <= buffer_data_3[151:144];
        layer3[13][55:48] <= 0;
        layer4[13][7:0] <= buffer_data_2[111:104];
        layer4[13][15:8] <= buffer_data_2[119:112];
        layer4[13][23:16] <= buffer_data_2[127:120];
        layer4[13][31:24] <= buffer_data_2[135:128];
        layer4[13][39:32] <= buffer_data_2[143:136];
        layer4[13][47:40] <= buffer_data_2[151:144];
        layer4[13][55:48] <= 0;
        layer5[13][7:0] <= buffer_data_1[111:104];
        layer5[13][15:8] <= buffer_data_1[119:112];
        layer5[13][23:16] <= buffer_data_1[127:120];
        layer5[13][31:24] <= buffer_data_1[135:128];
        layer5[13][39:32] <= buffer_data_1[143:136];
        layer5[13][47:40] <= buffer_data_1[151:144];
        layer5[13][55:48] <= 0;
        layer6[13][7:0] <= buffer_data_0[111:104];
        layer6[13][15:8] <= buffer_data_0[119:112];
        layer6[13][23:16] <= buffer_data_0[127:120];
        layer6[13][31:24] <= buffer_data_0[135:128];
        layer6[13][39:32] <= buffer_data_0[143:136];
        layer6[13][47:40] <= buffer_data_0[151:144];
        layer6[13][55:48] <= 0;
        layer0[14][7:0] <= buffer_data_6[119:112];
        layer0[14][15:8] <= buffer_data_6[127:120];
        layer0[14][23:16] <= buffer_data_6[135:128];
        layer0[14][31:24] <= buffer_data_6[143:136];
        layer0[14][39:32] <= buffer_data_6[151:144];
        layer0[14][47:40] <= 0;
        layer0[14][55:48] <= 0;
        layer1[14][7:0] <= buffer_data_5[119:112];
        layer1[14][15:8] <= buffer_data_5[127:120];
        layer1[14][23:16] <= buffer_data_5[135:128];
        layer1[14][31:24] <= buffer_data_5[143:136];
        layer1[14][39:32] <= buffer_data_5[151:144];
        layer1[14][47:40] <= 0;
        layer1[14][55:48] <= 0;
        layer2[14][7:0] <= buffer_data_4[119:112];
        layer2[14][15:8] <= buffer_data_4[127:120];
        layer2[14][23:16] <= buffer_data_4[135:128];
        layer2[14][31:24] <= buffer_data_4[143:136];
        layer2[14][39:32] <= buffer_data_4[151:144];
        layer2[14][47:40] <= 0;
        layer2[14][55:48] <= 0;
        layer3[14][7:0] <= buffer_data_3[119:112];
        layer3[14][15:8] <= buffer_data_3[127:120];
        layer3[14][23:16] <= buffer_data_3[135:128];
        layer3[14][31:24] <= buffer_data_3[143:136];
        layer3[14][39:32] <= buffer_data_3[151:144];
        layer3[14][47:40] <= 0;
        layer3[14][55:48] <= 0;
        layer4[14][7:0] <= buffer_data_2[119:112];
        layer4[14][15:8] <= buffer_data_2[127:120];
        layer4[14][23:16] <= buffer_data_2[135:128];
        layer4[14][31:24] <= buffer_data_2[143:136];
        layer4[14][39:32] <= buffer_data_2[151:144];
        layer4[14][47:40] <= 0;
        layer4[14][55:48] <= 0;
        layer5[14][7:0] <= buffer_data_1[119:112];
        layer5[14][15:8] <= buffer_data_1[127:120];
        layer5[14][23:16] <= buffer_data_1[135:128];
        layer5[14][31:24] <= buffer_data_1[143:136];
        layer5[14][39:32] <= buffer_data_1[151:144];
        layer5[14][47:40] <= 0;
        layer5[14][55:48] <= 0;
        layer6[14][7:0] <= buffer_data_0[119:112];
        layer6[14][15:8] <= buffer_data_0[127:120];
        layer6[14][23:16] <= buffer_data_0[135:128];
        layer6[14][31:24] <= buffer_data_0[143:136];
        layer6[14][39:32] <= buffer_data_0[151:144];
        layer6[14][47:40] <= 0;
        layer6[14][55:48] <= 0;
        layer0[15][7:0] <= buffer_data_6[127:120];
        layer0[15][15:8] <= buffer_data_6[135:128];
        layer0[15][23:16] <= buffer_data_6[143:136];
        layer0[15][31:24] <= buffer_data_6[151:144];
        layer0[15][39:32] <= 0;
        layer0[15][47:40] <= 0;
        layer0[15][55:48] <= 0;
        layer1[15][7:0] <= buffer_data_5[127:120];
        layer1[15][15:8] <= buffer_data_5[135:128];
        layer1[15][23:16] <= buffer_data_5[143:136];
        layer1[15][31:24] <= buffer_data_5[151:144];
        layer1[15][39:32] <= 0;
        layer1[15][47:40] <= 0;
        layer1[15][55:48] <= 0;
        layer2[15][7:0] <= buffer_data_4[127:120];
        layer2[15][15:8] <= buffer_data_4[135:128];
        layer2[15][23:16] <= buffer_data_4[143:136];
        layer2[15][31:24] <= buffer_data_4[151:144];
        layer2[15][39:32] <= 0;
        layer2[15][47:40] <= 0;
        layer2[15][55:48] <= 0;
        layer3[15][7:0] <= buffer_data_3[127:120];
        layer3[15][15:8] <= buffer_data_3[135:128];
        layer3[15][23:16] <= buffer_data_3[143:136];
        layer3[15][31:24] <= buffer_data_3[151:144];
        layer3[15][39:32] <= 0;
        layer3[15][47:40] <= 0;
        layer3[15][55:48] <= 0;
        layer4[15][7:0] <= buffer_data_2[127:120];
        layer4[15][15:8] <= buffer_data_2[135:128];
        layer4[15][23:16] <= buffer_data_2[143:136];
        layer4[15][31:24] <= buffer_data_2[151:144];
        layer4[15][39:32] <= 0;
        layer4[15][47:40] <= 0;
        layer4[15][55:48] <= 0;
        layer5[15][7:0] <= buffer_data_1[127:120];
        layer5[15][15:8] <= buffer_data_1[135:128];
        layer5[15][23:16] <= buffer_data_1[143:136];
        layer5[15][31:24] <= buffer_data_1[151:144];
        layer5[15][39:32] <= 0;
        layer5[15][47:40] <= 0;
        layer5[15][55:48] <= 0;
        layer6[15][7:0] <= buffer_data_0[127:120];
        layer6[15][15:8] <= buffer_data_0[135:128];
        layer6[15][23:16] <= buffer_data_0[143:136];
        layer6[15][31:24] <= buffer_data_0[151:144];
        layer6[15][39:32] <= 0;
        layer6[15][47:40] <= 0;
        layer6[15][55:48] <= 0;
    end
      default: begin
        layer0[0][7:0] <= 'd0;
        layer0[0][15:8] <= 'd0;
        layer0[0][23:16] <= 'd0;
        layer0[0][31:24] <= 'd0;
        layer0[0][39:32] <= 'd0;
        layer0[0][47:40] <= 'd0;
        layer0[0][55:48] <= 'd0;
        layer1[0][7:0] <= 'd0;
        layer1[0][15:8] <= 'd0;
        layer1[0][23:16] <= 'd0;
        layer1[0][31:24] <= 'd0;
        layer1[0][39:32] <= 'd0;
        layer1[0][47:40] <= 'd0;
        layer1[0][55:48] <= 'd0;
        layer2[0][7:0] <= 'd0;
        layer2[0][15:8] <= 'd0;
        layer2[0][23:16] <= 'd0;
        layer2[0][31:24] <= 'd0;
        layer2[0][39:32] <= 'd0;
        layer2[0][47:40] <= 'd0;
        layer2[0][55:48] <= 'd0;
        layer3[0][7:0] <= 'd0;
        layer3[0][15:8] <= 'd0;
        layer3[0][23:16] <= 'd0;
        layer3[0][31:24] <= 'd0;
        layer3[0][39:32] <= 'd0;
        layer3[0][47:40] <= 'd0;
        layer3[0][55:48] <= 'd0;
        layer4[0][7:0] <= 'd0;
        layer4[0][15:8] <= 'd0;
        layer4[0][23:16] <= 'd0;
        layer4[0][31:24] <= 'd0;
        layer4[0][39:32] <= 'd0;
        layer4[0][47:40] <= 'd0;
        layer4[0][55:48] <= 'd0;
        layer5[0][7:0] <= 'd0;
        layer5[0][15:8] <= 'd0;
        layer5[0][23:16] <= 'd0;
        layer5[0][31:24] <= 'd0;
        layer5[0][39:32] <= 'd0;
        layer5[0][47:40] <= 'd0;
        layer5[0][55:48] <= 'd0;
        layer6[0][7:0] <= 'd0;
        layer6[0][15:8] <= 'd0;
        layer6[0][23:16] <= 'd0;
        layer6[0][31:24] <= 'd0;
        layer6[0][39:32] <= 'd0;
        layer6[0][47:40] <= 'd0;
        layer6[0][55:48] <= 'd0;
        layer0[1][7:0] <= 'd0;
        layer0[1][15:8] <= 'd0;
        layer0[1][23:16] <= 'd0;
        layer0[1][31:24] <= 'd0;
        layer0[1][39:32] <= 'd0;
        layer0[1][47:40] <= 'd0;
        layer0[1][55:48] <= 'd0;
        layer1[1][7:0] <= 'd0;
        layer1[1][15:8] <= 'd0;
        layer1[1][23:16] <= 'd0;
        layer1[1][31:24] <= 'd0;
        layer1[1][39:32] <= 'd0;
        layer1[1][47:40] <= 'd0;
        layer1[1][55:48] <= 'd0;
        layer2[1][7:0] <= 'd0;
        layer2[1][15:8] <= 'd0;
        layer2[1][23:16] <= 'd0;
        layer2[1][31:24] <= 'd0;
        layer2[1][39:32] <= 'd0;
        layer2[1][47:40] <= 'd0;
        layer2[1][55:48] <= 'd0;
        layer3[1][7:0] <= 'd0;
        layer3[1][15:8] <= 'd0;
        layer3[1][23:16] <= 'd0;
        layer3[1][31:24] <= 'd0;
        layer3[1][39:32] <= 'd0;
        layer3[1][47:40] <= 'd0;
        layer3[1][55:48] <= 'd0;
        layer4[1][7:0] <= 'd0;
        layer4[1][15:8] <= 'd0;
        layer4[1][23:16] <= 'd0;
        layer4[1][31:24] <= 'd0;
        layer4[1][39:32] <= 'd0;
        layer4[1][47:40] <= 'd0;
        layer4[1][55:48] <= 'd0;
        layer5[1][7:0] <= 'd0;
        layer5[1][15:8] <= 'd0;
        layer5[1][23:16] <= 'd0;
        layer5[1][31:24] <= 'd0;
        layer5[1][39:32] <= 'd0;
        layer5[1][47:40] <= 'd0;
        layer5[1][55:48] <= 'd0;
        layer6[1][7:0] <= 'd0;
        layer6[1][15:8] <= 'd0;
        layer6[1][23:16] <= 'd0;
        layer6[1][31:24] <= 'd0;
        layer6[1][39:32] <= 'd0;
        layer6[1][47:40] <= 'd0;
        layer6[1][55:48] <= 'd0;
        layer0[2][7:0] <= 'd0;
        layer0[2][15:8] <= 'd0;
        layer0[2][23:16] <= 'd0;
        layer0[2][31:24] <= 'd0;
        layer0[2][39:32] <= 'd0;
        layer0[2][47:40] <= 'd0;
        layer0[2][55:48] <= 'd0;
        layer1[2][7:0] <= 'd0;
        layer1[2][15:8] <= 'd0;
        layer1[2][23:16] <= 'd0;
        layer1[2][31:24] <= 'd0;
        layer1[2][39:32] <= 'd0;
        layer1[2][47:40] <= 'd0;
        layer1[2][55:48] <= 'd0;
        layer2[2][7:0] <= 'd0;
        layer2[2][15:8] <= 'd0;
        layer2[2][23:16] <= 'd0;
        layer2[2][31:24] <= 'd0;
        layer2[2][39:32] <= 'd0;
        layer2[2][47:40] <= 'd0;
        layer2[2][55:48] <= 'd0;
        layer3[2][7:0] <= 'd0;
        layer3[2][15:8] <= 'd0;
        layer3[2][23:16] <= 'd0;
        layer3[2][31:24] <= 'd0;
        layer3[2][39:32] <= 'd0;
        layer3[2][47:40] <= 'd0;
        layer3[2][55:48] <= 'd0;
        layer4[2][7:0] <= 'd0;
        layer4[2][15:8] <= 'd0;
        layer4[2][23:16] <= 'd0;
        layer4[2][31:24] <= 'd0;
        layer4[2][39:32] <= 'd0;
        layer4[2][47:40] <= 'd0;
        layer4[2][55:48] <= 'd0;
        layer5[2][7:0] <= 'd0;
        layer5[2][15:8] <= 'd0;
        layer5[2][23:16] <= 'd0;
        layer5[2][31:24] <= 'd0;
        layer5[2][39:32] <= 'd0;
        layer5[2][47:40] <= 'd0;
        layer5[2][55:48] <= 'd0;
        layer6[2][7:0] <= 'd0;
        layer6[2][15:8] <= 'd0;
        layer6[2][23:16] <= 'd0;
        layer6[2][31:24] <= 'd0;
        layer6[2][39:32] <= 'd0;
        layer6[2][47:40] <= 'd0;
        layer6[2][55:48] <= 'd0;
        layer0[3][7:0] <= 'd0;
        layer0[3][15:8] <= 'd0;
        layer0[3][23:16] <= 'd0;
        layer0[3][31:24] <= 'd0;
        layer0[3][39:32] <= 'd0;
        layer0[3][47:40] <= 'd0;
        layer0[3][55:48] <= 'd0;
        layer1[3][7:0] <= 'd0;
        layer1[3][15:8] <= 'd0;
        layer1[3][23:16] <= 'd0;
        layer1[3][31:24] <= 'd0;
        layer1[3][39:32] <= 'd0;
        layer1[3][47:40] <= 'd0;
        layer1[3][55:48] <= 'd0;
        layer2[3][7:0] <= 'd0;
        layer2[3][15:8] <= 'd0;
        layer2[3][23:16] <= 'd0;
        layer2[3][31:24] <= 'd0;
        layer2[3][39:32] <= 'd0;
        layer2[3][47:40] <= 'd0;
        layer2[3][55:48] <= 'd0;
        layer3[3][7:0] <= 'd0;
        layer3[3][15:8] <= 'd0;
        layer3[3][23:16] <= 'd0;
        layer3[3][31:24] <= 'd0;
        layer3[3][39:32] <= 'd0;
        layer3[3][47:40] <= 'd0;
        layer3[3][55:48] <= 'd0;
        layer4[3][7:0] <= 'd0;
        layer4[3][15:8] <= 'd0;
        layer4[3][23:16] <= 'd0;
        layer4[3][31:24] <= 'd0;
        layer4[3][39:32] <= 'd0;
        layer4[3][47:40] <= 'd0;
        layer4[3][55:48] <= 'd0;
        layer5[3][7:0] <= 'd0;
        layer5[3][15:8] <= 'd0;
        layer5[3][23:16] <= 'd0;
        layer5[3][31:24] <= 'd0;
        layer5[3][39:32] <= 'd0;
        layer5[3][47:40] <= 'd0;
        layer5[3][55:48] <= 'd0;
        layer6[3][7:0] <= 'd0;
        layer6[3][15:8] <= 'd0;
        layer6[3][23:16] <= 'd0;
        layer6[3][31:24] <= 'd0;
        layer6[3][39:32] <= 'd0;
        layer6[3][47:40] <= 'd0;
        layer6[3][55:48] <= 'd0;
        layer0[4][7:0] <= 'd0;
        layer0[4][15:8] <= 'd0;
        layer0[4][23:16] <= 'd0;
        layer0[4][31:24] <= 'd0;
        layer0[4][39:32] <= 'd0;
        layer0[4][47:40] <= 'd0;
        layer0[4][55:48] <= 'd0;
        layer1[4][7:0] <= 'd0;
        layer1[4][15:8] <= 'd0;
        layer1[4][23:16] <= 'd0;
        layer1[4][31:24] <= 'd0;
        layer1[4][39:32] <= 'd0;
        layer1[4][47:40] <= 'd0;
        layer1[4][55:48] <= 'd0;
        layer2[4][7:0] <= 'd0;
        layer2[4][15:8] <= 'd0;
        layer2[4][23:16] <= 'd0;
        layer2[4][31:24] <= 'd0;
        layer2[4][39:32] <= 'd0;
        layer2[4][47:40] <= 'd0;
        layer2[4][55:48] <= 'd0;
        layer3[4][7:0] <= 'd0;
        layer3[4][15:8] <= 'd0;
        layer3[4][23:16] <= 'd0;
        layer3[4][31:24] <= 'd0;
        layer3[4][39:32] <= 'd0;
        layer3[4][47:40] <= 'd0;
        layer3[4][55:48] <= 'd0;
        layer4[4][7:0] <= 'd0;
        layer4[4][15:8] <= 'd0;
        layer4[4][23:16] <= 'd0;
        layer4[4][31:24] <= 'd0;
        layer4[4][39:32] <= 'd0;
        layer4[4][47:40] <= 'd0;
        layer4[4][55:48] <= 'd0;
        layer5[4][7:0] <= 'd0;
        layer5[4][15:8] <= 'd0;
        layer5[4][23:16] <= 'd0;
        layer5[4][31:24] <= 'd0;
        layer5[4][39:32] <= 'd0;
        layer5[4][47:40] <= 'd0;
        layer5[4][55:48] <= 'd0;
        layer6[4][7:0] <= 'd0;
        layer6[4][15:8] <= 'd0;
        layer6[4][23:16] <= 'd0;
        layer6[4][31:24] <= 'd0;
        layer6[4][39:32] <= 'd0;
        layer6[4][47:40] <= 'd0;
        layer6[4][55:48] <= 'd0;
        layer0[5][7:0] <= 'd0;
        layer0[5][15:8] <= 'd0;
        layer0[5][23:16] <= 'd0;
        layer0[5][31:24] <= 'd0;
        layer0[5][39:32] <= 'd0;
        layer0[5][47:40] <= 'd0;
        layer0[5][55:48] <= 'd0;
        layer1[5][7:0] <= 'd0;
        layer1[5][15:8] <= 'd0;
        layer1[5][23:16] <= 'd0;
        layer1[5][31:24] <= 'd0;
        layer1[5][39:32] <= 'd0;
        layer1[5][47:40] <= 'd0;
        layer1[5][55:48] <= 'd0;
        layer2[5][7:0] <= 'd0;
        layer2[5][15:8] <= 'd0;
        layer2[5][23:16] <= 'd0;
        layer2[5][31:24] <= 'd0;
        layer2[5][39:32] <= 'd0;
        layer2[5][47:40] <= 'd0;
        layer2[5][55:48] <= 'd0;
        layer3[5][7:0] <= 'd0;
        layer3[5][15:8] <= 'd0;
        layer3[5][23:16] <= 'd0;
        layer3[5][31:24] <= 'd0;
        layer3[5][39:32] <= 'd0;
        layer3[5][47:40] <= 'd0;
        layer3[5][55:48] <= 'd0;
        layer4[5][7:0] <= 'd0;
        layer4[5][15:8] <= 'd0;
        layer4[5][23:16] <= 'd0;
        layer4[5][31:24] <= 'd0;
        layer4[5][39:32] <= 'd0;
        layer4[5][47:40] <= 'd0;
        layer4[5][55:48] <= 'd0;
        layer5[5][7:0] <= 'd0;
        layer5[5][15:8] <= 'd0;
        layer5[5][23:16] <= 'd0;
        layer5[5][31:24] <= 'd0;
        layer5[5][39:32] <= 'd0;
        layer5[5][47:40] <= 'd0;
        layer5[5][55:48] <= 'd0;
        layer6[5][7:0] <= 'd0;
        layer6[5][15:8] <= 'd0;
        layer6[5][23:16] <= 'd0;
        layer6[5][31:24] <= 'd0;
        layer6[5][39:32] <= 'd0;
        layer6[5][47:40] <= 'd0;
        layer6[5][55:48] <= 'd0;
        layer0[6][7:0] <= 'd0;
        layer0[6][15:8] <= 'd0;
        layer0[6][23:16] <= 'd0;
        layer0[6][31:24] <= 'd0;
        layer0[6][39:32] <= 'd0;
        layer0[6][47:40] <= 'd0;
        layer0[6][55:48] <= 'd0;
        layer1[6][7:0] <= 'd0;
        layer1[6][15:8] <= 'd0;
        layer1[6][23:16] <= 'd0;
        layer1[6][31:24] <= 'd0;
        layer1[6][39:32] <= 'd0;
        layer1[6][47:40] <= 'd0;
        layer1[6][55:48] <= 'd0;
        layer2[6][7:0] <= 'd0;
        layer2[6][15:8] <= 'd0;
        layer2[6][23:16] <= 'd0;
        layer2[6][31:24] <= 'd0;
        layer2[6][39:32] <= 'd0;
        layer2[6][47:40] <= 'd0;
        layer2[6][55:48] <= 'd0;
        layer3[6][7:0] <= 'd0;
        layer3[6][15:8] <= 'd0;
        layer3[6][23:16] <= 'd0;
        layer3[6][31:24] <= 'd0;
        layer3[6][39:32] <= 'd0;
        layer3[6][47:40] <= 'd0;
        layer3[6][55:48] <= 'd0;
        layer4[6][7:0] <= 'd0;
        layer4[6][15:8] <= 'd0;
        layer4[6][23:16] <= 'd0;
        layer4[6][31:24] <= 'd0;
        layer4[6][39:32] <= 'd0;
        layer4[6][47:40] <= 'd0;
        layer4[6][55:48] <= 'd0;
        layer5[6][7:0] <= 'd0;
        layer5[6][15:8] <= 'd0;
        layer5[6][23:16] <= 'd0;
        layer5[6][31:24] <= 'd0;
        layer5[6][39:32] <= 'd0;
        layer5[6][47:40] <= 'd0;
        layer5[6][55:48] <= 'd0;
        layer6[6][7:0] <= 'd0;
        layer6[6][15:8] <= 'd0;
        layer6[6][23:16] <= 'd0;
        layer6[6][31:24] <= 'd0;
        layer6[6][39:32] <= 'd0;
        layer6[6][47:40] <= 'd0;
        layer6[6][55:48] <= 'd0;
        layer0[7][7:0] <= 'd0;
        layer0[7][15:8] <= 'd0;
        layer0[7][23:16] <= 'd0;
        layer0[7][31:24] <= 'd0;
        layer0[7][39:32] <= 'd0;
        layer0[7][47:40] <= 'd0;
        layer0[7][55:48] <= 'd0;
        layer1[7][7:0] <= 'd0;
        layer1[7][15:8] <= 'd0;
        layer1[7][23:16] <= 'd0;
        layer1[7][31:24] <= 'd0;
        layer1[7][39:32] <= 'd0;
        layer1[7][47:40] <= 'd0;
        layer1[7][55:48] <= 'd0;
        layer2[7][7:0] <= 'd0;
        layer2[7][15:8] <= 'd0;
        layer2[7][23:16] <= 'd0;
        layer2[7][31:24] <= 'd0;
        layer2[7][39:32] <= 'd0;
        layer2[7][47:40] <= 'd0;
        layer2[7][55:48] <= 'd0;
        layer3[7][7:0] <= 'd0;
        layer3[7][15:8] <= 'd0;
        layer3[7][23:16] <= 'd0;
        layer3[7][31:24] <= 'd0;
        layer3[7][39:32] <= 'd0;
        layer3[7][47:40] <= 'd0;
        layer3[7][55:48] <= 'd0;
        layer4[7][7:0] <= 'd0;
        layer4[7][15:8] <= 'd0;
        layer4[7][23:16] <= 'd0;
        layer4[7][31:24] <= 'd0;
        layer4[7][39:32] <= 'd0;
        layer4[7][47:40] <= 'd0;
        layer4[7][55:48] <= 'd0;
        layer5[7][7:0] <= 'd0;
        layer5[7][15:8] <= 'd0;
        layer5[7][23:16] <= 'd0;
        layer5[7][31:24] <= 'd0;
        layer5[7][39:32] <= 'd0;
        layer5[7][47:40] <= 'd0;
        layer5[7][55:48] <= 'd0;
        layer6[7][7:0] <= 'd0;
        layer6[7][15:8] <= 'd0;
        layer6[7][23:16] <= 'd0;
        layer6[7][31:24] <= 'd0;
        layer6[7][39:32] <= 'd0;
        layer6[7][47:40] <= 'd0;
        layer6[7][55:48] <= 'd0;
        layer0[8][7:0] <= 'd0;
        layer0[8][15:8] <= 'd0;
        layer0[8][23:16] <= 'd0;
        layer0[8][31:24] <= 'd0;
        layer0[8][39:32] <= 'd0;
        layer0[8][47:40] <= 'd0;
        layer0[8][55:48] <= 'd0;
        layer1[8][7:0] <= 'd0;
        layer1[8][15:8] <= 'd0;
        layer1[8][23:16] <= 'd0;
        layer1[8][31:24] <= 'd0;
        layer1[8][39:32] <= 'd0;
        layer1[8][47:40] <= 'd0;
        layer1[8][55:48] <= 'd0;
        layer2[8][7:0] <= 'd0;
        layer2[8][15:8] <= 'd0;
        layer2[8][23:16] <= 'd0;
        layer2[8][31:24] <= 'd0;
        layer2[8][39:32] <= 'd0;
        layer2[8][47:40] <= 'd0;
        layer2[8][55:48] <= 'd0;
        layer3[8][7:0] <= 'd0;
        layer3[8][15:8] <= 'd0;
        layer3[8][23:16] <= 'd0;
        layer3[8][31:24] <= 'd0;
        layer3[8][39:32] <= 'd0;
        layer3[8][47:40] <= 'd0;
        layer3[8][55:48] <= 'd0;
        layer4[8][7:0] <= 'd0;
        layer4[8][15:8] <= 'd0;
        layer4[8][23:16] <= 'd0;
        layer4[8][31:24] <= 'd0;
        layer4[8][39:32] <= 'd0;
        layer4[8][47:40] <= 'd0;
        layer4[8][55:48] <= 'd0;
        layer5[8][7:0] <= 'd0;
        layer5[8][15:8] <= 'd0;
        layer5[8][23:16] <= 'd0;
        layer5[8][31:24] <= 'd0;
        layer5[8][39:32] <= 'd0;
        layer5[8][47:40] <= 'd0;
        layer5[8][55:48] <= 'd0;
        layer6[8][7:0] <= 'd0;
        layer6[8][15:8] <= 'd0;
        layer6[8][23:16] <= 'd0;
        layer6[8][31:24] <= 'd0;
        layer6[8][39:32] <= 'd0;
        layer6[8][47:40] <= 'd0;
        layer6[8][55:48] <= 'd0;
        layer0[9][7:0] <= 'd0;
        layer0[9][15:8] <= 'd0;
        layer0[9][23:16] <= 'd0;
        layer0[9][31:24] <= 'd0;
        layer0[9][39:32] <= 'd0;
        layer0[9][47:40] <= 'd0;
        layer0[9][55:48] <= 'd0;
        layer1[9][7:0] <= 'd0;
        layer1[9][15:8] <= 'd0;
        layer1[9][23:16] <= 'd0;
        layer1[9][31:24] <= 'd0;
        layer1[9][39:32] <= 'd0;
        layer1[9][47:40] <= 'd0;
        layer1[9][55:48] <= 'd0;
        layer2[9][7:0] <= 'd0;
        layer2[9][15:8] <= 'd0;
        layer2[9][23:16] <= 'd0;
        layer2[9][31:24] <= 'd0;
        layer2[9][39:32] <= 'd0;
        layer2[9][47:40] <= 'd0;
        layer2[9][55:48] <= 'd0;
        layer3[9][7:0] <= 'd0;
        layer3[9][15:8] <= 'd0;
        layer3[9][23:16] <= 'd0;
        layer3[9][31:24] <= 'd0;
        layer3[9][39:32] <= 'd0;
        layer3[9][47:40] <= 'd0;
        layer3[9][55:48] <= 'd0;
        layer4[9][7:0] <= 'd0;
        layer4[9][15:8] <= 'd0;
        layer4[9][23:16] <= 'd0;
        layer4[9][31:24] <= 'd0;
        layer4[9][39:32] <= 'd0;
        layer4[9][47:40] <= 'd0;
        layer4[9][55:48] <= 'd0;
        layer5[9][7:0] <= 'd0;
        layer5[9][15:8] <= 'd0;
        layer5[9][23:16] <= 'd0;
        layer5[9][31:24] <= 'd0;
        layer5[9][39:32] <= 'd0;
        layer5[9][47:40] <= 'd0;
        layer5[9][55:48] <= 'd0;
        layer6[9][7:0] <= 'd0;
        layer6[9][15:8] <= 'd0;
        layer6[9][23:16] <= 'd0;
        layer6[9][31:24] <= 'd0;
        layer6[9][39:32] <= 'd0;
        layer6[9][47:40] <= 'd0;
        layer6[9][55:48] <= 'd0;
        layer0[10][7:0] <= 'd0;
        layer0[10][15:8] <= 'd0;
        layer0[10][23:16] <= 'd0;
        layer0[10][31:24] <= 'd0;
        layer0[10][39:32] <= 'd0;
        layer0[10][47:40] <= 'd0;
        layer0[10][55:48] <= 'd0;
        layer1[10][7:0] <= 'd0;
        layer1[10][15:8] <= 'd0;
        layer1[10][23:16] <= 'd0;
        layer1[10][31:24] <= 'd0;
        layer1[10][39:32] <= 'd0;
        layer1[10][47:40] <= 'd0;
        layer1[10][55:48] <= 'd0;
        layer2[10][7:0] <= 'd0;
        layer2[10][15:8] <= 'd0;
        layer2[10][23:16] <= 'd0;
        layer2[10][31:24] <= 'd0;
        layer2[10][39:32] <= 'd0;
        layer2[10][47:40] <= 'd0;
        layer2[10][55:48] <= 'd0;
        layer3[10][7:0] <= 'd0;
        layer3[10][15:8] <= 'd0;
        layer3[10][23:16] <= 'd0;
        layer3[10][31:24] <= 'd0;
        layer3[10][39:32] <= 'd0;
        layer3[10][47:40] <= 'd0;
        layer3[10][55:48] <= 'd0;
        layer4[10][7:0] <= 'd0;
        layer4[10][15:8] <= 'd0;
        layer4[10][23:16] <= 'd0;
        layer4[10][31:24] <= 'd0;
        layer4[10][39:32] <= 'd0;
        layer4[10][47:40] <= 'd0;
        layer4[10][55:48] <= 'd0;
        layer5[10][7:0] <= 'd0;
        layer5[10][15:8] <= 'd0;
        layer5[10][23:16] <= 'd0;
        layer5[10][31:24] <= 'd0;
        layer5[10][39:32] <= 'd0;
        layer5[10][47:40] <= 'd0;
        layer5[10][55:48] <= 'd0;
        layer6[10][7:0] <= 'd0;
        layer6[10][15:8] <= 'd0;
        layer6[10][23:16] <= 'd0;
        layer6[10][31:24] <= 'd0;
        layer6[10][39:32] <= 'd0;
        layer6[10][47:40] <= 'd0;
        layer6[10][55:48] <= 'd0;
        layer0[11][7:0] <= 'd0;
        layer0[11][15:8] <= 'd0;
        layer0[11][23:16] <= 'd0;
        layer0[11][31:24] <= 'd0;
        layer0[11][39:32] <= 'd0;
        layer0[11][47:40] <= 'd0;
        layer0[11][55:48] <= 'd0;
        layer1[11][7:0] <= 'd0;
        layer1[11][15:8] <= 'd0;
        layer1[11][23:16] <= 'd0;
        layer1[11][31:24] <= 'd0;
        layer1[11][39:32] <= 'd0;
        layer1[11][47:40] <= 'd0;
        layer1[11][55:48] <= 'd0;
        layer2[11][7:0] <= 'd0;
        layer2[11][15:8] <= 'd0;
        layer2[11][23:16] <= 'd0;
        layer2[11][31:24] <= 'd0;
        layer2[11][39:32] <= 'd0;
        layer2[11][47:40] <= 'd0;
        layer2[11][55:48] <= 'd0;
        layer3[11][7:0] <= 'd0;
        layer3[11][15:8] <= 'd0;
        layer3[11][23:16] <= 'd0;
        layer3[11][31:24] <= 'd0;
        layer3[11][39:32] <= 'd0;
        layer3[11][47:40] <= 'd0;
        layer3[11][55:48] <= 'd0;
        layer4[11][7:0] <= 'd0;
        layer4[11][15:8] <= 'd0;
        layer4[11][23:16] <= 'd0;
        layer4[11][31:24] <= 'd0;
        layer4[11][39:32] <= 'd0;
        layer4[11][47:40] <= 'd0;
        layer4[11][55:48] <= 'd0;
        layer5[11][7:0] <= 'd0;
        layer5[11][15:8] <= 'd0;
        layer5[11][23:16] <= 'd0;
        layer5[11][31:24] <= 'd0;
        layer5[11][39:32] <= 'd0;
        layer5[11][47:40] <= 'd0;
        layer5[11][55:48] <= 'd0;
        layer6[11][7:0] <= 'd0;
        layer6[11][15:8] <= 'd0;
        layer6[11][23:16] <= 'd0;
        layer6[11][31:24] <= 'd0;
        layer6[11][39:32] <= 'd0;
        layer6[11][47:40] <= 'd0;
        layer6[11][55:48] <= 'd0;
        layer0[12][7:0] <= 'd0;
        layer0[12][15:8] <= 'd0;
        layer0[12][23:16] <= 'd0;
        layer0[12][31:24] <= 'd0;
        layer0[12][39:32] <= 'd0;
        layer0[12][47:40] <= 'd0;
        layer0[12][55:48] <= 'd0;
        layer1[12][7:0] <= 'd0;
        layer1[12][15:8] <= 'd0;
        layer1[12][23:16] <= 'd0;
        layer1[12][31:24] <= 'd0;
        layer1[12][39:32] <= 'd0;
        layer1[12][47:40] <= 'd0;
        layer1[12][55:48] <= 'd0;
        layer2[12][7:0] <= 'd0;
        layer2[12][15:8] <= 'd0;
        layer2[12][23:16] <= 'd0;
        layer2[12][31:24] <= 'd0;
        layer2[12][39:32] <= 'd0;
        layer2[12][47:40] <= 'd0;
        layer2[12][55:48] <= 'd0;
        layer3[12][7:0] <= 'd0;
        layer3[12][15:8] <= 'd0;
        layer3[12][23:16] <= 'd0;
        layer3[12][31:24] <= 'd0;
        layer3[12][39:32] <= 'd0;
        layer3[12][47:40] <= 'd0;
        layer3[12][55:48] <= 'd0;
        layer4[12][7:0] <= 'd0;
        layer4[12][15:8] <= 'd0;
        layer4[12][23:16] <= 'd0;
        layer4[12][31:24] <= 'd0;
        layer4[12][39:32] <= 'd0;
        layer4[12][47:40] <= 'd0;
        layer4[12][55:48] <= 'd0;
        layer5[12][7:0] <= 'd0;
        layer5[12][15:8] <= 'd0;
        layer5[12][23:16] <= 'd0;
        layer5[12][31:24] <= 'd0;
        layer5[12][39:32] <= 'd0;
        layer5[12][47:40] <= 'd0;
        layer5[12][55:48] <= 'd0;
        layer6[12][7:0] <= 'd0;
        layer6[12][15:8] <= 'd0;
        layer6[12][23:16] <= 'd0;
        layer6[12][31:24] <= 'd0;
        layer6[12][39:32] <= 'd0;
        layer6[12][47:40] <= 'd0;
        layer6[12][55:48] <= 'd0;
        layer0[13][7:0] <= 'd0;
        layer0[13][15:8] <= 'd0;
        layer0[13][23:16] <= 'd0;
        layer0[13][31:24] <= 'd0;
        layer0[13][39:32] <= 'd0;
        layer0[13][47:40] <= 'd0;
        layer0[13][55:48] <= 'd0;
        layer1[13][7:0] <= 'd0;
        layer1[13][15:8] <= 'd0;
        layer1[13][23:16] <= 'd0;
        layer1[13][31:24] <= 'd0;
        layer1[13][39:32] <= 'd0;
        layer1[13][47:40] <= 'd0;
        layer1[13][55:48] <= 'd0;
        layer2[13][7:0] <= 'd0;
        layer2[13][15:8] <= 'd0;
        layer2[13][23:16] <= 'd0;
        layer2[13][31:24] <= 'd0;
        layer2[13][39:32] <= 'd0;
        layer2[13][47:40] <= 'd0;
        layer2[13][55:48] <= 'd0;
        layer3[13][7:0] <= 'd0;
        layer3[13][15:8] <= 'd0;
        layer3[13][23:16] <= 'd0;
        layer3[13][31:24] <= 'd0;
        layer3[13][39:32] <= 'd0;
        layer3[13][47:40] <= 'd0;
        layer3[13][55:48] <= 'd0;
        layer4[13][7:0] <= 'd0;
        layer4[13][15:8] <= 'd0;
        layer4[13][23:16] <= 'd0;
        layer4[13][31:24] <= 'd0;
        layer4[13][39:32] <= 'd0;
        layer4[13][47:40] <= 'd0;
        layer4[13][55:48] <= 'd0;
        layer5[13][7:0] <= 'd0;
        layer5[13][15:8] <= 'd0;
        layer5[13][23:16] <= 'd0;
        layer5[13][31:24] <= 'd0;
        layer5[13][39:32] <= 'd0;
        layer5[13][47:40] <= 'd0;
        layer5[13][55:48] <= 'd0;
        layer6[13][7:0] <= 'd0;
        layer6[13][15:8] <= 'd0;
        layer6[13][23:16] <= 'd0;
        layer6[13][31:24] <= 'd0;
        layer6[13][39:32] <= 'd0;
        layer6[13][47:40] <= 'd0;
        layer6[13][55:48] <= 'd0;
        layer0[14][7:0] <= 'd0;
        layer0[14][15:8] <= 'd0;
        layer0[14][23:16] <= 'd0;
        layer0[14][31:24] <= 'd0;
        layer0[14][39:32] <= 'd0;
        layer0[14][47:40] <= 'd0;
        layer0[14][55:48] <= 'd0;
        layer1[14][7:0] <= 'd0;
        layer1[14][15:8] <= 'd0;
        layer1[14][23:16] <= 'd0;
        layer1[14][31:24] <= 'd0;
        layer1[14][39:32] <= 'd0;
        layer1[14][47:40] <= 'd0;
        layer1[14][55:48] <= 'd0;
        layer2[14][7:0] <= 'd0;
        layer2[14][15:8] <= 'd0;
        layer2[14][23:16] <= 'd0;
        layer2[14][31:24] <= 'd0;
        layer2[14][39:32] <= 'd0;
        layer2[14][47:40] <= 'd0;
        layer2[14][55:48] <= 'd0;
        layer3[14][7:0] <= 'd0;
        layer3[14][15:8] <= 'd0;
        layer3[14][23:16] <= 'd0;
        layer3[14][31:24] <= 'd0;
        layer3[14][39:32] <= 'd0;
        layer3[14][47:40] <= 'd0;
        layer3[14][55:48] <= 'd0;
        layer4[14][7:0] <= 'd0;
        layer4[14][15:8] <= 'd0;
        layer4[14][23:16] <= 'd0;
        layer4[14][31:24] <= 'd0;
        layer4[14][39:32] <= 'd0;
        layer4[14][47:40] <= 'd0;
        layer4[14][55:48] <= 'd0;
        layer5[14][7:0] <= 'd0;
        layer5[14][15:8] <= 'd0;
        layer5[14][23:16] <= 'd0;
        layer5[14][31:24] <= 'd0;
        layer5[14][39:32] <= 'd0;
        layer5[14][47:40] <= 'd0;
        layer5[14][55:48] <= 'd0;
        layer6[14][7:0] <= 'd0;
        layer6[14][15:8] <= 'd0;
        layer6[14][23:16] <= 'd0;
        layer6[14][31:24] <= 'd0;
        layer6[14][39:32] <= 'd0;
        layer6[14][47:40] <= 'd0;
        layer6[14][55:48] <= 'd0;
        layer0[15][7:0] <= 'd0;
        layer0[15][15:8] <= 'd0;
        layer0[15][23:16] <= 'd0;
        layer0[15][31:24] <= 'd0;
        layer0[15][39:32] <= 'd0;
        layer0[15][47:40] <= 'd0;
        layer0[15][55:48] <= 'd0;
        layer1[15][7:0] <= 'd0;
        layer1[15][15:8] <= 'd0;
        layer1[15][23:16] <= 'd0;
        layer1[15][31:24] <= 'd0;
        layer1[15][39:32] <= 'd0;
        layer1[15][47:40] <= 'd0;
        layer1[15][55:48] <= 'd0;
        layer2[15][7:0] <= 'd0;
        layer2[15][15:8] <= 'd0;
        layer2[15][23:16] <= 'd0;
        layer2[15][31:24] <= 'd0;
        layer2[15][39:32] <= 'd0;
        layer2[15][47:40] <= 'd0;
        layer2[15][55:48] <= 'd0;
        layer3[15][7:0] <= 'd0;
        layer3[15][15:8] <= 'd0;
        layer3[15][23:16] <= 'd0;
        layer3[15][31:24] <= 'd0;
        layer3[15][39:32] <= 'd0;
        layer3[15][47:40] <= 'd0;
        layer3[15][55:48] <= 'd0;
        layer4[15][7:0] <= 'd0;
        layer4[15][15:8] <= 'd0;
        layer4[15][23:16] <= 'd0;
        layer4[15][31:24] <= 'd0;
        layer4[15][39:32] <= 'd0;
        layer4[15][47:40] <= 'd0;
        layer4[15][55:48] <= 'd0;
        layer5[15][7:0] <= 'd0;
        layer5[15][15:8] <= 'd0;
        layer5[15][23:16] <= 'd0;
        layer5[15][31:24] <= 'd0;
        layer5[15][39:32] <= 'd0;
        layer5[15][47:40] <= 'd0;
        layer5[15][55:48] <= 'd0;
        layer6[15][7:0] <= 'd0;
        layer6[15][15:8] <= 'd0;
        layer6[15][23:16] <= 'd0;
        layer6[15][31:24] <= 'd0;
        layer6[15][39:32] <= 'd0;
        layer6[15][47:40] <= 'd0;
        layer6[15][55:48] <= 'd0;
    end
  endcase
end

reg  [15:0]  kernel_img_mul_0[0:48];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_0[0] <= 'd0;
    kernel_img_mul_0[1] <= 'd0;
    kernel_img_mul_0[2] <= 'd0;
    kernel_img_mul_0[3] <= 'd0;
    kernel_img_mul_0[4] <= 'd0;
    kernel_img_mul_0[5] <= 'd0;
    kernel_img_mul_0[6] <= 'd0;
    kernel_img_mul_0[7] <= 'd0;
    kernel_img_mul_0[8] <= 'd0;
    kernel_img_mul_0[9] <= 'd0;
    kernel_img_mul_0[10] <= 'd0;
    kernel_img_mul_0[11] <= 'd0;
    kernel_img_mul_0[12] <= 'd0;
    kernel_img_mul_0[13] <= 'd0;
    kernel_img_mul_0[14] <= 'd0;
    kernel_img_mul_0[15] <= 'd0;
    kernel_img_mul_0[16] <= 'd0;
    kernel_img_mul_0[17] <= 'd0;
    kernel_img_mul_0[18] <= 'd0;
    kernel_img_mul_0[19] <= 'd0;
    kernel_img_mul_0[20] <= 'd0;
    kernel_img_mul_0[21] <= 'd0;
    kernel_img_mul_0[22] <= 'd0;
    kernel_img_mul_0[23] <= 'd0;
    kernel_img_mul_0[24] <= 'd0;
    kernel_img_mul_0[25] <= 'd0;
    kernel_img_mul_0[26] <= 'd0;
    kernel_img_mul_0[27] <= 'd0;
    kernel_img_mul_0[28] <= 'd0;
    kernel_img_mul_0[29] <= 'd0;
    kernel_img_mul_0[30] <= 'd0;
    kernel_img_mul_0[31] <= 'd0;
    kernel_img_mul_0[32] <= 'd0;
    kernel_img_mul_0[33] <= 'd0;
    kernel_img_mul_0[34] <= 'd0;
    kernel_img_mul_0[35] <= 'd0;
    kernel_img_mul_0[36] <= 'd0;
    kernel_img_mul_0[37] <= 'd0;
    kernel_img_mul_0[38] <= 'd0;
    kernel_img_mul_0[39] <= 'd0;
    kernel_img_mul_0[40] <= 'd0;
    kernel_img_mul_0[41] <= 'd0;
    kernel_img_mul_0[42] <= 'd0;
    kernel_img_mul_0[43] <= 'd0;
    kernel_img_mul_0[44] <= 'd0;
    kernel_img_mul_0[45] <= 'd0;
    kernel_img_mul_0[46] <= 'd0;
    kernel_img_mul_0[47] <= 'd0;
    kernel_img_mul_0[48] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_0[0] <= { {8{1'b0}},layer0[0][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_0[1] <= { {8{1'b0}},layer0[0][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_0[2] <= { {8{1'b0}},layer0[0][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_0[3] <= { {8{1'b0}},layer0[0][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_0[4] <= { {8{1'b0}},layer0[0][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_0[5] <= { {8{1'b0}},layer0[0][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_0[6] <= { {8{1'b0}},layer0[0][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
    kernel_img_mul_0[7] <= { {8{1'b0}},layer1[0][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_0[8] <= { {8{1'b0}},layer1[0][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_0[9] <= { {8{1'b0}},layer1[0][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_0[10] <= { {8{1'b0}},layer1[0][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_0[11] <= { {8{1'b0}},layer1[0][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_0[12] <= { {8{1'b0}},layer1[0][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_0[13] <= { {8{1'b0}},layer1[0][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_0[14] <= { {8{1'b0}},layer2[0][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_0[15] <= { {8{1'b0}},layer2[0][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_0[16] <= { {8{1'b0}},layer2[0][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_0[17] <= { {8{1'b0}},layer2[0][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_0[18] <= { {8{1'b0}},layer2[0][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_0[19] <= { {8{1'b0}},layer2[0][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_0[20] <= { {8{1'b0}},layer2[0][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_0[21] <= { {8{1'b0}},layer3[0][7:0]} * { {8{1'b0}}, G_Kernel_7x7_3[7:0]};
    kernel_img_mul_0[22] <= { {8{1'b0}},layer3[0][15:8]} * { {8{1'b0}}, G_Kernel_7x7_3[15:8]};
    kernel_img_mul_0[23] <= { {8{1'b0}},layer3[0][23:16]} * { {8{1'b0}}, G_Kernel_7x7_3[23:16]};
    kernel_img_mul_0[24] <= { {8{1'b0}},layer3[0][31:24]} * { {8{1'b0}}, G_Kernel_7x7_3[31:24]};
    kernel_img_mul_0[25] <= { {8{1'b0}},layer3[0][39:32]} * { {8{1'b0}}, G_Kernel_7x7_3[39:32]};
    kernel_img_mul_0[26] <= { {8{1'b0}},layer3[0][47:40]} * { {8{1'b0}}, G_Kernel_7x7_3[47:40]};
    kernel_img_mul_0[27] <= { {8{1'b0}},layer3[0][55:48]} * { {8{1'b0}}, G_Kernel_7x7_3[55:48]};
    kernel_img_mul_0[28] <= { {8{1'b0}},layer4[0][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_0[29] <= { {8{1'b0}},layer4[0][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_0[30] <= { {8{1'b0}},layer4[0][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_0[31] <= { {8{1'b0}},layer4[0][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_0[32] <= { {8{1'b0}},layer4[0][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_0[33] <= { {8{1'b0}},layer4[0][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_0[34] <= { {8{1'b0}},layer4[0][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_0[35] <= { {8{1'b0}},layer5[0][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_0[36] <= { {8{1'b0}},layer5[0][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_0[37] <= { {8{1'b0}},layer5[0][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_0[38] <= { {8{1'b0}},layer5[0][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_0[39] <= { {8{1'b0}},layer5[0][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_0[40] <= { {8{1'b0}},layer5[0][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_0[41] <= { {8{1'b0}},layer5[0][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_0[42] <= { {8{1'b0}},layer6[0][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_0[43] <= { {8{1'b0}},layer6[0][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_0[44] <= { {8{1'b0}},layer6[0][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_0[45] <= { {8{1'b0}},layer6[0][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_0[46] <= { {8{1'b0}},layer6[0][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_0[47] <= { {8{1'b0}},layer6[0][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_0[48] <= { {8{1'b0}},layer6[0][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
  end
end
reg  [15:0]  kernel_img_sum_1_0;
reg  [15:0]  kernel_img_sum_2_0;
reg  [15:0]  kernel_img_sum_3_0;
reg  [15:0]  kernel_img_sum_4_0;
reg  [15:0]  kernel_img_sum_5_0;
reg  [15:0]  kernel_img_sum_6_0;
reg  [15:0]  kernel_img_sum_7_0;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_0 <= kernel_img_mul_0[0] + kernel_img_mul_0[1] + kernel_img_mul_0[2] + kernel_img_mul_0[3] + kernel_img_mul_0[4] + kernel_img_mul_0[5] + kernel_img_mul_0[6] + kernel_img_mul_0[7] + kernel_img_mul_0[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_0 <= kernel_img_mul_0[9] + kernel_img_mul_0[10] + kernel_img_mul_0[11] + kernel_img_mul_0[12] + kernel_img_mul_0[13] + kernel_img_mul_0[14] + kernel_img_mul_0[15] + kernel_img_mul_0[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_0 <= kernel_img_mul_0[17] + kernel_img_mul_0[18] + kernel_img_mul_0[19] + kernel_img_mul_0[20] + kernel_img_mul_0[21] + kernel_img_mul_0[22] + kernel_img_mul_0[23] + kernel_img_mul_0[24];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_0 <= kernel_img_mul_0[25] + kernel_img_mul_0[26] + kernel_img_mul_0[27] + kernel_img_mul_0[28] + kernel_img_mul_0[29] + kernel_img_mul_0[30] + kernel_img_mul_0[31] + kernel_img_mul_0[32];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_0 <= kernel_img_mul_0[33] + kernel_img_mul_0[34] + kernel_img_mul_0[35] + kernel_img_mul_0[36] + kernel_img_mul_0[37] + kernel_img_mul_0[38] + kernel_img_mul_0[39] + kernel_img_mul_0[40];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_0 <= kernel_img_mul_0[41] + kernel_img_mul_0[42] + kernel_img_mul_0[43] + kernel_img_mul_0[44] + kernel_img_mul_0[45] + kernel_img_mul_0[46] + kernel_img_mul_0[47] + kernel_img_mul_0[48];
  end
end
always@(*) begin
  kernel_img_sum_7_0 = kernel_img_sum_1_0 + kernel_img_sum_2_0 + kernel_img_sum_3_0 + kernel_img_sum_4_0 + kernel_img_sum_5_0 + kernel_img_sum_6_0;
end
reg  [15:0]  kernel_img_mul_1[0:48];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_1[0] <= 'd0;
    kernel_img_mul_1[1] <= 'd0;
    kernel_img_mul_1[2] <= 'd0;
    kernel_img_mul_1[3] <= 'd0;
    kernel_img_mul_1[4] <= 'd0;
    kernel_img_mul_1[5] <= 'd0;
    kernel_img_mul_1[6] <= 'd0;
    kernel_img_mul_1[7] <= 'd0;
    kernel_img_mul_1[8] <= 'd0;
    kernel_img_mul_1[9] <= 'd0;
    kernel_img_mul_1[10] <= 'd0;
    kernel_img_mul_1[11] <= 'd0;
    kernel_img_mul_1[12] <= 'd0;
    kernel_img_mul_1[13] <= 'd0;
    kernel_img_mul_1[14] <= 'd0;
    kernel_img_mul_1[15] <= 'd0;
    kernel_img_mul_1[16] <= 'd0;
    kernel_img_mul_1[17] <= 'd0;
    kernel_img_mul_1[18] <= 'd0;
    kernel_img_mul_1[19] <= 'd0;
    kernel_img_mul_1[20] <= 'd0;
    kernel_img_mul_1[21] <= 'd0;
    kernel_img_mul_1[22] <= 'd0;
    kernel_img_mul_1[23] <= 'd0;
    kernel_img_mul_1[24] <= 'd0;
    kernel_img_mul_1[25] <= 'd0;
    kernel_img_mul_1[26] <= 'd0;
    kernel_img_mul_1[27] <= 'd0;
    kernel_img_mul_1[28] <= 'd0;
    kernel_img_mul_1[29] <= 'd0;
    kernel_img_mul_1[30] <= 'd0;
    kernel_img_mul_1[31] <= 'd0;
    kernel_img_mul_1[32] <= 'd0;
    kernel_img_mul_1[33] <= 'd0;
    kernel_img_mul_1[34] <= 'd0;
    kernel_img_mul_1[35] <= 'd0;
    kernel_img_mul_1[36] <= 'd0;
    kernel_img_mul_1[37] <= 'd0;
    kernel_img_mul_1[38] <= 'd0;
    kernel_img_mul_1[39] <= 'd0;
    kernel_img_mul_1[40] <= 'd0;
    kernel_img_mul_1[41] <= 'd0;
    kernel_img_mul_1[42] <= 'd0;
    kernel_img_mul_1[43] <= 'd0;
    kernel_img_mul_1[44] <= 'd0;
    kernel_img_mul_1[45] <= 'd0;
    kernel_img_mul_1[46] <= 'd0;
    kernel_img_mul_1[47] <= 'd0;
    kernel_img_mul_1[48] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_1[0] <= { {8{1'b0}},layer0[1][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_1[1] <= { {8{1'b0}},layer0[1][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_1[2] <= { {8{1'b0}},layer0[1][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_1[3] <= { {8{1'b0}},layer0[1][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_1[4] <= { {8{1'b0}},layer0[1][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_1[5] <= { {8{1'b0}},layer0[1][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_1[6] <= { {8{1'b0}},layer0[1][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
    kernel_img_mul_1[7] <= { {8{1'b0}},layer1[1][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_1[8] <= { {8{1'b0}},layer1[1][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_1[9] <= { {8{1'b0}},layer1[1][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_1[10] <= { {8{1'b0}},layer1[1][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_1[11] <= { {8{1'b0}},layer1[1][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_1[12] <= { {8{1'b0}},layer1[1][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_1[13] <= { {8{1'b0}},layer1[1][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_1[14] <= { {8{1'b0}},layer2[1][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_1[15] <= { {8{1'b0}},layer2[1][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_1[16] <= { {8{1'b0}},layer2[1][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_1[17] <= { {8{1'b0}},layer2[1][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_1[18] <= { {8{1'b0}},layer2[1][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_1[19] <= { {8{1'b0}},layer2[1][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_1[20] <= { {8{1'b0}},layer2[1][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_1[21] <= { {8{1'b0}},layer3[1][7:0]} * { {8{1'b0}}, G_Kernel_7x7_3[7:0]};
    kernel_img_mul_1[22] <= { {8{1'b0}},layer3[1][15:8]} * { {8{1'b0}}, G_Kernel_7x7_3[15:8]};
    kernel_img_mul_1[23] <= { {8{1'b0}},layer3[1][23:16]} * { {8{1'b0}}, G_Kernel_7x7_3[23:16]};
    kernel_img_mul_1[24] <= { {8{1'b0}},layer3[1][31:24]} * { {8{1'b0}}, G_Kernel_7x7_3[31:24]};
    kernel_img_mul_1[25] <= { {8{1'b0}},layer3[1][39:32]} * { {8{1'b0}}, G_Kernel_7x7_3[39:32]};
    kernel_img_mul_1[26] <= { {8{1'b0}},layer3[1][47:40]} * { {8{1'b0}}, G_Kernel_7x7_3[47:40]};
    kernel_img_mul_1[27] <= { {8{1'b0}},layer3[1][55:48]} * { {8{1'b0}}, G_Kernel_7x7_3[55:48]};
    kernel_img_mul_1[28] <= { {8{1'b0}},layer4[1][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_1[29] <= { {8{1'b0}},layer4[1][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_1[30] <= { {8{1'b0}},layer4[1][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_1[31] <= { {8{1'b0}},layer4[1][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_1[32] <= { {8{1'b0}},layer4[1][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_1[33] <= { {8{1'b0}},layer4[1][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_1[34] <= { {8{1'b0}},layer4[1][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_1[35] <= { {8{1'b0}},layer5[1][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_1[36] <= { {8{1'b0}},layer5[1][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_1[37] <= { {8{1'b0}},layer5[1][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_1[38] <= { {8{1'b0}},layer5[1][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_1[39] <= { {8{1'b0}},layer5[1][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_1[40] <= { {8{1'b0}},layer5[1][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_1[41] <= { {8{1'b0}},layer5[1][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_1[42] <= { {8{1'b0}},layer6[1][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_1[43] <= { {8{1'b0}},layer6[1][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_1[44] <= { {8{1'b0}},layer6[1][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_1[45] <= { {8{1'b0}},layer6[1][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_1[46] <= { {8{1'b0}},layer6[1][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_1[47] <= { {8{1'b0}},layer6[1][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_1[48] <= { {8{1'b0}},layer6[1][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
  end
end
reg  [15:0]  kernel_img_sum_1_1;
reg  [15:0]  kernel_img_sum_2_1;
reg  [15:0]  kernel_img_sum_3_1;
reg  [15:0]  kernel_img_sum_4_1;
reg  [15:0]  kernel_img_sum_5_1;
reg  [15:0]  kernel_img_sum_6_1;
reg  [15:0]  kernel_img_sum_7_1;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_1 <= kernel_img_mul_1[0] + kernel_img_mul_1[1] + kernel_img_mul_1[2] + kernel_img_mul_1[3] + kernel_img_mul_1[4] + kernel_img_mul_1[5] + kernel_img_mul_1[6] + kernel_img_mul_1[7] + kernel_img_mul_1[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_1 <= kernel_img_mul_1[9] + kernel_img_mul_1[10] + kernel_img_mul_1[11] + kernel_img_mul_1[12] + kernel_img_mul_1[13] + kernel_img_mul_1[14] + kernel_img_mul_1[15] + kernel_img_mul_1[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_1 <= kernel_img_mul_1[17] + kernel_img_mul_1[18] + kernel_img_mul_1[19] + kernel_img_mul_1[20] + kernel_img_mul_1[21] + kernel_img_mul_1[22] + kernel_img_mul_1[23] + kernel_img_mul_1[24];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_1 <= kernel_img_mul_1[25] + kernel_img_mul_1[26] + kernel_img_mul_1[27] + kernel_img_mul_1[28] + kernel_img_mul_1[29] + kernel_img_mul_1[30] + kernel_img_mul_1[31] + kernel_img_mul_1[32];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_1 <= kernel_img_mul_1[33] + kernel_img_mul_1[34] + kernel_img_mul_1[35] + kernel_img_mul_1[36] + kernel_img_mul_1[37] + kernel_img_mul_1[38] + kernel_img_mul_1[39] + kernel_img_mul_1[40];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_1 <= kernel_img_mul_1[41] + kernel_img_mul_1[42] + kernel_img_mul_1[43] + kernel_img_mul_1[44] + kernel_img_mul_1[45] + kernel_img_mul_1[46] + kernel_img_mul_1[47] + kernel_img_mul_1[48];
  end
end
always@(*) begin
  kernel_img_sum_7_1 = kernel_img_sum_1_1 + kernel_img_sum_2_1 + kernel_img_sum_3_1 + kernel_img_sum_4_1 + kernel_img_sum_5_1 + kernel_img_sum_6_1;
end
reg  [15:0]  kernel_img_mul_2[0:48];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_2[0] <= 'd0;
    kernel_img_mul_2[1] <= 'd0;
    kernel_img_mul_2[2] <= 'd0;
    kernel_img_mul_2[3] <= 'd0;
    kernel_img_mul_2[4] <= 'd0;
    kernel_img_mul_2[5] <= 'd0;
    kernel_img_mul_2[6] <= 'd0;
    kernel_img_mul_2[7] <= 'd0;
    kernel_img_mul_2[8] <= 'd0;
    kernel_img_mul_2[9] <= 'd0;
    kernel_img_mul_2[10] <= 'd0;
    kernel_img_mul_2[11] <= 'd0;
    kernel_img_mul_2[12] <= 'd0;
    kernel_img_mul_2[13] <= 'd0;
    kernel_img_mul_2[14] <= 'd0;
    kernel_img_mul_2[15] <= 'd0;
    kernel_img_mul_2[16] <= 'd0;
    kernel_img_mul_2[17] <= 'd0;
    kernel_img_mul_2[18] <= 'd0;
    kernel_img_mul_2[19] <= 'd0;
    kernel_img_mul_2[20] <= 'd0;
    kernel_img_mul_2[21] <= 'd0;
    kernel_img_mul_2[22] <= 'd0;
    kernel_img_mul_2[23] <= 'd0;
    kernel_img_mul_2[24] <= 'd0;
    kernel_img_mul_2[25] <= 'd0;
    kernel_img_mul_2[26] <= 'd0;
    kernel_img_mul_2[27] <= 'd0;
    kernel_img_mul_2[28] <= 'd0;
    kernel_img_mul_2[29] <= 'd0;
    kernel_img_mul_2[30] <= 'd0;
    kernel_img_mul_2[31] <= 'd0;
    kernel_img_mul_2[32] <= 'd0;
    kernel_img_mul_2[33] <= 'd0;
    kernel_img_mul_2[34] <= 'd0;
    kernel_img_mul_2[35] <= 'd0;
    kernel_img_mul_2[36] <= 'd0;
    kernel_img_mul_2[37] <= 'd0;
    kernel_img_mul_2[38] <= 'd0;
    kernel_img_mul_2[39] <= 'd0;
    kernel_img_mul_2[40] <= 'd0;
    kernel_img_mul_2[41] <= 'd0;
    kernel_img_mul_2[42] <= 'd0;
    kernel_img_mul_2[43] <= 'd0;
    kernel_img_mul_2[44] <= 'd0;
    kernel_img_mul_2[45] <= 'd0;
    kernel_img_mul_2[46] <= 'd0;
    kernel_img_mul_2[47] <= 'd0;
    kernel_img_mul_2[48] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_2[0] <= { {8{1'b0}},layer0[2][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_2[1] <= { {8{1'b0}},layer0[2][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_2[2] <= { {8{1'b0}},layer0[2][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_2[3] <= { {8{1'b0}},layer0[2][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_2[4] <= { {8{1'b0}},layer0[2][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_2[5] <= { {8{1'b0}},layer0[2][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_2[6] <= { {8{1'b0}},layer0[2][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
    kernel_img_mul_2[7] <= { {8{1'b0}},layer1[2][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_2[8] <= { {8{1'b0}},layer1[2][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_2[9] <= { {8{1'b0}},layer1[2][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_2[10] <= { {8{1'b0}},layer1[2][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_2[11] <= { {8{1'b0}},layer1[2][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_2[12] <= { {8{1'b0}},layer1[2][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_2[13] <= { {8{1'b0}},layer1[2][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_2[14] <= { {8{1'b0}},layer2[2][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_2[15] <= { {8{1'b0}},layer2[2][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_2[16] <= { {8{1'b0}},layer2[2][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_2[17] <= { {8{1'b0}},layer2[2][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_2[18] <= { {8{1'b0}},layer2[2][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_2[19] <= { {8{1'b0}},layer2[2][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_2[20] <= { {8{1'b0}},layer2[2][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_2[21] <= { {8{1'b0}},layer3[2][7:0]} * { {8{1'b0}}, G_Kernel_7x7_3[7:0]};
    kernel_img_mul_2[22] <= { {8{1'b0}},layer3[2][15:8]} * { {8{1'b0}}, G_Kernel_7x7_3[15:8]};
    kernel_img_mul_2[23] <= { {8{1'b0}},layer3[2][23:16]} * { {8{1'b0}}, G_Kernel_7x7_3[23:16]};
    kernel_img_mul_2[24] <= { {8{1'b0}},layer3[2][31:24]} * { {8{1'b0}}, G_Kernel_7x7_3[31:24]};
    kernel_img_mul_2[25] <= { {8{1'b0}},layer3[2][39:32]} * { {8{1'b0}}, G_Kernel_7x7_3[39:32]};
    kernel_img_mul_2[26] <= { {8{1'b0}},layer3[2][47:40]} * { {8{1'b0}}, G_Kernel_7x7_3[47:40]};
    kernel_img_mul_2[27] <= { {8{1'b0}},layer3[2][55:48]} * { {8{1'b0}}, G_Kernel_7x7_3[55:48]};
    kernel_img_mul_2[28] <= { {8{1'b0}},layer4[2][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_2[29] <= { {8{1'b0}},layer4[2][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_2[30] <= { {8{1'b0}},layer4[2][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_2[31] <= { {8{1'b0}},layer4[2][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_2[32] <= { {8{1'b0}},layer4[2][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_2[33] <= { {8{1'b0}},layer4[2][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_2[34] <= { {8{1'b0}},layer4[2][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_2[35] <= { {8{1'b0}},layer5[2][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_2[36] <= { {8{1'b0}},layer5[2][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_2[37] <= { {8{1'b0}},layer5[2][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_2[38] <= { {8{1'b0}},layer5[2][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_2[39] <= { {8{1'b0}},layer5[2][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_2[40] <= { {8{1'b0}},layer5[2][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_2[41] <= { {8{1'b0}},layer5[2][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_2[42] <= { {8{1'b0}},layer6[2][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_2[43] <= { {8{1'b0}},layer6[2][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_2[44] <= { {8{1'b0}},layer6[2][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_2[45] <= { {8{1'b0}},layer6[2][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_2[46] <= { {8{1'b0}},layer6[2][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_2[47] <= { {8{1'b0}},layer6[2][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_2[48] <= { {8{1'b0}},layer6[2][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
  end
end
reg  [15:0]  kernel_img_sum_1_2;
reg  [15:0]  kernel_img_sum_2_2;
reg  [15:0]  kernel_img_sum_3_2;
reg  [15:0]  kernel_img_sum_4_2;
reg  [15:0]  kernel_img_sum_5_2;
reg  [15:0]  kernel_img_sum_6_2;
reg  [15:0]  kernel_img_sum_7_2;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_2 <= kernel_img_mul_2[0] + kernel_img_mul_2[1] + kernel_img_mul_2[2] + kernel_img_mul_2[3] + kernel_img_mul_2[4] + kernel_img_mul_2[5] + kernel_img_mul_2[6] + kernel_img_mul_2[7] + kernel_img_mul_2[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_2 <= kernel_img_mul_2[9] + kernel_img_mul_2[10] + kernel_img_mul_2[11] + kernel_img_mul_2[12] + kernel_img_mul_2[13] + kernel_img_mul_2[14] + kernel_img_mul_2[15] + kernel_img_mul_2[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_2 <= kernel_img_mul_2[17] + kernel_img_mul_2[18] + kernel_img_mul_2[19] + kernel_img_mul_2[20] + kernel_img_mul_2[21] + kernel_img_mul_2[22] + kernel_img_mul_2[23] + kernel_img_mul_2[24];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_2 <= kernel_img_mul_2[25] + kernel_img_mul_2[26] + kernel_img_mul_2[27] + kernel_img_mul_2[28] + kernel_img_mul_2[29] + kernel_img_mul_2[30] + kernel_img_mul_2[31] + kernel_img_mul_2[32];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_2 <= kernel_img_mul_2[33] + kernel_img_mul_2[34] + kernel_img_mul_2[35] + kernel_img_mul_2[36] + kernel_img_mul_2[37] + kernel_img_mul_2[38] + kernel_img_mul_2[39] + kernel_img_mul_2[40];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_2 <= kernel_img_mul_2[41] + kernel_img_mul_2[42] + kernel_img_mul_2[43] + kernel_img_mul_2[44] + kernel_img_mul_2[45] + kernel_img_mul_2[46] + kernel_img_mul_2[47] + kernel_img_mul_2[48];
  end
end
always@(*) begin
  kernel_img_sum_7_2 = kernel_img_sum_1_2 + kernel_img_sum_2_2 + kernel_img_sum_3_2 + kernel_img_sum_4_2 + kernel_img_sum_5_2 + kernel_img_sum_6_2;
end
reg  [15:0]  kernel_img_mul_3[0:48];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_3[0] <= 'd0;
    kernel_img_mul_3[1] <= 'd0;
    kernel_img_mul_3[2] <= 'd0;
    kernel_img_mul_3[3] <= 'd0;
    kernel_img_mul_3[4] <= 'd0;
    kernel_img_mul_3[5] <= 'd0;
    kernel_img_mul_3[6] <= 'd0;
    kernel_img_mul_3[7] <= 'd0;
    kernel_img_mul_3[8] <= 'd0;
    kernel_img_mul_3[9] <= 'd0;
    kernel_img_mul_3[10] <= 'd0;
    kernel_img_mul_3[11] <= 'd0;
    kernel_img_mul_3[12] <= 'd0;
    kernel_img_mul_3[13] <= 'd0;
    kernel_img_mul_3[14] <= 'd0;
    kernel_img_mul_3[15] <= 'd0;
    kernel_img_mul_3[16] <= 'd0;
    kernel_img_mul_3[17] <= 'd0;
    kernel_img_mul_3[18] <= 'd0;
    kernel_img_mul_3[19] <= 'd0;
    kernel_img_mul_3[20] <= 'd0;
    kernel_img_mul_3[21] <= 'd0;
    kernel_img_mul_3[22] <= 'd0;
    kernel_img_mul_3[23] <= 'd0;
    kernel_img_mul_3[24] <= 'd0;
    kernel_img_mul_3[25] <= 'd0;
    kernel_img_mul_3[26] <= 'd0;
    kernel_img_mul_3[27] <= 'd0;
    kernel_img_mul_3[28] <= 'd0;
    kernel_img_mul_3[29] <= 'd0;
    kernel_img_mul_3[30] <= 'd0;
    kernel_img_mul_3[31] <= 'd0;
    kernel_img_mul_3[32] <= 'd0;
    kernel_img_mul_3[33] <= 'd0;
    kernel_img_mul_3[34] <= 'd0;
    kernel_img_mul_3[35] <= 'd0;
    kernel_img_mul_3[36] <= 'd0;
    kernel_img_mul_3[37] <= 'd0;
    kernel_img_mul_3[38] <= 'd0;
    kernel_img_mul_3[39] <= 'd0;
    kernel_img_mul_3[40] <= 'd0;
    kernel_img_mul_3[41] <= 'd0;
    kernel_img_mul_3[42] <= 'd0;
    kernel_img_mul_3[43] <= 'd0;
    kernel_img_mul_3[44] <= 'd0;
    kernel_img_mul_3[45] <= 'd0;
    kernel_img_mul_3[46] <= 'd0;
    kernel_img_mul_3[47] <= 'd0;
    kernel_img_mul_3[48] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_3[0] <= { {8{1'b0}},layer0[3][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_3[1] <= { {8{1'b0}},layer0[3][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_3[2] <= { {8{1'b0}},layer0[3][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_3[3] <= { {8{1'b0}},layer0[3][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_3[4] <= { {8{1'b0}},layer0[3][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_3[5] <= { {8{1'b0}},layer0[3][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_3[6] <= { {8{1'b0}},layer0[3][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
    kernel_img_mul_3[7] <= { {8{1'b0}},layer1[3][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_3[8] <= { {8{1'b0}},layer1[3][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_3[9] <= { {8{1'b0}},layer1[3][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_3[10] <= { {8{1'b0}},layer1[3][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_3[11] <= { {8{1'b0}},layer1[3][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_3[12] <= { {8{1'b0}},layer1[3][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_3[13] <= { {8{1'b0}},layer1[3][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_3[14] <= { {8{1'b0}},layer2[3][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_3[15] <= { {8{1'b0}},layer2[3][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_3[16] <= { {8{1'b0}},layer2[3][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_3[17] <= { {8{1'b0}},layer2[3][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_3[18] <= { {8{1'b0}},layer2[3][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_3[19] <= { {8{1'b0}},layer2[3][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_3[20] <= { {8{1'b0}},layer2[3][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_3[21] <= { {8{1'b0}},layer3[3][7:0]} * { {8{1'b0}}, G_Kernel_7x7_3[7:0]};
    kernel_img_mul_3[22] <= { {8{1'b0}},layer3[3][15:8]} * { {8{1'b0}}, G_Kernel_7x7_3[15:8]};
    kernel_img_mul_3[23] <= { {8{1'b0}},layer3[3][23:16]} * { {8{1'b0}}, G_Kernel_7x7_3[23:16]};
    kernel_img_mul_3[24] <= { {8{1'b0}},layer3[3][31:24]} * { {8{1'b0}}, G_Kernel_7x7_3[31:24]};
    kernel_img_mul_3[25] <= { {8{1'b0}},layer3[3][39:32]} * { {8{1'b0}}, G_Kernel_7x7_3[39:32]};
    kernel_img_mul_3[26] <= { {8{1'b0}},layer3[3][47:40]} * { {8{1'b0}}, G_Kernel_7x7_3[47:40]};
    kernel_img_mul_3[27] <= { {8{1'b0}},layer3[3][55:48]} * { {8{1'b0}}, G_Kernel_7x7_3[55:48]};
    kernel_img_mul_3[28] <= { {8{1'b0}},layer4[3][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_3[29] <= { {8{1'b0}},layer4[3][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_3[30] <= { {8{1'b0}},layer4[3][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_3[31] <= { {8{1'b0}},layer4[3][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_3[32] <= { {8{1'b0}},layer4[3][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_3[33] <= { {8{1'b0}},layer4[3][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_3[34] <= { {8{1'b0}},layer4[3][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_3[35] <= { {8{1'b0}},layer5[3][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_3[36] <= { {8{1'b0}},layer5[3][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_3[37] <= { {8{1'b0}},layer5[3][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_3[38] <= { {8{1'b0}},layer5[3][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_3[39] <= { {8{1'b0}},layer5[3][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_3[40] <= { {8{1'b0}},layer5[3][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_3[41] <= { {8{1'b0}},layer5[3][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_3[42] <= { {8{1'b0}},layer6[3][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_3[43] <= { {8{1'b0}},layer6[3][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_3[44] <= { {8{1'b0}},layer6[3][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_3[45] <= { {8{1'b0}},layer6[3][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_3[46] <= { {8{1'b0}},layer6[3][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_3[47] <= { {8{1'b0}},layer6[3][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_3[48] <= { {8{1'b0}},layer6[3][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
  end
end
reg  [15:0]  kernel_img_sum_1_3;
reg  [15:0]  kernel_img_sum_2_3;
reg  [15:0]  kernel_img_sum_3_3;
reg  [15:0]  kernel_img_sum_4_3;
reg  [15:0]  kernel_img_sum_5_3;
reg  [15:0]  kernel_img_sum_6_3;
reg  [15:0]  kernel_img_sum_7_3;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_3 <= kernel_img_mul_3[0] + kernel_img_mul_3[1] + kernel_img_mul_3[2] + kernel_img_mul_3[3] + kernel_img_mul_3[4] + kernel_img_mul_3[5] + kernel_img_mul_3[6] + kernel_img_mul_3[7] + kernel_img_mul_3[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_3 <= kernel_img_mul_3[9] + kernel_img_mul_3[10] + kernel_img_mul_3[11] + kernel_img_mul_3[12] + kernel_img_mul_3[13] + kernel_img_mul_3[14] + kernel_img_mul_3[15] + kernel_img_mul_3[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_3 <= kernel_img_mul_3[17] + kernel_img_mul_3[18] + kernel_img_mul_3[19] + kernel_img_mul_3[20] + kernel_img_mul_3[21] + kernel_img_mul_3[22] + kernel_img_mul_3[23] + kernel_img_mul_3[24];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_3 <= kernel_img_mul_3[25] + kernel_img_mul_3[26] + kernel_img_mul_3[27] + kernel_img_mul_3[28] + kernel_img_mul_3[29] + kernel_img_mul_3[30] + kernel_img_mul_3[31] + kernel_img_mul_3[32];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_3 <= kernel_img_mul_3[33] + kernel_img_mul_3[34] + kernel_img_mul_3[35] + kernel_img_mul_3[36] + kernel_img_mul_3[37] + kernel_img_mul_3[38] + kernel_img_mul_3[39] + kernel_img_mul_3[40];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_3 <= kernel_img_mul_3[41] + kernel_img_mul_3[42] + kernel_img_mul_3[43] + kernel_img_mul_3[44] + kernel_img_mul_3[45] + kernel_img_mul_3[46] + kernel_img_mul_3[47] + kernel_img_mul_3[48];
  end
end
always@(*) begin
  kernel_img_sum_7_3 = kernel_img_sum_1_3 + kernel_img_sum_2_3 + kernel_img_sum_3_3 + kernel_img_sum_4_3 + kernel_img_sum_5_3 + kernel_img_sum_6_3;
end
reg  [15:0]  kernel_img_mul_4[0:48];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_4[0] <= 'd0;
    kernel_img_mul_4[1] <= 'd0;
    kernel_img_mul_4[2] <= 'd0;
    kernel_img_mul_4[3] <= 'd0;
    kernel_img_mul_4[4] <= 'd0;
    kernel_img_mul_4[5] <= 'd0;
    kernel_img_mul_4[6] <= 'd0;
    kernel_img_mul_4[7] <= 'd0;
    kernel_img_mul_4[8] <= 'd0;
    kernel_img_mul_4[9] <= 'd0;
    kernel_img_mul_4[10] <= 'd0;
    kernel_img_mul_4[11] <= 'd0;
    kernel_img_mul_4[12] <= 'd0;
    kernel_img_mul_4[13] <= 'd0;
    kernel_img_mul_4[14] <= 'd0;
    kernel_img_mul_4[15] <= 'd0;
    kernel_img_mul_4[16] <= 'd0;
    kernel_img_mul_4[17] <= 'd0;
    kernel_img_mul_4[18] <= 'd0;
    kernel_img_mul_4[19] <= 'd0;
    kernel_img_mul_4[20] <= 'd0;
    kernel_img_mul_4[21] <= 'd0;
    kernel_img_mul_4[22] <= 'd0;
    kernel_img_mul_4[23] <= 'd0;
    kernel_img_mul_4[24] <= 'd0;
    kernel_img_mul_4[25] <= 'd0;
    kernel_img_mul_4[26] <= 'd0;
    kernel_img_mul_4[27] <= 'd0;
    kernel_img_mul_4[28] <= 'd0;
    kernel_img_mul_4[29] <= 'd0;
    kernel_img_mul_4[30] <= 'd0;
    kernel_img_mul_4[31] <= 'd0;
    kernel_img_mul_4[32] <= 'd0;
    kernel_img_mul_4[33] <= 'd0;
    kernel_img_mul_4[34] <= 'd0;
    kernel_img_mul_4[35] <= 'd0;
    kernel_img_mul_4[36] <= 'd0;
    kernel_img_mul_4[37] <= 'd0;
    kernel_img_mul_4[38] <= 'd0;
    kernel_img_mul_4[39] <= 'd0;
    kernel_img_mul_4[40] <= 'd0;
    kernel_img_mul_4[41] <= 'd0;
    kernel_img_mul_4[42] <= 'd0;
    kernel_img_mul_4[43] <= 'd0;
    kernel_img_mul_4[44] <= 'd0;
    kernel_img_mul_4[45] <= 'd0;
    kernel_img_mul_4[46] <= 'd0;
    kernel_img_mul_4[47] <= 'd0;
    kernel_img_mul_4[48] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_4[0] <= { {8{1'b0}},layer0[4][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_4[1] <= { {8{1'b0}},layer0[4][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_4[2] <= { {8{1'b0}},layer0[4][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_4[3] <= { {8{1'b0}},layer0[4][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_4[4] <= { {8{1'b0}},layer0[4][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_4[5] <= { {8{1'b0}},layer0[4][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_4[6] <= { {8{1'b0}},layer0[4][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
    kernel_img_mul_4[7] <= { {8{1'b0}},layer1[4][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_4[8] <= { {8{1'b0}},layer1[4][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_4[9] <= { {8{1'b0}},layer1[4][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_4[10] <= { {8{1'b0}},layer1[4][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_4[11] <= { {8{1'b0}},layer1[4][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_4[12] <= { {8{1'b0}},layer1[4][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_4[13] <= { {8{1'b0}},layer1[4][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_4[14] <= { {8{1'b0}},layer2[4][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_4[15] <= { {8{1'b0}},layer2[4][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_4[16] <= { {8{1'b0}},layer2[4][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_4[17] <= { {8{1'b0}},layer2[4][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_4[18] <= { {8{1'b0}},layer2[4][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_4[19] <= { {8{1'b0}},layer2[4][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_4[20] <= { {8{1'b0}},layer2[4][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_4[21] <= { {8{1'b0}},layer3[4][7:0]} * { {8{1'b0}}, G_Kernel_7x7_3[7:0]};
    kernel_img_mul_4[22] <= { {8{1'b0}},layer3[4][15:8]} * { {8{1'b0}}, G_Kernel_7x7_3[15:8]};
    kernel_img_mul_4[23] <= { {8{1'b0}},layer3[4][23:16]} * { {8{1'b0}}, G_Kernel_7x7_3[23:16]};
    kernel_img_mul_4[24] <= { {8{1'b0}},layer3[4][31:24]} * { {8{1'b0}}, G_Kernel_7x7_3[31:24]};
    kernel_img_mul_4[25] <= { {8{1'b0}},layer3[4][39:32]} * { {8{1'b0}}, G_Kernel_7x7_3[39:32]};
    kernel_img_mul_4[26] <= { {8{1'b0}},layer3[4][47:40]} * { {8{1'b0}}, G_Kernel_7x7_3[47:40]};
    kernel_img_mul_4[27] <= { {8{1'b0}},layer3[4][55:48]} * { {8{1'b0}}, G_Kernel_7x7_3[55:48]};
    kernel_img_mul_4[28] <= { {8{1'b0}},layer4[4][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_4[29] <= { {8{1'b0}},layer4[4][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_4[30] <= { {8{1'b0}},layer4[4][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_4[31] <= { {8{1'b0}},layer4[4][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_4[32] <= { {8{1'b0}},layer4[4][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_4[33] <= { {8{1'b0}},layer4[4][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_4[34] <= { {8{1'b0}},layer4[4][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_4[35] <= { {8{1'b0}},layer5[4][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_4[36] <= { {8{1'b0}},layer5[4][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_4[37] <= { {8{1'b0}},layer5[4][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_4[38] <= { {8{1'b0}},layer5[4][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_4[39] <= { {8{1'b0}},layer5[4][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_4[40] <= { {8{1'b0}},layer5[4][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_4[41] <= { {8{1'b0}},layer5[4][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_4[42] <= { {8{1'b0}},layer6[4][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_4[43] <= { {8{1'b0}},layer6[4][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_4[44] <= { {8{1'b0}},layer6[4][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_4[45] <= { {8{1'b0}},layer6[4][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_4[46] <= { {8{1'b0}},layer6[4][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_4[47] <= { {8{1'b0}},layer6[4][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_4[48] <= { {8{1'b0}},layer6[4][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
  end
end
reg  [15:0]  kernel_img_sum_1_4;
reg  [15:0]  kernel_img_sum_2_4;
reg  [15:0]  kernel_img_sum_3_4;
reg  [15:0]  kernel_img_sum_4_4;
reg  [15:0]  kernel_img_sum_5_4;
reg  [15:0]  kernel_img_sum_6_4;
reg  [15:0]  kernel_img_sum_7_4;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_4 <= kernel_img_mul_4[0] + kernel_img_mul_4[1] + kernel_img_mul_4[2] + kernel_img_mul_4[3] + kernel_img_mul_4[4] + kernel_img_mul_4[5] + kernel_img_mul_4[6] + kernel_img_mul_4[7] + kernel_img_mul_4[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_4 <= kernel_img_mul_4[9] + kernel_img_mul_4[10] + kernel_img_mul_4[11] + kernel_img_mul_4[12] + kernel_img_mul_4[13] + kernel_img_mul_4[14] + kernel_img_mul_4[15] + kernel_img_mul_4[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_4 <= kernel_img_mul_4[17] + kernel_img_mul_4[18] + kernel_img_mul_4[19] + kernel_img_mul_4[20] + kernel_img_mul_4[21] + kernel_img_mul_4[22] + kernel_img_mul_4[23] + kernel_img_mul_4[24];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_4 <= kernel_img_mul_4[25] + kernel_img_mul_4[26] + kernel_img_mul_4[27] + kernel_img_mul_4[28] + kernel_img_mul_4[29] + kernel_img_mul_4[30] + kernel_img_mul_4[31] + kernel_img_mul_4[32];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_4 <= kernel_img_mul_4[33] + kernel_img_mul_4[34] + kernel_img_mul_4[35] + kernel_img_mul_4[36] + kernel_img_mul_4[37] + kernel_img_mul_4[38] + kernel_img_mul_4[39] + kernel_img_mul_4[40];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_4 <= kernel_img_mul_4[41] + kernel_img_mul_4[42] + kernel_img_mul_4[43] + kernel_img_mul_4[44] + kernel_img_mul_4[45] + kernel_img_mul_4[46] + kernel_img_mul_4[47] + kernel_img_mul_4[48];
  end
end
always@(*) begin
  kernel_img_sum_7_4 = kernel_img_sum_1_4 + kernel_img_sum_2_4 + kernel_img_sum_3_4 + kernel_img_sum_4_4 + kernel_img_sum_5_4 + kernel_img_sum_6_4;
end
reg  [15:0]  kernel_img_mul_5[0:48];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_5[0] <= 'd0;
    kernel_img_mul_5[1] <= 'd0;
    kernel_img_mul_5[2] <= 'd0;
    kernel_img_mul_5[3] <= 'd0;
    kernel_img_mul_5[4] <= 'd0;
    kernel_img_mul_5[5] <= 'd0;
    kernel_img_mul_5[6] <= 'd0;
    kernel_img_mul_5[7] <= 'd0;
    kernel_img_mul_5[8] <= 'd0;
    kernel_img_mul_5[9] <= 'd0;
    kernel_img_mul_5[10] <= 'd0;
    kernel_img_mul_5[11] <= 'd0;
    kernel_img_mul_5[12] <= 'd0;
    kernel_img_mul_5[13] <= 'd0;
    kernel_img_mul_5[14] <= 'd0;
    kernel_img_mul_5[15] <= 'd0;
    kernel_img_mul_5[16] <= 'd0;
    kernel_img_mul_5[17] <= 'd0;
    kernel_img_mul_5[18] <= 'd0;
    kernel_img_mul_5[19] <= 'd0;
    kernel_img_mul_5[20] <= 'd0;
    kernel_img_mul_5[21] <= 'd0;
    kernel_img_mul_5[22] <= 'd0;
    kernel_img_mul_5[23] <= 'd0;
    kernel_img_mul_5[24] <= 'd0;
    kernel_img_mul_5[25] <= 'd0;
    kernel_img_mul_5[26] <= 'd0;
    kernel_img_mul_5[27] <= 'd0;
    kernel_img_mul_5[28] <= 'd0;
    kernel_img_mul_5[29] <= 'd0;
    kernel_img_mul_5[30] <= 'd0;
    kernel_img_mul_5[31] <= 'd0;
    kernel_img_mul_5[32] <= 'd0;
    kernel_img_mul_5[33] <= 'd0;
    kernel_img_mul_5[34] <= 'd0;
    kernel_img_mul_5[35] <= 'd0;
    kernel_img_mul_5[36] <= 'd0;
    kernel_img_mul_5[37] <= 'd0;
    kernel_img_mul_5[38] <= 'd0;
    kernel_img_mul_5[39] <= 'd0;
    kernel_img_mul_5[40] <= 'd0;
    kernel_img_mul_5[41] <= 'd0;
    kernel_img_mul_5[42] <= 'd0;
    kernel_img_mul_5[43] <= 'd0;
    kernel_img_mul_5[44] <= 'd0;
    kernel_img_mul_5[45] <= 'd0;
    kernel_img_mul_5[46] <= 'd0;
    kernel_img_mul_5[47] <= 'd0;
    kernel_img_mul_5[48] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_5[0] <= { {8{1'b0}},layer0[5][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_5[1] <= { {8{1'b0}},layer0[5][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_5[2] <= { {8{1'b0}},layer0[5][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_5[3] <= { {8{1'b0}},layer0[5][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_5[4] <= { {8{1'b0}},layer0[5][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_5[5] <= { {8{1'b0}},layer0[5][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_5[6] <= { {8{1'b0}},layer0[5][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
    kernel_img_mul_5[7] <= { {8{1'b0}},layer1[5][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_5[8] <= { {8{1'b0}},layer1[5][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_5[9] <= { {8{1'b0}},layer1[5][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_5[10] <= { {8{1'b0}},layer1[5][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_5[11] <= { {8{1'b0}},layer1[5][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_5[12] <= { {8{1'b0}},layer1[5][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_5[13] <= { {8{1'b0}},layer1[5][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_5[14] <= { {8{1'b0}},layer2[5][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_5[15] <= { {8{1'b0}},layer2[5][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_5[16] <= { {8{1'b0}},layer2[5][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_5[17] <= { {8{1'b0}},layer2[5][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_5[18] <= { {8{1'b0}},layer2[5][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_5[19] <= { {8{1'b0}},layer2[5][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_5[20] <= { {8{1'b0}},layer2[5][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_5[21] <= { {8{1'b0}},layer3[5][7:0]} * { {8{1'b0}}, G_Kernel_7x7_3[7:0]};
    kernel_img_mul_5[22] <= { {8{1'b0}},layer3[5][15:8]} * { {8{1'b0}}, G_Kernel_7x7_3[15:8]};
    kernel_img_mul_5[23] <= { {8{1'b0}},layer3[5][23:16]} * { {8{1'b0}}, G_Kernel_7x7_3[23:16]};
    kernel_img_mul_5[24] <= { {8{1'b0}},layer3[5][31:24]} * { {8{1'b0}}, G_Kernel_7x7_3[31:24]};
    kernel_img_mul_5[25] <= { {8{1'b0}},layer3[5][39:32]} * { {8{1'b0}}, G_Kernel_7x7_3[39:32]};
    kernel_img_mul_5[26] <= { {8{1'b0}},layer3[5][47:40]} * { {8{1'b0}}, G_Kernel_7x7_3[47:40]};
    kernel_img_mul_5[27] <= { {8{1'b0}},layer3[5][55:48]} * { {8{1'b0}}, G_Kernel_7x7_3[55:48]};
    kernel_img_mul_5[28] <= { {8{1'b0}},layer4[5][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_5[29] <= { {8{1'b0}},layer4[5][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_5[30] <= { {8{1'b0}},layer4[5][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_5[31] <= { {8{1'b0}},layer4[5][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_5[32] <= { {8{1'b0}},layer4[5][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_5[33] <= { {8{1'b0}},layer4[5][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_5[34] <= { {8{1'b0}},layer4[5][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_5[35] <= { {8{1'b0}},layer5[5][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_5[36] <= { {8{1'b0}},layer5[5][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_5[37] <= { {8{1'b0}},layer5[5][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_5[38] <= { {8{1'b0}},layer5[5][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_5[39] <= { {8{1'b0}},layer5[5][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_5[40] <= { {8{1'b0}},layer5[5][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_5[41] <= { {8{1'b0}},layer5[5][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_5[42] <= { {8{1'b0}},layer6[5][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_5[43] <= { {8{1'b0}},layer6[5][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_5[44] <= { {8{1'b0}},layer6[5][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_5[45] <= { {8{1'b0}},layer6[5][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_5[46] <= { {8{1'b0}},layer6[5][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_5[47] <= { {8{1'b0}},layer6[5][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_5[48] <= { {8{1'b0}},layer6[5][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
  end
end
reg  [15:0]  kernel_img_sum_1_5;
reg  [15:0]  kernel_img_sum_2_5;
reg  [15:0]  kernel_img_sum_3_5;
reg  [15:0]  kernel_img_sum_4_5;
reg  [15:0]  kernel_img_sum_5_5;
reg  [15:0]  kernel_img_sum_6_5;
reg  [15:0]  kernel_img_sum_7_5;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_5 <= kernel_img_mul_5[0] + kernel_img_mul_5[1] + kernel_img_mul_5[2] + kernel_img_mul_5[3] + kernel_img_mul_5[4] + kernel_img_mul_5[5] + kernel_img_mul_5[6] + kernel_img_mul_5[7] + kernel_img_mul_5[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_5 <= kernel_img_mul_5[9] + kernel_img_mul_5[10] + kernel_img_mul_5[11] + kernel_img_mul_5[12] + kernel_img_mul_5[13] + kernel_img_mul_5[14] + kernel_img_mul_5[15] + kernel_img_mul_5[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_5 <= kernel_img_mul_5[17] + kernel_img_mul_5[18] + kernel_img_mul_5[19] + kernel_img_mul_5[20] + kernel_img_mul_5[21] + kernel_img_mul_5[22] + kernel_img_mul_5[23] + kernel_img_mul_5[24];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_5 <= kernel_img_mul_5[25] + kernel_img_mul_5[26] + kernel_img_mul_5[27] + kernel_img_mul_5[28] + kernel_img_mul_5[29] + kernel_img_mul_5[30] + kernel_img_mul_5[31] + kernel_img_mul_5[32];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_5 <= kernel_img_mul_5[33] + kernel_img_mul_5[34] + kernel_img_mul_5[35] + kernel_img_mul_5[36] + kernel_img_mul_5[37] + kernel_img_mul_5[38] + kernel_img_mul_5[39] + kernel_img_mul_5[40];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_5 <= kernel_img_mul_5[41] + kernel_img_mul_5[42] + kernel_img_mul_5[43] + kernel_img_mul_5[44] + kernel_img_mul_5[45] + kernel_img_mul_5[46] + kernel_img_mul_5[47] + kernel_img_mul_5[48];
  end
end
always@(*) begin
  kernel_img_sum_7_5 = kernel_img_sum_1_5 + kernel_img_sum_2_5 + kernel_img_sum_3_5 + kernel_img_sum_4_5 + kernel_img_sum_5_5 + kernel_img_sum_6_5;
end
reg  [15:0]  kernel_img_mul_6[0:48];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_6[0] <= 'd0;
    kernel_img_mul_6[1] <= 'd0;
    kernel_img_mul_6[2] <= 'd0;
    kernel_img_mul_6[3] <= 'd0;
    kernel_img_mul_6[4] <= 'd0;
    kernel_img_mul_6[5] <= 'd0;
    kernel_img_mul_6[6] <= 'd0;
    kernel_img_mul_6[7] <= 'd0;
    kernel_img_mul_6[8] <= 'd0;
    kernel_img_mul_6[9] <= 'd0;
    kernel_img_mul_6[10] <= 'd0;
    kernel_img_mul_6[11] <= 'd0;
    kernel_img_mul_6[12] <= 'd0;
    kernel_img_mul_6[13] <= 'd0;
    kernel_img_mul_6[14] <= 'd0;
    kernel_img_mul_6[15] <= 'd0;
    kernel_img_mul_6[16] <= 'd0;
    kernel_img_mul_6[17] <= 'd0;
    kernel_img_mul_6[18] <= 'd0;
    kernel_img_mul_6[19] <= 'd0;
    kernel_img_mul_6[20] <= 'd0;
    kernel_img_mul_6[21] <= 'd0;
    kernel_img_mul_6[22] <= 'd0;
    kernel_img_mul_6[23] <= 'd0;
    kernel_img_mul_6[24] <= 'd0;
    kernel_img_mul_6[25] <= 'd0;
    kernel_img_mul_6[26] <= 'd0;
    kernel_img_mul_6[27] <= 'd0;
    kernel_img_mul_6[28] <= 'd0;
    kernel_img_mul_6[29] <= 'd0;
    kernel_img_mul_6[30] <= 'd0;
    kernel_img_mul_6[31] <= 'd0;
    kernel_img_mul_6[32] <= 'd0;
    kernel_img_mul_6[33] <= 'd0;
    kernel_img_mul_6[34] <= 'd0;
    kernel_img_mul_6[35] <= 'd0;
    kernel_img_mul_6[36] <= 'd0;
    kernel_img_mul_6[37] <= 'd0;
    kernel_img_mul_6[38] <= 'd0;
    kernel_img_mul_6[39] <= 'd0;
    kernel_img_mul_6[40] <= 'd0;
    kernel_img_mul_6[41] <= 'd0;
    kernel_img_mul_6[42] <= 'd0;
    kernel_img_mul_6[43] <= 'd0;
    kernel_img_mul_6[44] <= 'd0;
    kernel_img_mul_6[45] <= 'd0;
    kernel_img_mul_6[46] <= 'd0;
    kernel_img_mul_6[47] <= 'd0;
    kernel_img_mul_6[48] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_6[0] <= { {8{1'b0}},layer0[6][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_6[1] <= { {8{1'b0}},layer0[6][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_6[2] <= { {8{1'b0}},layer0[6][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_6[3] <= { {8{1'b0}},layer0[6][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_6[4] <= { {8{1'b0}},layer0[6][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_6[5] <= { {8{1'b0}},layer0[6][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_6[6] <= { {8{1'b0}},layer0[6][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
    kernel_img_mul_6[7] <= { {8{1'b0}},layer1[6][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_6[8] <= { {8{1'b0}},layer1[6][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_6[9] <= { {8{1'b0}},layer1[6][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_6[10] <= { {8{1'b0}},layer1[6][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_6[11] <= { {8{1'b0}},layer1[6][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_6[12] <= { {8{1'b0}},layer1[6][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_6[13] <= { {8{1'b0}},layer1[6][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_6[14] <= { {8{1'b0}},layer2[6][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_6[15] <= { {8{1'b0}},layer2[6][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_6[16] <= { {8{1'b0}},layer2[6][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_6[17] <= { {8{1'b0}},layer2[6][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_6[18] <= { {8{1'b0}},layer2[6][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_6[19] <= { {8{1'b0}},layer2[6][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_6[20] <= { {8{1'b0}},layer2[6][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_6[21] <= { {8{1'b0}},layer3[6][7:0]} * { {8{1'b0}}, G_Kernel_7x7_3[7:0]};
    kernel_img_mul_6[22] <= { {8{1'b0}},layer3[6][15:8]} * { {8{1'b0}}, G_Kernel_7x7_3[15:8]};
    kernel_img_mul_6[23] <= { {8{1'b0}},layer3[6][23:16]} * { {8{1'b0}}, G_Kernel_7x7_3[23:16]};
    kernel_img_mul_6[24] <= { {8{1'b0}},layer3[6][31:24]} * { {8{1'b0}}, G_Kernel_7x7_3[31:24]};
    kernel_img_mul_6[25] <= { {8{1'b0}},layer3[6][39:32]} * { {8{1'b0}}, G_Kernel_7x7_3[39:32]};
    kernel_img_mul_6[26] <= { {8{1'b0}},layer3[6][47:40]} * { {8{1'b0}}, G_Kernel_7x7_3[47:40]};
    kernel_img_mul_6[27] <= { {8{1'b0}},layer3[6][55:48]} * { {8{1'b0}}, G_Kernel_7x7_3[55:48]};
    kernel_img_mul_6[28] <= { {8{1'b0}},layer4[6][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_6[29] <= { {8{1'b0}},layer4[6][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_6[30] <= { {8{1'b0}},layer4[6][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_6[31] <= { {8{1'b0}},layer4[6][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_6[32] <= { {8{1'b0}},layer4[6][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_6[33] <= { {8{1'b0}},layer4[6][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_6[34] <= { {8{1'b0}},layer4[6][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_6[35] <= { {8{1'b0}},layer5[6][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_6[36] <= { {8{1'b0}},layer5[6][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_6[37] <= { {8{1'b0}},layer5[6][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_6[38] <= { {8{1'b0}},layer5[6][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_6[39] <= { {8{1'b0}},layer5[6][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_6[40] <= { {8{1'b0}},layer5[6][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_6[41] <= { {8{1'b0}},layer5[6][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_6[42] <= { {8{1'b0}},layer6[6][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_6[43] <= { {8{1'b0}},layer6[6][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_6[44] <= { {8{1'b0}},layer6[6][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_6[45] <= { {8{1'b0}},layer6[6][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_6[46] <= { {8{1'b0}},layer6[6][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_6[47] <= { {8{1'b0}},layer6[6][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_6[48] <= { {8{1'b0}},layer6[6][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
  end
end
reg  [15:0]  kernel_img_sum_1_6;
reg  [15:0]  kernel_img_sum_2_6;
reg  [15:0]  kernel_img_sum_3_6;
reg  [15:0]  kernel_img_sum_4_6;
reg  [15:0]  kernel_img_sum_5_6;
reg  [15:0]  kernel_img_sum_6_6;
reg  [15:0]  kernel_img_sum_7_6;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_6 <= kernel_img_mul_6[0] + kernel_img_mul_6[1] + kernel_img_mul_6[2] + kernel_img_mul_6[3] + kernel_img_mul_6[4] + kernel_img_mul_6[5] + kernel_img_mul_6[6] + kernel_img_mul_6[7] + kernel_img_mul_6[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_6 <= kernel_img_mul_6[9] + kernel_img_mul_6[10] + kernel_img_mul_6[11] + kernel_img_mul_6[12] + kernel_img_mul_6[13] + kernel_img_mul_6[14] + kernel_img_mul_6[15] + kernel_img_mul_6[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_6 <= kernel_img_mul_6[17] + kernel_img_mul_6[18] + kernel_img_mul_6[19] + kernel_img_mul_6[20] + kernel_img_mul_6[21] + kernel_img_mul_6[22] + kernel_img_mul_6[23] + kernel_img_mul_6[24];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_6 <= kernel_img_mul_6[25] + kernel_img_mul_6[26] + kernel_img_mul_6[27] + kernel_img_mul_6[28] + kernel_img_mul_6[29] + kernel_img_mul_6[30] + kernel_img_mul_6[31] + kernel_img_mul_6[32];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_6 <= kernel_img_mul_6[33] + kernel_img_mul_6[34] + kernel_img_mul_6[35] + kernel_img_mul_6[36] + kernel_img_mul_6[37] + kernel_img_mul_6[38] + kernel_img_mul_6[39] + kernel_img_mul_6[40];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_6 <= kernel_img_mul_6[41] + kernel_img_mul_6[42] + kernel_img_mul_6[43] + kernel_img_mul_6[44] + kernel_img_mul_6[45] + kernel_img_mul_6[46] + kernel_img_mul_6[47] + kernel_img_mul_6[48];
  end
end
always@(*) begin
  kernel_img_sum_7_6 = kernel_img_sum_1_6 + kernel_img_sum_2_6 + kernel_img_sum_3_6 + kernel_img_sum_4_6 + kernel_img_sum_5_6 + kernel_img_sum_6_6;
end
reg  [15:0]  kernel_img_mul_7[0:48];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_7[0] <= 'd0;
    kernel_img_mul_7[1] <= 'd0;
    kernel_img_mul_7[2] <= 'd0;
    kernel_img_mul_7[3] <= 'd0;
    kernel_img_mul_7[4] <= 'd0;
    kernel_img_mul_7[5] <= 'd0;
    kernel_img_mul_7[6] <= 'd0;
    kernel_img_mul_7[7] <= 'd0;
    kernel_img_mul_7[8] <= 'd0;
    kernel_img_mul_7[9] <= 'd0;
    kernel_img_mul_7[10] <= 'd0;
    kernel_img_mul_7[11] <= 'd0;
    kernel_img_mul_7[12] <= 'd0;
    kernel_img_mul_7[13] <= 'd0;
    kernel_img_mul_7[14] <= 'd0;
    kernel_img_mul_7[15] <= 'd0;
    kernel_img_mul_7[16] <= 'd0;
    kernel_img_mul_7[17] <= 'd0;
    kernel_img_mul_7[18] <= 'd0;
    kernel_img_mul_7[19] <= 'd0;
    kernel_img_mul_7[20] <= 'd0;
    kernel_img_mul_7[21] <= 'd0;
    kernel_img_mul_7[22] <= 'd0;
    kernel_img_mul_7[23] <= 'd0;
    kernel_img_mul_7[24] <= 'd0;
    kernel_img_mul_7[25] <= 'd0;
    kernel_img_mul_7[26] <= 'd0;
    kernel_img_mul_7[27] <= 'd0;
    kernel_img_mul_7[28] <= 'd0;
    kernel_img_mul_7[29] <= 'd0;
    kernel_img_mul_7[30] <= 'd0;
    kernel_img_mul_7[31] <= 'd0;
    kernel_img_mul_7[32] <= 'd0;
    kernel_img_mul_7[33] <= 'd0;
    kernel_img_mul_7[34] <= 'd0;
    kernel_img_mul_7[35] <= 'd0;
    kernel_img_mul_7[36] <= 'd0;
    kernel_img_mul_7[37] <= 'd0;
    kernel_img_mul_7[38] <= 'd0;
    kernel_img_mul_7[39] <= 'd0;
    kernel_img_mul_7[40] <= 'd0;
    kernel_img_mul_7[41] <= 'd0;
    kernel_img_mul_7[42] <= 'd0;
    kernel_img_mul_7[43] <= 'd0;
    kernel_img_mul_7[44] <= 'd0;
    kernel_img_mul_7[45] <= 'd0;
    kernel_img_mul_7[46] <= 'd0;
    kernel_img_mul_7[47] <= 'd0;
    kernel_img_mul_7[48] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_7[0] <= { {8{1'b0}},layer0[7][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_7[1] <= { {8{1'b0}},layer0[7][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_7[2] <= { {8{1'b0}},layer0[7][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_7[3] <= { {8{1'b0}},layer0[7][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_7[4] <= { {8{1'b0}},layer0[7][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_7[5] <= { {8{1'b0}},layer0[7][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_7[6] <= { {8{1'b0}},layer0[7][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
    kernel_img_mul_7[7] <= { {8{1'b0}},layer1[7][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_7[8] <= { {8{1'b0}},layer1[7][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_7[9] <= { {8{1'b0}},layer1[7][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_7[10] <= { {8{1'b0}},layer1[7][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_7[11] <= { {8{1'b0}},layer1[7][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_7[12] <= { {8{1'b0}},layer1[7][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_7[13] <= { {8{1'b0}},layer1[7][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_7[14] <= { {8{1'b0}},layer2[7][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_7[15] <= { {8{1'b0}},layer2[7][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_7[16] <= { {8{1'b0}},layer2[7][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_7[17] <= { {8{1'b0}},layer2[7][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_7[18] <= { {8{1'b0}},layer2[7][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_7[19] <= { {8{1'b0}},layer2[7][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_7[20] <= { {8{1'b0}},layer2[7][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_7[21] <= { {8{1'b0}},layer3[7][7:0]} * { {8{1'b0}}, G_Kernel_7x7_3[7:0]};
    kernel_img_mul_7[22] <= { {8{1'b0}},layer3[7][15:8]} * { {8{1'b0}}, G_Kernel_7x7_3[15:8]};
    kernel_img_mul_7[23] <= { {8{1'b0}},layer3[7][23:16]} * { {8{1'b0}}, G_Kernel_7x7_3[23:16]};
    kernel_img_mul_7[24] <= { {8{1'b0}},layer3[7][31:24]} * { {8{1'b0}}, G_Kernel_7x7_3[31:24]};
    kernel_img_mul_7[25] <= { {8{1'b0}},layer3[7][39:32]} * { {8{1'b0}}, G_Kernel_7x7_3[39:32]};
    kernel_img_mul_7[26] <= { {8{1'b0}},layer3[7][47:40]} * { {8{1'b0}}, G_Kernel_7x7_3[47:40]};
    kernel_img_mul_7[27] <= { {8{1'b0}},layer3[7][55:48]} * { {8{1'b0}}, G_Kernel_7x7_3[55:48]};
    kernel_img_mul_7[28] <= { {8{1'b0}},layer4[7][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_7[29] <= { {8{1'b0}},layer4[7][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_7[30] <= { {8{1'b0}},layer4[7][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_7[31] <= { {8{1'b0}},layer4[7][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_7[32] <= { {8{1'b0}},layer4[7][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_7[33] <= { {8{1'b0}},layer4[7][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_7[34] <= { {8{1'b0}},layer4[7][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_7[35] <= { {8{1'b0}},layer5[7][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_7[36] <= { {8{1'b0}},layer5[7][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_7[37] <= { {8{1'b0}},layer5[7][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_7[38] <= { {8{1'b0}},layer5[7][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_7[39] <= { {8{1'b0}},layer5[7][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_7[40] <= { {8{1'b0}},layer5[7][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_7[41] <= { {8{1'b0}},layer5[7][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_7[42] <= { {8{1'b0}},layer6[7][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_7[43] <= { {8{1'b0}},layer6[7][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_7[44] <= { {8{1'b0}},layer6[7][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_7[45] <= { {8{1'b0}},layer6[7][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_7[46] <= { {8{1'b0}},layer6[7][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_7[47] <= { {8{1'b0}},layer6[7][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_7[48] <= { {8{1'b0}},layer6[7][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
  end
end
reg  [15:0]  kernel_img_sum_1_7;
reg  [15:0]  kernel_img_sum_2_7;
reg  [15:0]  kernel_img_sum_3_7;
reg  [15:0]  kernel_img_sum_4_7;
reg  [15:0]  kernel_img_sum_5_7;
reg  [15:0]  kernel_img_sum_6_7;
reg  [15:0]  kernel_img_sum_7_7;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_7 <= kernel_img_mul_7[0] + kernel_img_mul_7[1] + kernel_img_mul_7[2] + kernel_img_mul_7[3] + kernel_img_mul_7[4] + kernel_img_mul_7[5] + kernel_img_mul_7[6] + kernel_img_mul_7[7] + kernel_img_mul_7[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_7 <= kernel_img_mul_7[9] + kernel_img_mul_7[10] + kernel_img_mul_7[11] + kernel_img_mul_7[12] + kernel_img_mul_7[13] + kernel_img_mul_7[14] + kernel_img_mul_7[15] + kernel_img_mul_7[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_7 <= kernel_img_mul_7[17] + kernel_img_mul_7[18] + kernel_img_mul_7[19] + kernel_img_mul_7[20] + kernel_img_mul_7[21] + kernel_img_mul_7[22] + kernel_img_mul_7[23] + kernel_img_mul_7[24];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_7 <= kernel_img_mul_7[25] + kernel_img_mul_7[26] + kernel_img_mul_7[27] + kernel_img_mul_7[28] + kernel_img_mul_7[29] + kernel_img_mul_7[30] + kernel_img_mul_7[31] + kernel_img_mul_7[32];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_7 <= kernel_img_mul_7[33] + kernel_img_mul_7[34] + kernel_img_mul_7[35] + kernel_img_mul_7[36] + kernel_img_mul_7[37] + kernel_img_mul_7[38] + kernel_img_mul_7[39] + kernel_img_mul_7[40];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_7 <= kernel_img_mul_7[41] + kernel_img_mul_7[42] + kernel_img_mul_7[43] + kernel_img_mul_7[44] + kernel_img_mul_7[45] + kernel_img_mul_7[46] + kernel_img_mul_7[47] + kernel_img_mul_7[48];
  end
end
always@(*) begin
  kernel_img_sum_7_7 = kernel_img_sum_1_7 + kernel_img_sum_2_7 + kernel_img_sum_3_7 + kernel_img_sum_4_7 + kernel_img_sum_5_7 + kernel_img_sum_6_7;
end
reg  [15:0]  kernel_img_mul_8[0:48];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_8[0] <= 'd0;
    kernel_img_mul_8[1] <= 'd0;
    kernel_img_mul_8[2] <= 'd0;
    kernel_img_mul_8[3] <= 'd0;
    kernel_img_mul_8[4] <= 'd0;
    kernel_img_mul_8[5] <= 'd0;
    kernel_img_mul_8[6] <= 'd0;
    kernel_img_mul_8[7] <= 'd0;
    kernel_img_mul_8[8] <= 'd0;
    kernel_img_mul_8[9] <= 'd0;
    kernel_img_mul_8[10] <= 'd0;
    kernel_img_mul_8[11] <= 'd0;
    kernel_img_mul_8[12] <= 'd0;
    kernel_img_mul_8[13] <= 'd0;
    kernel_img_mul_8[14] <= 'd0;
    kernel_img_mul_8[15] <= 'd0;
    kernel_img_mul_8[16] <= 'd0;
    kernel_img_mul_8[17] <= 'd0;
    kernel_img_mul_8[18] <= 'd0;
    kernel_img_mul_8[19] <= 'd0;
    kernel_img_mul_8[20] <= 'd0;
    kernel_img_mul_8[21] <= 'd0;
    kernel_img_mul_8[22] <= 'd0;
    kernel_img_mul_8[23] <= 'd0;
    kernel_img_mul_8[24] <= 'd0;
    kernel_img_mul_8[25] <= 'd0;
    kernel_img_mul_8[26] <= 'd0;
    kernel_img_mul_8[27] <= 'd0;
    kernel_img_mul_8[28] <= 'd0;
    kernel_img_mul_8[29] <= 'd0;
    kernel_img_mul_8[30] <= 'd0;
    kernel_img_mul_8[31] <= 'd0;
    kernel_img_mul_8[32] <= 'd0;
    kernel_img_mul_8[33] <= 'd0;
    kernel_img_mul_8[34] <= 'd0;
    kernel_img_mul_8[35] <= 'd0;
    kernel_img_mul_8[36] <= 'd0;
    kernel_img_mul_8[37] <= 'd0;
    kernel_img_mul_8[38] <= 'd0;
    kernel_img_mul_8[39] <= 'd0;
    kernel_img_mul_8[40] <= 'd0;
    kernel_img_mul_8[41] <= 'd0;
    kernel_img_mul_8[42] <= 'd0;
    kernel_img_mul_8[43] <= 'd0;
    kernel_img_mul_8[44] <= 'd0;
    kernel_img_mul_8[45] <= 'd0;
    kernel_img_mul_8[46] <= 'd0;
    kernel_img_mul_8[47] <= 'd0;
    kernel_img_mul_8[48] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_8[0] <= { {8{1'b0}},layer0[8][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_8[1] <= { {8{1'b0}},layer0[8][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_8[2] <= { {8{1'b0}},layer0[8][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_8[3] <= { {8{1'b0}},layer0[8][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_8[4] <= { {8{1'b0}},layer0[8][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_8[5] <= { {8{1'b0}},layer0[8][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_8[6] <= { {8{1'b0}},layer0[8][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
    kernel_img_mul_8[7] <= { {8{1'b0}},layer1[8][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_8[8] <= { {8{1'b0}},layer1[8][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_8[9] <= { {8{1'b0}},layer1[8][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_8[10] <= { {8{1'b0}},layer1[8][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_8[11] <= { {8{1'b0}},layer1[8][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_8[12] <= { {8{1'b0}},layer1[8][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_8[13] <= { {8{1'b0}},layer1[8][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_8[14] <= { {8{1'b0}},layer2[8][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_8[15] <= { {8{1'b0}},layer2[8][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_8[16] <= { {8{1'b0}},layer2[8][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_8[17] <= { {8{1'b0}},layer2[8][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_8[18] <= { {8{1'b0}},layer2[8][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_8[19] <= { {8{1'b0}},layer2[8][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_8[20] <= { {8{1'b0}},layer2[8][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_8[21] <= { {8{1'b0}},layer3[8][7:0]} * { {8{1'b0}}, G_Kernel_7x7_3[7:0]};
    kernel_img_mul_8[22] <= { {8{1'b0}},layer3[8][15:8]} * { {8{1'b0}}, G_Kernel_7x7_3[15:8]};
    kernel_img_mul_8[23] <= { {8{1'b0}},layer3[8][23:16]} * { {8{1'b0}}, G_Kernel_7x7_3[23:16]};
    kernel_img_mul_8[24] <= { {8{1'b0}},layer3[8][31:24]} * { {8{1'b0}}, G_Kernel_7x7_3[31:24]};
    kernel_img_mul_8[25] <= { {8{1'b0}},layer3[8][39:32]} * { {8{1'b0}}, G_Kernel_7x7_3[39:32]};
    kernel_img_mul_8[26] <= { {8{1'b0}},layer3[8][47:40]} * { {8{1'b0}}, G_Kernel_7x7_3[47:40]};
    kernel_img_mul_8[27] <= { {8{1'b0}},layer3[8][55:48]} * { {8{1'b0}}, G_Kernel_7x7_3[55:48]};
    kernel_img_mul_8[28] <= { {8{1'b0}},layer4[8][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_8[29] <= { {8{1'b0}},layer4[8][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_8[30] <= { {8{1'b0}},layer4[8][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_8[31] <= { {8{1'b0}},layer4[8][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_8[32] <= { {8{1'b0}},layer4[8][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_8[33] <= { {8{1'b0}},layer4[8][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_8[34] <= { {8{1'b0}},layer4[8][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_8[35] <= { {8{1'b0}},layer5[8][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_8[36] <= { {8{1'b0}},layer5[8][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_8[37] <= { {8{1'b0}},layer5[8][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_8[38] <= { {8{1'b0}},layer5[8][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_8[39] <= { {8{1'b0}},layer5[8][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_8[40] <= { {8{1'b0}},layer5[8][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_8[41] <= { {8{1'b0}},layer5[8][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_8[42] <= { {8{1'b0}},layer6[8][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_8[43] <= { {8{1'b0}},layer6[8][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_8[44] <= { {8{1'b0}},layer6[8][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_8[45] <= { {8{1'b0}},layer6[8][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_8[46] <= { {8{1'b0}},layer6[8][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_8[47] <= { {8{1'b0}},layer6[8][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_8[48] <= { {8{1'b0}},layer6[8][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
  end
end
reg  [15:0]  kernel_img_sum_1_8;
reg  [15:0]  kernel_img_sum_2_8;
reg  [15:0]  kernel_img_sum_3_8;
reg  [15:0]  kernel_img_sum_4_8;
reg  [15:0]  kernel_img_sum_5_8;
reg  [15:0]  kernel_img_sum_6_8;
reg  [15:0]  kernel_img_sum_7_8;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_8 <= kernel_img_mul_8[0] + kernel_img_mul_8[1] + kernel_img_mul_8[2] + kernel_img_mul_8[3] + kernel_img_mul_8[4] + kernel_img_mul_8[5] + kernel_img_mul_8[6] + kernel_img_mul_8[7] + kernel_img_mul_8[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_8 <= kernel_img_mul_8[9] + kernel_img_mul_8[10] + kernel_img_mul_8[11] + kernel_img_mul_8[12] + kernel_img_mul_8[13] + kernel_img_mul_8[14] + kernel_img_mul_8[15] + kernel_img_mul_8[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_8 <= kernel_img_mul_8[17] + kernel_img_mul_8[18] + kernel_img_mul_8[19] + kernel_img_mul_8[20] + kernel_img_mul_8[21] + kernel_img_mul_8[22] + kernel_img_mul_8[23] + kernel_img_mul_8[24];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_8 <= kernel_img_mul_8[25] + kernel_img_mul_8[26] + kernel_img_mul_8[27] + kernel_img_mul_8[28] + kernel_img_mul_8[29] + kernel_img_mul_8[30] + kernel_img_mul_8[31] + kernel_img_mul_8[32];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_8 <= kernel_img_mul_8[33] + kernel_img_mul_8[34] + kernel_img_mul_8[35] + kernel_img_mul_8[36] + kernel_img_mul_8[37] + kernel_img_mul_8[38] + kernel_img_mul_8[39] + kernel_img_mul_8[40];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_8 <= kernel_img_mul_8[41] + kernel_img_mul_8[42] + kernel_img_mul_8[43] + kernel_img_mul_8[44] + kernel_img_mul_8[45] + kernel_img_mul_8[46] + kernel_img_mul_8[47] + kernel_img_mul_8[48];
  end
end
always@(*) begin
  kernel_img_sum_7_8 = kernel_img_sum_1_8 + kernel_img_sum_2_8 + kernel_img_sum_3_8 + kernel_img_sum_4_8 + kernel_img_sum_5_8 + kernel_img_sum_6_8;
end
reg  [15:0]  kernel_img_mul_9[0:48];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_9[0] <= 'd0;
    kernel_img_mul_9[1] <= 'd0;
    kernel_img_mul_9[2] <= 'd0;
    kernel_img_mul_9[3] <= 'd0;
    kernel_img_mul_9[4] <= 'd0;
    kernel_img_mul_9[5] <= 'd0;
    kernel_img_mul_9[6] <= 'd0;
    kernel_img_mul_9[7] <= 'd0;
    kernel_img_mul_9[8] <= 'd0;
    kernel_img_mul_9[9] <= 'd0;
    kernel_img_mul_9[10] <= 'd0;
    kernel_img_mul_9[11] <= 'd0;
    kernel_img_mul_9[12] <= 'd0;
    kernel_img_mul_9[13] <= 'd0;
    kernel_img_mul_9[14] <= 'd0;
    kernel_img_mul_9[15] <= 'd0;
    kernel_img_mul_9[16] <= 'd0;
    kernel_img_mul_9[17] <= 'd0;
    kernel_img_mul_9[18] <= 'd0;
    kernel_img_mul_9[19] <= 'd0;
    kernel_img_mul_9[20] <= 'd0;
    kernel_img_mul_9[21] <= 'd0;
    kernel_img_mul_9[22] <= 'd0;
    kernel_img_mul_9[23] <= 'd0;
    kernel_img_mul_9[24] <= 'd0;
    kernel_img_mul_9[25] <= 'd0;
    kernel_img_mul_9[26] <= 'd0;
    kernel_img_mul_9[27] <= 'd0;
    kernel_img_mul_9[28] <= 'd0;
    kernel_img_mul_9[29] <= 'd0;
    kernel_img_mul_9[30] <= 'd0;
    kernel_img_mul_9[31] <= 'd0;
    kernel_img_mul_9[32] <= 'd0;
    kernel_img_mul_9[33] <= 'd0;
    kernel_img_mul_9[34] <= 'd0;
    kernel_img_mul_9[35] <= 'd0;
    kernel_img_mul_9[36] <= 'd0;
    kernel_img_mul_9[37] <= 'd0;
    kernel_img_mul_9[38] <= 'd0;
    kernel_img_mul_9[39] <= 'd0;
    kernel_img_mul_9[40] <= 'd0;
    kernel_img_mul_9[41] <= 'd0;
    kernel_img_mul_9[42] <= 'd0;
    kernel_img_mul_9[43] <= 'd0;
    kernel_img_mul_9[44] <= 'd0;
    kernel_img_mul_9[45] <= 'd0;
    kernel_img_mul_9[46] <= 'd0;
    kernel_img_mul_9[47] <= 'd0;
    kernel_img_mul_9[48] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_9[0] <= { {8{1'b0}},layer0[9][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_9[1] <= { {8{1'b0}},layer0[9][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_9[2] <= { {8{1'b0}},layer0[9][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_9[3] <= { {8{1'b0}},layer0[9][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_9[4] <= { {8{1'b0}},layer0[9][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_9[5] <= { {8{1'b0}},layer0[9][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_9[6] <= { {8{1'b0}},layer0[9][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
    kernel_img_mul_9[7] <= { {8{1'b0}},layer1[9][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_9[8] <= { {8{1'b0}},layer1[9][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_9[9] <= { {8{1'b0}},layer1[9][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_9[10] <= { {8{1'b0}},layer1[9][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_9[11] <= { {8{1'b0}},layer1[9][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_9[12] <= { {8{1'b0}},layer1[9][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_9[13] <= { {8{1'b0}},layer1[9][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_9[14] <= { {8{1'b0}},layer2[9][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_9[15] <= { {8{1'b0}},layer2[9][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_9[16] <= { {8{1'b0}},layer2[9][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_9[17] <= { {8{1'b0}},layer2[9][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_9[18] <= { {8{1'b0}},layer2[9][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_9[19] <= { {8{1'b0}},layer2[9][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_9[20] <= { {8{1'b0}},layer2[9][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_9[21] <= { {8{1'b0}},layer3[9][7:0]} * { {8{1'b0}}, G_Kernel_7x7_3[7:0]};
    kernel_img_mul_9[22] <= { {8{1'b0}},layer3[9][15:8]} * { {8{1'b0}}, G_Kernel_7x7_3[15:8]};
    kernel_img_mul_9[23] <= { {8{1'b0}},layer3[9][23:16]} * { {8{1'b0}}, G_Kernel_7x7_3[23:16]};
    kernel_img_mul_9[24] <= { {8{1'b0}},layer3[9][31:24]} * { {8{1'b0}}, G_Kernel_7x7_3[31:24]};
    kernel_img_mul_9[25] <= { {8{1'b0}},layer3[9][39:32]} * { {8{1'b0}}, G_Kernel_7x7_3[39:32]};
    kernel_img_mul_9[26] <= { {8{1'b0}},layer3[9][47:40]} * { {8{1'b0}}, G_Kernel_7x7_3[47:40]};
    kernel_img_mul_9[27] <= { {8{1'b0}},layer3[9][55:48]} * { {8{1'b0}}, G_Kernel_7x7_3[55:48]};
    kernel_img_mul_9[28] <= { {8{1'b0}},layer4[9][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_9[29] <= { {8{1'b0}},layer4[9][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_9[30] <= { {8{1'b0}},layer4[9][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_9[31] <= { {8{1'b0}},layer4[9][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_9[32] <= { {8{1'b0}},layer4[9][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_9[33] <= { {8{1'b0}},layer4[9][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_9[34] <= { {8{1'b0}},layer4[9][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_9[35] <= { {8{1'b0}},layer5[9][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_9[36] <= { {8{1'b0}},layer5[9][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_9[37] <= { {8{1'b0}},layer5[9][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_9[38] <= { {8{1'b0}},layer5[9][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_9[39] <= { {8{1'b0}},layer5[9][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_9[40] <= { {8{1'b0}},layer5[9][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_9[41] <= { {8{1'b0}},layer5[9][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_9[42] <= { {8{1'b0}},layer6[9][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_9[43] <= { {8{1'b0}},layer6[9][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_9[44] <= { {8{1'b0}},layer6[9][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_9[45] <= { {8{1'b0}},layer6[9][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_9[46] <= { {8{1'b0}},layer6[9][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_9[47] <= { {8{1'b0}},layer6[9][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_9[48] <= { {8{1'b0}},layer6[9][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
  end
end
reg  [15:0]  kernel_img_sum_1_9;
reg  [15:0]  kernel_img_sum_2_9;
reg  [15:0]  kernel_img_sum_3_9;
reg  [15:0]  kernel_img_sum_4_9;
reg  [15:0]  kernel_img_sum_5_9;
reg  [15:0]  kernel_img_sum_6_9;
reg  [15:0]  kernel_img_sum_7_9;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_9 <= kernel_img_mul_9[0] + kernel_img_mul_9[1] + kernel_img_mul_9[2] + kernel_img_mul_9[3] + kernel_img_mul_9[4] + kernel_img_mul_9[5] + kernel_img_mul_9[6] + kernel_img_mul_9[7] + kernel_img_mul_9[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_9 <= kernel_img_mul_9[9] + kernel_img_mul_9[10] + kernel_img_mul_9[11] + kernel_img_mul_9[12] + kernel_img_mul_9[13] + kernel_img_mul_9[14] + kernel_img_mul_9[15] + kernel_img_mul_9[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_9 <= kernel_img_mul_9[17] + kernel_img_mul_9[18] + kernel_img_mul_9[19] + kernel_img_mul_9[20] + kernel_img_mul_9[21] + kernel_img_mul_9[22] + kernel_img_mul_9[23] + kernel_img_mul_9[24];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_9 <= kernel_img_mul_9[25] + kernel_img_mul_9[26] + kernel_img_mul_9[27] + kernel_img_mul_9[28] + kernel_img_mul_9[29] + kernel_img_mul_9[30] + kernel_img_mul_9[31] + kernel_img_mul_9[32];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_9 <= kernel_img_mul_9[33] + kernel_img_mul_9[34] + kernel_img_mul_9[35] + kernel_img_mul_9[36] + kernel_img_mul_9[37] + kernel_img_mul_9[38] + kernel_img_mul_9[39] + kernel_img_mul_9[40];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_9 <= kernel_img_mul_9[41] + kernel_img_mul_9[42] + kernel_img_mul_9[43] + kernel_img_mul_9[44] + kernel_img_mul_9[45] + kernel_img_mul_9[46] + kernel_img_mul_9[47] + kernel_img_mul_9[48];
  end
end
always@(*) begin
  kernel_img_sum_7_9 = kernel_img_sum_1_9 + kernel_img_sum_2_9 + kernel_img_sum_3_9 + kernel_img_sum_4_9 + kernel_img_sum_5_9 + kernel_img_sum_6_9;
end
reg  [15:0]  kernel_img_mul_10[0:48];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_10[0] <= 'd0;
    kernel_img_mul_10[1] <= 'd0;
    kernel_img_mul_10[2] <= 'd0;
    kernel_img_mul_10[3] <= 'd0;
    kernel_img_mul_10[4] <= 'd0;
    kernel_img_mul_10[5] <= 'd0;
    kernel_img_mul_10[6] <= 'd0;
    kernel_img_mul_10[7] <= 'd0;
    kernel_img_mul_10[8] <= 'd0;
    kernel_img_mul_10[9] <= 'd0;
    kernel_img_mul_10[10] <= 'd0;
    kernel_img_mul_10[11] <= 'd0;
    kernel_img_mul_10[12] <= 'd0;
    kernel_img_mul_10[13] <= 'd0;
    kernel_img_mul_10[14] <= 'd0;
    kernel_img_mul_10[15] <= 'd0;
    kernel_img_mul_10[16] <= 'd0;
    kernel_img_mul_10[17] <= 'd0;
    kernel_img_mul_10[18] <= 'd0;
    kernel_img_mul_10[19] <= 'd0;
    kernel_img_mul_10[20] <= 'd0;
    kernel_img_mul_10[21] <= 'd0;
    kernel_img_mul_10[22] <= 'd0;
    kernel_img_mul_10[23] <= 'd0;
    kernel_img_mul_10[24] <= 'd0;
    kernel_img_mul_10[25] <= 'd0;
    kernel_img_mul_10[26] <= 'd0;
    kernel_img_mul_10[27] <= 'd0;
    kernel_img_mul_10[28] <= 'd0;
    kernel_img_mul_10[29] <= 'd0;
    kernel_img_mul_10[30] <= 'd0;
    kernel_img_mul_10[31] <= 'd0;
    kernel_img_mul_10[32] <= 'd0;
    kernel_img_mul_10[33] <= 'd0;
    kernel_img_mul_10[34] <= 'd0;
    kernel_img_mul_10[35] <= 'd0;
    kernel_img_mul_10[36] <= 'd0;
    kernel_img_mul_10[37] <= 'd0;
    kernel_img_mul_10[38] <= 'd0;
    kernel_img_mul_10[39] <= 'd0;
    kernel_img_mul_10[40] <= 'd0;
    kernel_img_mul_10[41] <= 'd0;
    kernel_img_mul_10[42] <= 'd0;
    kernel_img_mul_10[43] <= 'd0;
    kernel_img_mul_10[44] <= 'd0;
    kernel_img_mul_10[45] <= 'd0;
    kernel_img_mul_10[46] <= 'd0;
    kernel_img_mul_10[47] <= 'd0;
    kernel_img_mul_10[48] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_10[0] <= { {8{1'b0}},layer0[10][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_10[1] <= { {8{1'b0}},layer0[10][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_10[2] <= { {8{1'b0}},layer0[10][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_10[3] <= { {8{1'b0}},layer0[10][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_10[4] <= { {8{1'b0}},layer0[10][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_10[5] <= { {8{1'b0}},layer0[10][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_10[6] <= { {8{1'b0}},layer0[10][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
    kernel_img_mul_10[7] <= { {8{1'b0}},layer1[10][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_10[8] <= { {8{1'b0}},layer1[10][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_10[9] <= { {8{1'b0}},layer1[10][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_10[10] <= { {8{1'b0}},layer1[10][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_10[11] <= { {8{1'b0}},layer1[10][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_10[12] <= { {8{1'b0}},layer1[10][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_10[13] <= { {8{1'b0}},layer1[10][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_10[14] <= { {8{1'b0}},layer2[10][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_10[15] <= { {8{1'b0}},layer2[10][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_10[16] <= { {8{1'b0}},layer2[10][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_10[17] <= { {8{1'b0}},layer2[10][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_10[18] <= { {8{1'b0}},layer2[10][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_10[19] <= { {8{1'b0}},layer2[10][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_10[20] <= { {8{1'b0}},layer2[10][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_10[21] <= { {8{1'b0}},layer3[10][7:0]} * { {8{1'b0}}, G_Kernel_7x7_3[7:0]};
    kernel_img_mul_10[22] <= { {8{1'b0}},layer3[10][15:8]} * { {8{1'b0}}, G_Kernel_7x7_3[15:8]};
    kernel_img_mul_10[23] <= { {8{1'b0}},layer3[10][23:16]} * { {8{1'b0}}, G_Kernel_7x7_3[23:16]};
    kernel_img_mul_10[24] <= { {8{1'b0}},layer3[10][31:24]} * { {8{1'b0}}, G_Kernel_7x7_3[31:24]};
    kernel_img_mul_10[25] <= { {8{1'b0}},layer3[10][39:32]} * { {8{1'b0}}, G_Kernel_7x7_3[39:32]};
    kernel_img_mul_10[26] <= { {8{1'b0}},layer3[10][47:40]} * { {8{1'b0}}, G_Kernel_7x7_3[47:40]};
    kernel_img_mul_10[27] <= { {8{1'b0}},layer3[10][55:48]} * { {8{1'b0}}, G_Kernel_7x7_3[55:48]};
    kernel_img_mul_10[28] <= { {8{1'b0}},layer4[10][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_10[29] <= { {8{1'b0}},layer4[10][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_10[30] <= { {8{1'b0}},layer4[10][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_10[31] <= { {8{1'b0}},layer4[10][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_10[32] <= { {8{1'b0}},layer4[10][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_10[33] <= { {8{1'b0}},layer4[10][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_10[34] <= { {8{1'b0}},layer4[10][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_10[35] <= { {8{1'b0}},layer5[10][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_10[36] <= { {8{1'b0}},layer5[10][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_10[37] <= { {8{1'b0}},layer5[10][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_10[38] <= { {8{1'b0}},layer5[10][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_10[39] <= { {8{1'b0}},layer5[10][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_10[40] <= { {8{1'b0}},layer5[10][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_10[41] <= { {8{1'b0}},layer5[10][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_10[42] <= { {8{1'b0}},layer6[10][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_10[43] <= { {8{1'b0}},layer6[10][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_10[44] <= { {8{1'b0}},layer6[10][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_10[45] <= { {8{1'b0}},layer6[10][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_10[46] <= { {8{1'b0}},layer6[10][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_10[47] <= { {8{1'b0}},layer6[10][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_10[48] <= { {8{1'b0}},layer6[10][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
  end
end
reg  [15:0]  kernel_img_sum_1_10;
reg  [15:0]  kernel_img_sum_2_10;
reg  [15:0]  kernel_img_sum_3_10;
reg  [15:0]  kernel_img_sum_4_10;
reg  [15:0]  kernel_img_sum_5_10;
reg  [15:0]  kernel_img_sum_6_10;
reg  [15:0]  kernel_img_sum_7_10;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_10 <= kernel_img_mul_10[0] + kernel_img_mul_10[1] + kernel_img_mul_10[2] + kernel_img_mul_10[3] + kernel_img_mul_10[4] + kernel_img_mul_10[5] + kernel_img_mul_10[6] + kernel_img_mul_10[7] + kernel_img_mul_10[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_10 <= kernel_img_mul_10[9] + kernel_img_mul_10[10] + kernel_img_mul_10[11] + kernel_img_mul_10[12] + kernel_img_mul_10[13] + kernel_img_mul_10[14] + kernel_img_mul_10[15] + kernel_img_mul_10[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_10 <= kernel_img_mul_10[17] + kernel_img_mul_10[18] + kernel_img_mul_10[19] + kernel_img_mul_10[20] + kernel_img_mul_10[21] + kernel_img_mul_10[22] + kernel_img_mul_10[23] + kernel_img_mul_10[24];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_10 <= kernel_img_mul_10[25] + kernel_img_mul_10[26] + kernel_img_mul_10[27] + kernel_img_mul_10[28] + kernel_img_mul_10[29] + kernel_img_mul_10[30] + kernel_img_mul_10[31] + kernel_img_mul_10[32];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_10 <= kernel_img_mul_10[33] + kernel_img_mul_10[34] + kernel_img_mul_10[35] + kernel_img_mul_10[36] + kernel_img_mul_10[37] + kernel_img_mul_10[38] + kernel_img_mul_10[39] + kernel_img_mul_10[40];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_10 <= kernel_img_mul_10[41] + kernel_img_mul_10[42] + kernel_img_mul_10[43] + kernel_img_mul_10[44] + kernel_img_mul_10[45] + kernel_img_mul_10[46] + kernel_img_mul_10[47] + kernel_img_mul_10[48];
  end
end
always@(*) begin
  kernel_img_sum_7_10 = kernel_img_sum_1_10 + kernel_img_sum_2_10 + kernel_img_sum_3_10 + kernel_img_sum_4_10 + kernel_img_sum_5_10 + kernel_img_sum_6_10;
end
reg  [15:0]  kernel_img_mul_11[0:48];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_11[0] <= 'd0;
    kernel_img_mul_11[1] <= 'd0;
    kernel_img_mul_11[2] <= 'd0;
    kernel_img_mul_11[3] <= 'd0;
    kernel_img_mul_11[4] <= 'd0;
    kernel_img_mul_11[5] <= 'd0;
    kernel_img_mul_11[6] <= 'd0;
    kernel_img_mul_11[7] <= 'd0;
    kernel_img_mul_11[8] <= 'd0;
    kernel_img_mul_11[9] <= 'd0;
    kernel_img_mul_11[10] <= 'd0;
    kernel_img_mul_11[11] <= 'd0;
    kernel_img_mul_11[12] <= 'd0;
    kernel_img_mul_11[13] <= 'd0;
    kernel_img_mul_11[14] <= 'd0;
    kernel_img_mul_11[15] <= 'd0;
    kernel_img_mul_11[16] <= 'd0;
    kernel_img_mul_11[17] <= 'd0;
    kernel_img_mul_11[18] <= 'd0;
    kernel_img_mul_11[19] <= 'd0;
    kernel_img_mul_11[20] <= 'd0;
    kernel_img_mul_11[21] <= 'd0;
    kernel_img_mul_11[22] <= 'd0;
    kernel_img_mul_11[23] <= 'd0;
    kernel_img_mul_11[24] <= 'd0;
    kernel_img_mul_11[25] <= 'd0;
    kernel_img_mul_11[26] <= 'd0;
    kernel_img_mul_11[27] <= 'd0;
    kernel_img_mul_11[28] <= 'd0;
    kernel_img_mul_11[29] <= 'd0;
    kernel_img_mul_11[30] <= 'd0;
    kernel_img_mul_11[31] <= 'd0;
    kernel_img_mul_11[32] <= 'd0;
    kernel_img_mul_11[33] <= 'd0;
    kernel_img_mul_11[34] <= 'd0;
    kernel_img_mul_11[35] <= 'd0;
    kernel_img_mul_11[36] <= 'd0;
    kernel_img_mul_11[37] <= 'd0;
    kernel_img_mul_11[38] <= 'd0;
    kernel_img_mul_11[39] <= 'd0;
    kernel_img_mul_11[40] <= 'd0;
    kernel_img_mul_11[41] <= 'd0;
    kernel_img_mul_11[42] <= 'd0;
    kernel_img_mul_11[43] <= 'd0;
    kernel_img_mul_11[44] <= 'd0;
    kernel_img_mul_11[45] <= 'd0;
    kernel_img_mul_11[46] <= 'd0;
    kernel_img_mul_11[47] <= 'd0;
    kernel_img_mul_11[48] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_11[0] <= { {8{1'b0}},layer0[11][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_11[1] <= { {8{1'b0}},layer0[11][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_11[2] <= { {8{1'b0}},layer0[11][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_11[3] <= { {8{1'b0}},layer0[11][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_11[4] <= { {8{1'b0}},layer0[11][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_11[5] <= { {8{1'b0}},layer0[11][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_11[6] <= { {8{1'b0}},layer0[11][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
    kernel_img_mul_11[7] <= { {8{1'b0}},layer1[11][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_11[8] <= { {8{1'b0}},layer1[11][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_11[9] <= { {8{1'b0}},layer1[11][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_11[10] <= { {8{1'b0}},layer1[11][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_11[11] <= { {8{1'b0}},layer1[11][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_11[12] <= { {8{1'b0}},layer1[11][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_11[13] <= { {8{1'b0}},layer1[11][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_11[14] <= { {8{1'b0}},layer2[11][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_11[15] <= { {8{1'b0}},layer2[11][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_11[16] <= { {8{1'b0}},layer2[11][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_11[17] <= { {8{1'b0}},layer2[11][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_11[18] <= { {8{1'b0}},layer2[11][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_11[19] <= { {8{1'b0}},layer2[11][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_11[20] <= { {8{1'b0}},layer2[11][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_11[21] <= { {8{1'b0}},layer3[11][7:0]} * { {8{1'b0}}, G_Kernel_7x7_3[7:0]};
    kernel_img_mul_11[22] <= { {8{1'b0}},layer3[11][15:8]} * { {8{1'b0}}, G_Kernel_7x7_3[15:8]};
    kernel_img_mul_11[23] <= { {8{1'b0}},layer3[11][23:16]} * { {8{1'b0}}, G_Kernel_7x7_3[23:16]};
    kernel_img_mul_11[24] <= { {8{1'b0}},layer3[11][31:24]} * { {8{1'b0}}, G_Kernel_7x7_3[31:24]};
    kernel_img_mul_11[25] <= { {8{1'b0}},layer3[11][39:32]} * { {8{1'b0}}, G_Kernel_7x7_3[39:32]};
    kernel_img_mul_11[26] <= { {8{1'b0}},layer3[11][47:40]} * { {8{1'b0}}, G_Kernel_7x7_3[47:40]};
    kernel_img_mul_11[27] <= { {8{1'b0}},layer3[11][55:48]} * { {8{1'b0}}, G_Kernel_7x7_3[55:48]};
    kernel_img_mul_11[28] <= { {8{1'b0}},layer4[11][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_11[29] <= { {8{1'b0}},layer4[11][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_11[30] <= { {8{1'b0}},layer4[11][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_11[31] <= { {8{1'b0}},layer4[11][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_11[32] <= { {8{1'b0}},layer4[11][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_11[33] <= { {8{1'b0}},layer4[11][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_11[34] <= { {8{1'b0}},layer4[11][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_11[35] <= { {8{1'b0}},layer5[11][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_11[36] <= { {8{1'b0}},layer5[11][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_11[37] <= { {8{1'b0}},layer5[11][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_11[38] <= { {8{1'b0}},layer5[11][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_11[39] <= { {8{1'b0}},layer5[11][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_11[40] <= { {8{1'b0}},layer5[11][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_11[41] <= { {8{1'b0}},layer5[11][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_11[42] <= { {8{1'b0}},layer6[11][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_11[43] <= { {8{1'b0}},layer6[11][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_11[44] <= { {8{1'b0}},layer6[11][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_11[45] <= { {8{1'b0}},layer6[11][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_11[46] <= { {8{1'b0}},layer6[11][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_11[47] <= { {8{1'b0}},layer6[11][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_11[48] <= { {8{1'b0}},layer6[11][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
  end
end
reg  [15:0]  kernel_img_sum_1_11;
reg  [15:0]  kernel_img_sum_2_11;
reg  [15:0]  kernel_img_sum_3_11;
reg  [15:0]  kernel_img_sum_4_11;
reg  [15:0]  kernel_img_sum_5_11;
reg  [15:0]  kernel_img_sum_6_11;
reg  [15:0]  kernel_img_sum_7_11;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_11 <= kernel_img_mul_11[0] + kernel_img_mul_11[1] + kernel_img_mul_11[2] + kernel_img_mul_11[3] + kernel_img_mul_11[4] + kernel_img_mul_11[5] + kernel_img_mul_11[6] + kernel_img_mul_11[7] + kernel_img_mul_11[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_11 <= kernel_img_mul_11[9] + kernel_img_mul_11[10] + kernel_img_mul_11[11] + kernel_img_mul_11[12] + kernel_img_mul_11[13] + kernel_img_mul_11[14] + kernel_img_mul_11[15] + kernel_img_mul_11[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_11 <= kernel_img_mul_11[17] + kernel_img_mul_11[18] + kernel_img_mul_11[19] + kernel_img_mul_11[20] + kernel_img_mul_11[21] + kernel_img_mul_11[22] + kernel_img_mul_11[23] + kernel_img_mul_11[24];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_11 <= kernel_img_mul_11[25] + kernel_img_mul_11[26] + kernel_img_mul_11[27] + kernel_img_mul_11[28] + kernel_img_mul_11[29] + kernel_img_mul_11[30] + kernel_img_mul_11[31] + kernel_img_mul_11[32];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_11 <= kernel_img_mul_11[33] + kernel_img_mul_11[34] + kernel_img_mul_11[35] + kernel_img_mul_11[36] + kernel_img_mul_11[37] + kernel_img_mul_11[38] + kernel_img_mul_11[39] + kernel_img_mul_11[40];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_11 <= kernel_img_mul_11[41] + kernel_img_mul_11[42] + kernel_img_mul_11[43] + kernel_img_mul_11[44] + kernel_img_mul_11[45] + kernel_img_mul_11[46] + kernel_img_mul_11[47] + kernel_img_mul_11[48];
  end
end
always@(*) begin
  kernel_img_sum_7_11 = kernel_img_sum_1_11 + kernel_img_sum_2_11 + kernel_img_sum_3_11 + kernel_img_sum_4_11 + kernel_img_sum_5_11 + kernel_img_sum_6_11;
end
reg  [15:0]  kernel_img_mul_12[0:48];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_12[0] <= 'd0;
    kernel_img_mul_12[1] <= 'd0;
    kernel_img_mul_12[2] <= 'd0;
    kernel_img_mul_12[3] <= 'd0;
    kernel_img_mul_12[4] <= 'd0;
    kernel_img_mul_12[5] <= 'd0;
    kernel_img_mul_12[6] <= 'd0;
    kernel_img_mul_12[7] <= 'd0;
    kernel_img_mul_12[8] <= 'd0;
    kernel_img_mul_12[9] <= 'd0;
    kernel_img_mul_12[10] <= 'd0;
    kernel_img_mul_12[11] <= 'd0;
    kernel_img_mul_12[12] <= 'd0;
    kernel_img_mul_12[13] <= 'd0;
    kernel_img_mul_12[14] <= 'd0;
    kernel_img_mul_12[15] <= 'd0;
    kernel_img_mul_12[16] <= 'd0;
    kernel_img_mul_12[17] <= 'd0;
    kernel_img_mul_12[18] <= 'd0;
    kernel_img_mul_12[19] <= 'd0;
    kernel_img_mul_12[20] <= 'd0;
    kernel_img_mul_12[21] <= 'd0;
    kernel_img_mul_12[22] <= 'd0;
    kernel_img_mul_12[23] <= 'd0;
    kernel_img_mul_12[24] <= 'd0;
    kernel_img_mul_12[25] <= 'd0;
    kernel_img_mul_12[26] <= 'd0;
    kernel_img_mul_12[27] <= 'd0;
    kernel_img_mul_12[28] <= 'd0;
    kernel_img_mul_12[29] <= 'd0;
    kernel_img_mul_12[30] <= 'd0;
    kernel_img_mul_12[31] <= 'd0;
    kernel_img_mul_12[32] <= 'd0;
    kernel_img_mul_12[33] <= 'd0;
    kernel_img_mul_12[34] <= 'd0;
    kernel_img_mul_12[35] <= 'd0;
    kernel_img_mul_12[36] <= 'd0;
    kernel_img_mul_12[37] <= 'd0;
    kernel_img_mul_12[38] <= 'd0;
    kernel_img_mul_12[39] <= 'd0;
    kernel_img_mul_12[40] <= 'd0;
    kernel_img_mul_12[41] <= 'd0;
    kernel_img_mul_12[42] <= 'd0;
    kernel_img_mul_12[43] <= 'd0;
    kernel_img_mul_12[44] <= 'd0;
    kernel_img_mul_12[45] <= 'd0;
    kernel_img_mul_12[46] <= 'd0;
    kernel_img_mul_12[47] <= 'd0;
    kernel_img_mul_12[48] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_12[0] <= { {8{1'b0}},layer0[12][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_12[1] <= { {8{1'b0}},layer0[12][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_12[2] <= { {8{1'b0}},layer0[12][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_12[3] <= { {8{1'b0}},layer0[12][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_12[4] <= { {8{1'b0}},layer0[12][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_12[5] <= { {8{1'b0}},layer0[12][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_12[6] <= { {8{1'b0}},layer0[12][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
    kernel_img_mul_12[7] <= { {8{1'b0}},layer1[12][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_12[8] <= { {8{1'b0}},layer1[12][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_12[9] <= { {8{1'b0}},layer1[12][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_12[10] <= { {8{1'b0}},layer1[12][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_12[11] <= { {8{1'b0}},layer1[12][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_12[12] <= { {8{1'b0}},layer1[12][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_12[13] <= { {8{1'b0}},layer1[12][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_12[14] <= { {8{1'b0}},layer2[12][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_12[15] <= { {8{1'b0}},layer2[12][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_12[16] <= { {8{1'b0}},layer2[12][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_12[17] <= { {8{1'b0}},layer2[12][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_12[18] <= { {8{1'b0}},layer2[12][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_12[19] <= { {8{1'b0}},layer2[12][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_12[20] <= { {8{1'b0}},layer2[12][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_12[21] <= { {8{1'b0}},layer3[12][7:0]} * { {8{1'b0}}, G_Kernel_7x7_3[7:0]};
    kernel_img_mul_12[22] <= { {8{1'b0}},layer3[12][15:8]} * { {8{1'b0}}, G_Kernel_7x7_3[15:8]};
    kernel_img_mul_12[23] <= { {8{1'b0}},layer3[12][23:16]} * { {8{1'b0}}, G_Kernel_7x7_3[23:16]};
    kernel_img_mul_12[24] <= { {8{1'b0}},layer3[12][31:24]} * { {8{1'b0}}, G_Kernel_7x7_3[31:24]};
    kernel_img_mul_12[25] <= { {8{1'b0}},layer3[12][39:32]} * { {8{1'b0}}, G_Kernel_7x7_3[39:32]};
    kernel_img_mul_12[26] <= { {8{1'b0}},layer3[12][47:40]} * { {8{1'b0}}, G_Kernel_7x7_3[47:40]};
    kernel_img_mul_12[27] <= { {8{1'b0}},layer3[12][55:48]} * { {8{1'b0}}, G_Kernel_7x7_3[55:48]};
    kernel_img_mul_12[28] <= { {8{1'b0}},layer4[12][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_12[29] <= { {8{1'b0}},layer4[12][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_12[30] <= { {8{1'b0}},layer4[12][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_12[31] <= { {8{1'b0}},layer4[12][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_12[32] <= { {8{1'b0}},layer4[12][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_12[33] <= { {8{1'b0}},layer4[12][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_12[34] <= { {8{1'b0}},layer4[12][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_12[35] <= { {8{1'b0}},layer5[12][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_12[36] <= { {8{1'b0}},layer5[12][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_12[37] <= { {8{1'b0}},layer5[12][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_12[38] <= { {8{1'b0}},layer5[12][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_12[39] <= { {8{1'b0}},layer5[12][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_12[40] <= { {8{1'b0}},layer5[12][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_12[41] <= { {8{1'b0}},layer5[12][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_12[42] <= { {8{1'b0}},layer6[12][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_12[43] <= { {8{1'b0}},layer6[12][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_12[44] <= { {8{1'b0}},layer6[12][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_12[45] <= { {8{1'b0}},layer6[12][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_12[46] <= { {8{1'b0}},layer6[12][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_12[47] <= { {8{1'b0}},layer6[12][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_12[48] <= { {8{1'b0}},layer6[12][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
  end
end
reg  [15:0]  kernel_img_sum_1_12;
reg  [15:0]  kernel_img_sum_2_12;
reg  [15:0]  kernel_img_sum_3_12;
reg  [15:0]  kernel_img_sum_4_12;
reg  [15:0]  kernel_img_sum_5_12;
reg  [15:0]  kernel_img_sum_6_12;
reg  [15:0]  kernel_img_sum_7_12;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_12 <= kernel_img_mul_12[0] + kernel_img_mul_12[1] + kernel_img_mul_12[2] + kernel_img_mul_12[3] + kernel_img_mul_12[4] + kernel_img_mul_12[5] + kernel_img_mul_12[6] + kernel_img_mul_12[7] + kernel_img_mul_12[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_12 <= kernel_img_mul_12[9] + kernel_img_mul_12[10] + kernel_img_mul_12[11] + kernel_img_mul_12[12] + kernel_img_mul_12[13] + kernel_img_mul_12[14] + kernel_img_mul_12[15] + kernel_img_mul_12[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_12 <= kernel_img_mul_12[17] + kernel_img_mul_12[18] + kernel_img_mul_12[19] + kernel_img_mul_12[20] + kernel_img_mul_12[21] + kernel_img_mul_12[22] + kernel_img_mul_12[23] + kernel_img_mul_12[24];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_12 <= kernel_img_mul_12[25] + kernel_img_mul_12[26] + kernel_img_mul_12[27] + kernel_img_mul_12[28] + kernel_img_mul_12[29] + kernel_img_mul_12[30] + kernel_img_mul_12[31] + kernel_img_mul_12[32];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_12 <= kernel_img_mul_12[33] + kernel_img_mul_12[34] + kernel_img_mul_12[35] + kernel_img_mul_12[36] + kernel_img_mul_12[37] + kernel_img_mul_12[38] + kernel_img_mul_12[39] + kernel_img_mul_12[40];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_12 <= kernel_img_mul_12[41] + kernel_img_mul_12[42] + kernel_img_mul_12[43] + kernel_img_mul_12[44] + kernel_img_mul_12[45] + kernel_img_mul_12[46] + kernel_img_mul_12[47] + kernel_img_mul_12[48];
  end
end
always@(*) begin
  kernel_img_sum_7_12 = kernel_img_sum_1_12 + kernel_img_sum_2_12 + kernel_img_sum_3_12 + kernel_img_sum_4_12 + kernel_img_sum_5_12 + kernel_img_sum_6_12;
end
reg  [15:0]  kernel_img_mul_13[0:48];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_13[0] <= 'd0;
    kernel_img_mul_13[1] <= 'd0;
    kernel_img_mul_13[2] <= 'd0;
    kernel_img_mul_13[3] <= 'd0;
    kernel_img_mul_13[4] <= 'd0;
    kernel_img_mul_13[5] <= 'd0;
    kernel_img_mul_13[6] <= 'd0;
    kernel_img_mul_13[7] <= 'd0;
    kernel_img_mul_13[8] <= 'd0;
    kernel_img_mul_13[9] <= 'd0;
    kernel_img_mul_13[10] <= 'd0;
    kernel_img_mul_13[11] <= 'd0;
    kernel_img_mul_13[12] <= 'd0;
    kernel_img_mul_13[13] <= 'd0;
    kernel_img_mul_13[14] <= 'd0;
    kernel_img_mul_13[15] <= 'd0;
    kernel_img_mul_13[16] <= 'd0;
    kernel_img_mul_13[17] <= 'd0;
    kernel_img_mul_13[18] <= 'd0;
    kernel_img_mul_13[19] <= 'd0;
    kernel_img_mul_13[20] <= 'd0;
    kernel_img_mul_13[21] <= 'd0;
    kernel_img_mul_13[22] <= 'd0;
    kernel_img_mul_13[23] <= 'd0;
    kernel_img_mul_13[24] <= 'd0;
    kernel_img_mul_13[25] <= 'd0;
    kernel_img_mul_13[26] <= 'd0;
    kernel_img_mul_13[27] <= 'd0;
    kernel_img_mul_13[28] <= 'd0;
    kernel_img_mul_13[29] <= 'd0;
    kernel_img_mul_13[30] <= 'd0;
    kernel_img_mul_13[31] <= 'd0;
    kernel_img_mul_13[32] <= 'd0;
    kernel_img_mul_13[33] <= 'd0;
    kernel_img_mul_13[34] <= 'd0;
    kernel_img_mul_13[35] <= 'd0;
    kernel_img_mul_13[36] <= 'd0;
    kernel_img_mul_13[37] <= 'd0;
    kernel_img_mul_13[38] <= 'd0;
    kernel_img_mul_13[39] <= 'd0;
    kernel_img_mul_13[40] <= 'd0;
    kernel_img_mul_13[41] <= 'd0;
    kernel_img_mul_13[42] <= 'd0;
    kernel_img_mul_13[43] <= 'd0;
    kernel_img_mul_13[44] <= 'd0;
    kernel_img_mul_13[45] <= 'd0;
    kernel_img_mul_13[46] <= 'd0;
    kernel_img_mul_13[47] <= 'd0;
    kernel_img_mul_13[48] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_13[0] <= { {8{1'b0}},layer0[13][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_13[1] <= { {8{1'b0}},layer0[13][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_13[2] <= { {8{1'b0}},layer0[13][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_13[3] <= { {8{1'b0}},layer0[13][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_13[4] <= { {8{1'b0}},layer0[13][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_13[5] <= { {8{1'b0}},layer0[13][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_13[6] <= { {8{1'b0}},layer0[13][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
    kernel_img_mul_13[7] <= { {8{1'b0}},layer1[13][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_13[8] <= { {8{1'b0}},layer1[13][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_13[9] <= { {8{1'b0}},layer1[13][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_13[10] <= { {8{1'b0}},layer1[13][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_13[11] <= { {8{1'b0}},layer1[13][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_13[12] <= { {8{1'b0}},layer1[13][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_13[13] <= { {8{1'b0}},layer1[13][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_13[14] <= { {8{1'b0}},layer2[13][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_13[15] <= { {8{1'b0}},layer2[13][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_13[16] <= { {8{1'b0}},layer2[13][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_13[17] <= { {8{1'b0}},layer2[13][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_13[18] <= { {8{1'b0}},layer2[13][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_13[19] <= { {8{1'b0}},layer2[13][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_13[20] <= { {8{1'b0}},layer2[13][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_13[21] <= { {8{1'b0}},layer3[13][7:0]} * { {8{1'b0}}, G_Kernel_7x7_3[7:0]};
    kernel_img_mul_13[22] <= { {8{1'b0}},layer3[13][15:8]} * { {8{1'b0}}, G_Kernel_7x7_3[15:8]};
    kernel_img_mul_13[23] <= { {8{1'b0}},layer3[13][23:16]} * { {8{1'b0}}, G_Kernel_7x7_3[23:16]};
    kernel_img_mul_13[24] <= { {8{1'b0}},layer3[13][31:24]} * { {8{1'b0}}, G_Kernel_7x7_3[31:24]};
    kernel_img_mul_13[25] <= { {8{1'b0}},layer3[13][39:32]} * { {8{1'b0}}, G_Kernel_7x7_3[39:32]};
    kernel_img_mul_13[26] <= { {8{1'b0}},layer3[13][47:40]} * { {8{1'b0}}, G_Kernel_7x7_3[47:40]};
    kernel_img_mul_13[27] <= { {8{1'b0}},layer3[13][55:48]} * { {8{1'b0}}, G_Kernel_7x7_3[55:48]};
    kernel_img_mul_13[28] <= { {8{1'b0}},layer4[13][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_13[29] <= { {8{1'b0}},layer4[13][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_13[30] <= { {8{1'b0}},layer4[13][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_13[31] <= { {8{1'b0}},layer4[13][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_13[32] <= { {8{1'b0}},layer4[13][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_13[33] <= { {8{1'b0}},layer4[13][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_13[34] <= { {8{1'b0}},layer4[13][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_13[35] <= { {8{1'b0}},layer5[13][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_13[36] <= { {8{1'b0}},layer5[13][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_13[37] <= { {8{1'b0}},layer5[13][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_13[38] <= { {8{1'b0}},layer5[13][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_13[39] <= { {8{1'b0}},layer5[13][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_13[40] <= { {8{1'b0}},layer5[13][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_13[41] <= { {8{1'b0}},layer5[13][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_13[42] <= { {8{1'b0}},layer6[13][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_13[43] <= { {8{1'b0}},layer6[13][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_13[44] <= { {8{1'b0}},layer6[13][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_13[45] <= { {8{1'b0}},layer6[13][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_13[46] <= { {8{1'b0}},layer6[13][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_13[47] <= { {8{1'b0}},layer6[13][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_13[48] <= { {8{1'b0}},layer6[13][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
  end
end
reg  [15:0]  kernel_img_sum_1_13;
reg  [15:0]  kernel_img_sum_2_13;
reg  [15:0]  kernel_img_sum_3_13;
reg  [15:0]  kernel_img_sum_4_13;
reg  [15:0]  kernel_img_sum_5_13;
reg  [15:0]  kernel_img_sum_6_13;
reg  [15:0]  kernel_img_sum_7_13;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_13 <= kernel_img_mul_13[0] + kernel_img_mul_13[1] + kernel_img_mul_13[2] + kernel_img_mul_13[3] + kernel_img_mul_13[4] + kernel_img_mul_13[5] + kernel_img_mul_13[6] + kernel_img_mul_13[7] + kernel_img_mul_13[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_13 <= kernel_img_mul_13[9] + kernel_img_mul_13[10] + kernel_img_mul_13[11] + kernel_img_mul_13[12] + kernel_img_mul_13[13] + kernel_img_mul_13[14] + kernel_img_mul_13[15] + kernel_img_mul_13[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_13 <= kernel_img_mul_13[17] + kernel_img_mul_13[18] + kernel_img_mul_13[19] + kernel_img_mul_13[20] + kernel_img_mul_13[21] + kernel_img_mul_13[22] + kernel_img_mul_13[23] + kernel_img_mul_13[24];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_13 <= kernel_img_mul_13[25] + kernel_img_mul_13[26] + kernel_img_mul_13[27] + kernel_img_mul_13[28] + kernel_img_mul_13[29] + kernel_img_mul_13[30] + kernel_img_mul_13[31] + kernel_img_mul_13[32];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_13 <= kernel_img_mul_13[33] + kernel_img_mul_13[34] + kernel_img_mul_13[35] + kernel_img_mul_13[36] + kernel_img_mul_13[37] + kernel_img_mul_13[38] + kernel_img_mul_13[39] + kernel_img_mul_13[40];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_13 <= kernel_img_mul_13[41] + kernel_img_mul_13[42] + kernel_img_mul_13[43] + kernel_img_mul_13[44] + kernel_img_mul_13[45] + kernel_img_mul_13[46] + kernel_img_mul_13[47] + kernel_img_mul_13[48];
  end
end
always@(*) begin
  kernel_img_sum_7_13 = kernel_img_sum_1_13 + kernel_img_sum_2_13 + kernel_img_sum_3_13 + kernel_img_sum_4_13 + kernel_img_sum_5_13 + kernel_img_sum_6_13;
end
reg  [15:0]  kernel_img_mul_14[0:48];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_14[0] <= 'd0;
    kernel_img_mul_14[1] <= 'd0;
    kernel_img_mul_14[2] <= 'd0;
    kernel_img_mul_14[3] <= 'd0;
    kernel_img_mul_14[4] <= 'd0;
    kernel_img_mul_14[5] <= 'd0;
    kernel_img_mul_14[6] <= 'd0;
    kernel_img_mul_14[7] <= 'd0;
    kernel_img_mul_14[8] <= 'd0;
    kernel_img_mul_14[9] <= 'd0;
    kernel_img_mul_14[10] <= 'd0;
    kernel_img_mul_14[11] <= 'd0;
    kernel_img_mul_14[12] <= 'd0;
    kernel_img_mul_14[13] <= 'd0;
    kernel_img_mul_14[14] <= 'd0;
    kernel_img_mul_14[15] <= 'd0;
    kernel_img_mul_14[16] <= 'd0;
    kernel_img_mul_14[17] <= 'd0;
    kernel_img_mul_14[18] <= 'd0;
    kernel_img_mul_14[19] <= 'd0;
    kernel_img_mul_14[20] <= 'd0;
    kernel_img_mul_14[21] <= 'd0;
    kernel_img_mul_14[22] <= 'd0;
    kernel_img_mul_14[23] <= 'd0;
    kernel_img_mul_14[24] <= 'd0;
    kernel_img_mul_14[25] <= 'd0;
    kernel_img_mul_14[26] <= 'd0;
    kernel_img_mul_14[27] <= 'd0;
    kernel_img_mul_14[28] <= 'd0;
    kernel_img_mul_14[29] <= 'd0;
    kernel_img_mul_14[30] <= 'd0;
    kernel_img_mul_14[31] <= 'd0;
    kernel_img_mul_14[32] <= 'd0;
    kernel_img_mul_14[33] <= 'd0;
    kernel_img_mul_14[34] <= 'd0;
    kernel_img_mul_14[35] <= 'd0;
    kernel_img_mul_14[36] <= 'd0;
    kernel_img_mul_14[37] <= 'd0;
    kernel_img_mul_14[38] <= 'd0;
    kernel_img_mul_14[39] <= 'd0;
    kernel_img_mul_14[40] <= 'd0;
    kernel_img_mul_14[41] <= 'd0;
    kernel_img_mul_14[42] <= 'd0;
    kernel_img_mul_14[43] <= 'd0;
    kernel_img_mul_14[44] <= 'd0;
    kernel_img_mul_14[45] <= 'd0;
    kernel_img_mul_14[46] <= 'd0;
    kernel_img_mul_14[47] <= 'd0;
    kernel_img_mul_14[48] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_14[0] <= { {8{1'b0}},layer0[14][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_14[1] <= { {8{1'b0}},layer0[14][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_14[2] <= { {8{1'b0}},layer0[14][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_14[3] <= { {8{1'b0}},layer0[14][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_14[4] <= { {8{1'b0}},layer0[14][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_14[5] <= { {8{1'b0}},layer0[14][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_14[6] <= { {8{1'b0}},layer0[14][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
    kernel_img_mul_14[7] <= { {8{1'b0}},layer1[14][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_14[8] <= { {8{1'b0}},layer1[14][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_14[9] <= { {8{1'b0}},layer1[14][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_14[10] <= { {8{1'b0}},layer1[14][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_14[11] <= { {8{1'b0}},layer1[14][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_14[12] <= { {8{1'b0}},layer1[14][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_14[13] <= { {8{1'b0}},layer1[14][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_14[14] <= { {8{1'b0}},layer2[14][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_14[15] <= { {8{1'b0}},layer2[14][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_14[16] <= { {8{1'b0}},layer2[14][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_14[17] <= { {8{1'b0}},layer2[14][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_14[18] <= { {8{1'b0}},layer2[14][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_14[19] <= { {8{1'b0}},layer2[14][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_14[20] <= { {8{1'b0}},layer2[14][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_14[21] <= { {8{1'b0}},layer3[14][7:0]} * { {8{1'b0}}, G_Kernel_7x7_3[7:0]};
    kernel_img_mul_14[22] <= { {8{1'b0}},layer3[14][15:8]} * { {8{1'b0}}, G_Kernel_7x7_3[15:8]};
    kernel_img_mul_14[23] <= { {8{1'b0}},layer3[14][23:16]} * { {8{1'b0}}, G_Kernel_7x7_3[23:16]};
    kernel_img_mul_14[24] <= { {8{1'b0}},layer3[14][31:24]} * { {8{1'b0}}, G_Kernel_7x7_3[31:24]};
    kernel_img_mul_14[25] <= { {8{1'b0}},layer3[14][39:32]} * { {8{1'b0}}, G_Kernel_7x7_3[39:32]};
    kernel_img_mul_14[26] <= { {8{1'b0}},layer3[14][47:40]} * { {8{1'b0}}, G_Kernel_7x7_3[47:40]};
    kernel_img_mul_14[27] <= { {8{1'b0}},layer3[14][55:48]} * { {8{1'b0}}, G_Kernel_7x7_3[55:48]};
    kernel_img_mul_14[28] <= { {8{1'b0}},layer4[14][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_14[29] <= { {8{1'b0}},layer4[14][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_14[30] <= { {8{1'b0}},layer4[14][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_14[31] <= { {8{1'b0}},layer4[14][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_14[32] <= { {8{1'b0}},layer4[14][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_14[33] <= { {8{1'b0}},layer4[14][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_14[34] <= { {8{1'b0}},layer4[14][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_14[35] <= { {8{1'b0}},layer5[14][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_14[36] <= { {8{1'b0}},layer5[14][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_14[37] <= { {8{1'b0}},layer5[14][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_14[38] <= { {8{1'b0}},layer5[14][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_14[39] <= { {8{1'b0}},layer5[14][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_14[40] <= { {8{1'b0}},layer5[14][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_14[41] <= { {8{1'b0}},layer5[14][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_14[42] <= { {8{1'b0}},layer6[14][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_14[43] <= { {8{1'b0}},layer6[14][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_14[44] <= { {8{1'b0}},layer6[14][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_14[45] <= { {8{1'b0}},layer6[14][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_14[46] <= { {8{1'b0}},layer6[14][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_14[47] <= { {8{1'b0}},layer6[14][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_14[48] <= { {8{1'b0}},layer6[14][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
  end
end
reg  [15:0]  kernel_img_sum_1_14;
reg  [15:0]  kernel_img_sum_2_14;
reg  [15:0]  kernel_img_sum_3_14;
reg  [15:0]  kernel_img_sum_4_14;
reg  [15:0]  kernel_img_sum_5_14;
reg  [15:0]  kernel_img_sum_6_14;
reg  [15:0]  kernel_img_sum_7_14;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_14 <= kernel_img_mul_14[0] + kernel_img_mul_14[1] + kernel_img_mul_14[2] + kernel_img_mul_14[3] + kernel_img_mul_14[4] + kernel_img_mul_14[5] + kernel_img_mul_14[6] + kernel_img_mul_14[7] + kernel_img_mul_14[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_14 <= kernel_img_mul_14[9] + kernel_img_mul_14[10] + kernel_img_mul_14[11] + kernel_img_mul_14[12] + kernel_img_mul_14[13] + kernel_img_mul_14[14] + kernel_img_mul_14[15] + kernel_img_mul_14[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_14 <= kernel_img_mul_14[17] + kernel_img_mul_14[18] + kernel_img_mul_14[19] + kernel_img_mul_14[20] + kernel_img_mul_14[21] + kernel_img_mul_14[22] + kernel_img_mul_14[23] + kernel_img_mul_14[24];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_14 <= kernel_img_mul_14[25] + kernel_img_mul_14[26] + kernel_img_mul_14[27] + kernel_img_mul_14[28] + kernel_img_mul_14[29] + kernel_img_mul_14[30] + kernel_img_mul_14[31] + kernel_img_mul_14[32];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_14 <= kernel_img_mul_14[33] + kernel_img_mul_14[34] + kernel_img_mul_14[35] + kernel_img_mul_14[36] + kernel_img_mul_14[37] + kernel_img_mul_14[38] + kernel_img_mul_14[39] + kernel_img_mul_14[40];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_14 <= kernel_img_mul_14[41] + kernel_img_mul_14[42] + kernel_img_mul_14[43] + kernel_img_mul_14[44] + kernel_img_mul_14[45] + kernel_img_mul_14[46] + kernel_img_mul_14[47] + kernel_img_mul_14[48];
  end
end
always@(*) begin
  kernel_img_sum_7_14 = kernel_img_sum_1_14 + kernel_img_sum_2_14 + kernel_img_sum_3_14 + kernel_img_sum_4_14 + kernel_img_sum_5_14 + kernel_img_sum_6_14;
end
reg  [15:0]  kernel_img_mul_15[0:48];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_15[0] <= 'd0;
    kernel_img_mul_15[1] <= 'd0;
    kernel_img_mul_15[2] <= 'd0;
    kernel_img_mul_15[3] <= 'd0;
    kernel_img_mul_15[4] <= 'd0;
    kernel_img_mul_15[5] <= 'd0;
    kernel_img_mul_15[6] <= 'd0;
    kernel_img_mul_15[7] <= 'd0;
    kernel_img_mul_15[8] <= 'd0;
    kernel_img_mul_15[9] <= 'd0;
    kernel_img_mul_15[10] <= 'd0;
    kernel_img_mul_15[11] <= 'd0;
    kernel_img_mul_15[12] <= 'd0;
    kernel_img_mul_15[13] <= 'd0;
    kernel_img_mul_15[14] <= 'd0;
    kernel_img_mul_15[15] <= 'd0;
    kernel_img_mul_15[16] <= 'd0;
    kernel_img_mul_15[17] <= 'd0;
    kernel_img_mul_15[18] <= 'd0;
    kernel_img_mul_15[19] <= 'd0;
    kernel_img_mul_15[20] <= 'd0;
    kernel_img_mul_15[21] <= 'd0;
    kernel_img_mul_15[22] <= 'd0;
    kernel_img_mul_15[23] <= 'd0;
    kernel_img_mul_15[24] <= 'd0;
    kernel_img_mul_15[25] <= 'd0;
    kernel_img_mul_15[26] <= 'd0;
    kernel_img_mul_15[27] <= 'd0;
    kernel_img_mul_15[28] <= 'd0;
    kernel_img_mul_15[29] <= 'd0;
    kernel_img_mul_15[30] <= 'd0;
    kernel_img_mul_15[31] <= 'd0;
    kernel_img_mul_15[32] <= 'd0;
    kernel_img_mul_15[33] <= 'd0;
    kernel_img_mul_15[34] <= 'd0;
    kernel_img_mul_15[35] <= 'd0;
    kernel_img_mul_15[36] <= 'd0;
    kernel_img_mul_15[37] <= 'd0;
    kernel_img_mul_15[38] <= 'd0;
    kernel_img_mul_15[39] <= 'd0;
    kernel_img_mul_15[40] <= 'd0;
    kernel_img_mul_15[41] <= 'd0;
    kernel_img_mul_15[42] <= 'd0;
    kernel_img_mul_15[43] <= 'd0;
    kernel_img_mul_15[44] <= 'd0;
    kernel_img_mul_15[45] <= 'd0;
    kernel_img_mul_15[46] <= 'd0;
    kernel_img_mul_15[47] <= 'd0;
    kernel_img_mul_15[48] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_15[0] <= { {8{1'b0}},layer0[15][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_15[1] <= { {8{1'b0}},layer0[15][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_15[2] <= { {8{1'b0}},layer0[15][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_15[3] <= { {8{1'b0}},layer0[15][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_15[4] <= { {8{1'b0}},layer0[15][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_15[5] <= { {8{1'b0}},layer0[15][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_15[6] <= { {8{1'b0}},layer0[15][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
    kernel_img_mul_15[7] <= { {8{1'b0}},layer1[15][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_15[8] <= { {8{1'b0}},layer1[15][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_15[9] <= { {8{1'b0}},layer1[15][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_15[10] <= { {8{1'b0}},layer1[15][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_15[11] <= { {8{1'b0}},layer1[15][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_15[12] <= { {8{1'b0}},layer1[15][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_15[13] <= { {8{1'b0}},layer1[15][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_15[14] <= { {8{1'b0}},layer2[15][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_15[15] <= { {8{1'b0}},layer2[15][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_15[16] <= { {8{1'b0}},layer2[15][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_15[17] <= { {8{1'b0}},layer2[15][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_15[18] <= { {8{1'b0}},layer2[15][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_15[19] <= { {8{1'b0}},layer2[15][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_15[20] <= { {8{1'b0}},layer2[15][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_15[21] <= { {8{1'b0}},layer3[15][7:0]} * { {8{1'b0}}, G_Kernel_7x7_3[7:0]};
    kernel_img_mul_15[22] <= { {8{1'b0}},layer3[15][15:8]} * { {8{1'b0}}, G_Kernel_7x7_3[15:8]};
    kernel_img_mul_15[23] <= { {8{1'b0}},layer3[15][23:16]} * { {8{1'b0}}, G_Kernel_7x7_3[23:16]};
    kernel_img_mul_15[24] <= { {8{1'b0}},layer3[15][31:24]} * { {8{1'b0}}, G_Kernel_7x7_3[31:24]};
    kernel_img_mul_15[25] <= { {8{1'b0}},layer3[15][39:32]} * { {8{1'b0}}, G_Kernel_7x7_3[39:32]};
    kernel_img_mul_15[26] <= { {8{1'b0}},layer3[15][47:40]} * { {8{1'b0}}, G_Kernel_7x7_3[47:40]};
    kernel_img_mul_15[27] <= { {8{1'b0}},layer3[15][55:48]} * { {8{1'b0}}, G_Kernel_7x7_3[55:48]};
    kernel_img_mul_15[28] <= { {8{1'b0}},layer4[15][7:0]} * { {8{1'b0}}, G_Kernel_7x7_2[7:0]};
    kernel_img_mul_15[29] <= { {8{1'b0}},layer4[15][15:8]} * { {8{1'b0}}, G_Kernel_7x7_2[15:8]};
    kernel_img_mul_15[30] <= { {8{1'b0}},layer4[15][23:16]} * { {8{1'b0}}, G_Kernel_7x7_2[23:16]};
    kernel_img_mul_15[31] <= { {8{1'b0}},layer4[15][31:24]} * { {8{1'b0}}, G_Kernel_7x7_2[31:24]};
    kernel_img_mul_15[32] <= { {8{1'b0}},layer4[15][39:32]} * { {8{1'b0}}, G_Kernel_7x7_2[39:32]};
    kernel_img_mul_15[33] <= { {8{1'b0}},layer4[15][47:40]} * { {8{1'b0}}, G_Kernel_7x7_2[47:40]};
    kernel_img_mul_15[34] <= { {8{1'b0}},layer4[15][55:48]} * { {8{1'b0}}, G_Kernel_7x7_2[55:48]};
    kernel_img_mul_15[35] <= { {8{1'b0}},layer5[15][7:0]} * { {8{1'b0}}, G_Kernel_7x7_1[7:0]};
    kernel_img_mul_15[36] <= { {8{1'b0}},layer5[15][15:8]} * { {8{1'b0}}, G_Kernel_7x7_1[15:8]};
    kernel_img_mul_15[37] <= { {8{1'b0}},layer5[15][23:16]} * { {8{1'b0}}, G_Kernel_7x7_1[23:16]};
    kernel_img_mul_15[38] <= { {8{1'b0}},layer5[15][31:24]} * { {8{1'b0}}, G_Kernel_7x7_1[31:24]};
    kernel_img_mul_15[39] <= { {8{1'b0}},layer5[15][39:32]} * { {8{1'b0}}, G_Kernel_7x7_1[39:32]};
    kernel_img_mul_15[40] <= { {8{1'b0}},layer5[15][47:40]} * { {8{1'b0}}, G_Kernel_7x7_1[47:40]};
    kernel_img_mul_15[41] <= { {8{1'b0}},layer5[15][55:48]} * { {8{1'b0}}, G_Kernel_7x7_1[55:48]};
    kernel_img_mul_15[42] <= { {8{1'b0}},layer6[15][7:0]} * { {8{1'b0}}, G_Kernel_7x7_0[7:0]};
    kernel_img_mul_15[43] <= { {8{1'b0}},layer6[15][15:8]} * { {8{1'b0}}, G_Kernel_7x7_0[15:8]};
    kernel_img_mul_15[44] <= { {8{1'b0}},layer6[15][23:16]} * { {8{1'b0}}, G_Kernel_7x7_0[23:16]};
    kernel_img_mul_15[45] <= { {8{1'b0}},layer6[15][31:24]} * { {8{1'b0}}, G_Kernel_7x7_0[31:24]};
    kernel_img_mul_15[46] <= { {8{1'b0}},layer6[15][39:32]} * { {8{1'b0}}, G_Kernel_7x7_0[39:32]};
    kernel_img_mul_15[47] <= { {8{1'b0}},layer6[15][47:40]} * { {8{1'b0}}, G_Kernel_7x7_0[47:40]};
    kernel_img_mul_15[48] <= { {8{1'b0}},layer6[15][55:48]} * { {8{1'b0}}, G_Kernel_7x7_0[55:48]};
  end
end
reg  [15:0]  kernel_img_sum_1_15;
reg  [15:0]  kernel_img_sum_2_15;
reg  [15:0]  kernel_img_sum_3_15;
reg  [15:0]  kernel_img_sum_4_15;
reg  [15:0]  kernel_img_sum_5_15;
reg  [15:0]  kernel_img_sum_6_15;
reg  [15:0]  kernel_img_sum_7_15;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_15 <= kernel_img_mul_15[0] + kernel_img_mul_15[1] + kernel_img_mul_15[2] + kernel_img_mul_15[3] + kernel_img_mul_15[4] + kernel_img_mul_15[5] + kernel_img_mul_15[6] + kernel_img_mul_15[7] + kernel_img_mul_15[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_15 <= kernel_img_mul_15[9] + kernel_img_mul_15[10] + kernel_img_mul_15[11] + kernel_img_mul_15[12] + kernel_img_mul_15[13] + kernel_img_mul_15[14] + kernel_img_mul_15[15] + kernel_img_mul_15[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_15 <= kernel_img_mul_15[17] + kernel_img_mul_15[18] + kernel_img_mul_15[19] + kernel_img_mul_15[20] + kernel_img_mul_15[21] + kernel_img_mul_15[22] + kernel_img_mul_15[23] + kernel_img_mul_15[24];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_15 <= kernel_img_mul_15[25] + kernel_img_mul_15[26] + kernel_img_mul_15[27] + kernel_img_mul_15[28] + kernel_img_mul_15[29] + kernel_img_mul_15[30] + kernel_img_mul_15[31] + kernel_img_mul_15[32];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_15 <= kernel_img_mul_15[33] + kernel_img_mul_15[34] + kernel_img_mul_15[35] + kernel_img_mul_15[36] + kernel_img_mul_15[37] + kernel_img_mul_15[38] + kernel_img_mul_15[39] + kernel_img_mul_15[40];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_15 <= kernel_img_mul_15[41] + kernel_img_mul_15[42] + kernel_img_mul_15[43] + kernel_img_mul_15[44] + kernel_img_mul_15[45] + kernel_img_mul_15[46] + kernel_img_mul_15[47] + kernel_img_mul_15[48];
  end
end
always@(*) begin
  kernel_img_sum_7_15 = kernel_img_sum_1_15 + kernel_img_sum_2_15 + kernel_img_sum_3_15 + kernel_img_sum_4_15 + kernel_img_sum_5_15 + kernel_img_sum_6_15;
end
always @(posedge clk) begin
  if(!rst_n) begin
    blur_out[7:0] <= 'd0;
    blur_out[15:8] <= 'd0;
    blur_out[23:16] <= 'd0;
    blur_out[31:24] <= 'd0;
    blur_out[39:32] <= 'd0;
    blur_out[47:40] <= 'd0;
    blur_out[55:48] <= 'd0;
    blur_out[63:56] <= 'd0;
    blur_out[71:64] <= 'd0;
    blur_out[79:72] <= 'd0;
    blur_out[87:80] <= 'd0;
    blur_out[95:88] <= 'd0;
    blur_out[103:96] <= 'd0;
    blur_out[111:104] <= 'd0;
    blur_out[119:112] <= 'd0;
    blur_out[127:120] <= 'd0;
  end
  else if(current_state==ST_UPDATE) begin
    blur_out[7:0] <= kernel_img_sum_7_0[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[15:8] <= kernel_img_sum_7_1[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[23:16] <= kernel_img_sum_7_2[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[31:24] <= kernel_img_sum_7_3[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[39:32] <= kernel_img_sum_7_4[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[47:40] <= kernel_img_sum_7_5[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[55:48] <= kernel_img_sum_7_6[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[63:56] <= kernel_img_sum_7_7[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[71:64] <= kernel_img_sum_7_8[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[79:72] <= kernel_img_sum_7_9[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[87:80] <= kernel_img_sum_7_10[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[95:88] <= kernel_img_sum_7_11[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[103:96] <= kernel_img_sum_7_12[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[111:104] <= kernel_img_sum_7_13[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[119:112] <= kernel_img_sum_7_14[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[127:120] <= kernel_img_sum_7_15[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
  end
end

/*
 *  FSM
 *
 */
always @(posedge clk) begin
  if (!rst_n) begin
    current_state <= ST_MUX;    
  end
  else begin
    current_state <= next_state;
  end
end
always @(*) begin
  case(current_state)
    ST_MUX: begin
      if(start)
        next_state = ST_MUL;
      else
        next_state = ST_MUX;
    end
    ST_MUL: begin
      if(current_state==ST_MUL)
        next_state = ST_ADD;
      else 
        next_state = ST_MUL;
    end
    ST_ADD: begin
      if(current_state==ST_ADD)
        next_state = ST_UPDATE;
      else 
        next_state = ST_ADD;
    end
    ST_UPDATE: begin
      if(current_state==ST_UPDATE)
        next_state = ST_MUL;
      else 
        next_state = ST_UPDATE;
    end
    default:
      next_state = ST_MUL;
  endcase
end

endmodule