module Gaussian_Blur_5x5_1(
  clk,
  rst_n,
  buffer_data_0,
  buffer_data_1,
  buffer_data_2,
  buffer_data_3,
  buffer_data_4,
  current_col,
  blur_out,
  start,
  done
);

input                 clk;
input                 rst_n;
input                 start;
output                done;
input         [5:0]   current_col;
input       [175:0]   buffer_data_0;
input       [175:0]   buffer_data_1;
input       [175:0]   buffer_data_2;
input       [175:0]   buffer_data_3;
input       [175:0]   buffer_data_4;
output reg  [127:0]   blur_out; // wire

parameter  ST_MUX         = 0,
           ST_MUL         = 1,
           ST_ADD         = 2,
           ST_UPDATE      = 3;
reg     [2:0] current_state,
              next_state;
assign done = (current_state==ST_UPDATE) ? 1 : 0;

wire       [39:0]  G_Kernel_5x5_0;
wire       [39:0]  G_Kernel_5x5_1;
wire       [39:0]  G_Kernel_5x5_2;
assign  G_Kernel_5x5_0[7:0]   = 8'h07; //E31AF6; //18'b000001111110001100;//'d030809;
assign  G_Kernel_5x5_0[15:8]  = 8'h09; //83EB80; //18'b000010011000001111;//'d037169;
assign  G_Kernel_5x5_0[23:16] = 8'h0A; //212B91; //18'b000010100010000100;//'d039568;
assign  G_Kernel_5x5_0[31:24] = 8'h09; //83EB80; //18'b000010011000001111;//'d037169;
assign  G_Kernel_5x5_0[39:32] = 8'h07; //E31AF6; //18'b000001111110001100;//'d030809;
assign  G_Kernel_5x5_1[7:0]   = 8'h09; //83EB80; //18'b000010011000001111;//'d037169;
assign  G_Kernel_5x5_1[15:8]  = 8'h0B; //7AC7A0; //18'b000010110111101011;//'d044842;
assign  G_Kernel_5x5_1[23:16] = 8'h0C; //387DF7; //18'b000011000011100001;//'d047737;
assign  G_Kernel_5x5_1[31:24] = 8'h0B; //7AC7A0; //18'b000010110111101011;//'d044842;
assign  G_Kernel_5x5_1[39:32] = 8'h09; //83EB80; //18'b000010011000001111;//'d037169;
assign  G_Kernel_5x5_2[7:0]   = 8'h0A; //212B91; //18'b000010100010000100;//'d039568;
assign  G_Kernel_5x5_2[15:8]  = 8'h0C; //387DF7; //18'b000011000011100001;//'d047737;
assign  G_Kernel_5x5_2[23:16] = 8'h0D; //02737E; //18'b000011010000001001;//'d050818;
assign  G_Kernel_5x5_2[31:24] = 8'h0C; //387DF7; //18'b000011000011100001;//'d047737;
assign  G_Kernel_5x5_2[39:32] = 8'h0A; //212B91; //18'b000010100010000100;//'d039568;

reg    [39:0]    layer0_0;
reg    [39:0]    layer0_1;
reg    [39:0]    layer0_2;
reg    [39:0]    layer0_3;
reg    [39:0]    layer0_4;
reg    [39:0]    layer0_5;
reg    [39:0]    layer0_6;
reg    [39:0]    layer0_7;
reg    [39:0]    layer0_8;
reg    [39:0]    layer0_9;
reg    [39:0]    layer0_10;
reg    [39:0]    layer0_11;
reg    [39:0]    layer0_12;
reg    [39:0]    layer0_13;
reg    [39:0]    layer0_14;
reg    [39:0]    layer0_15;
reg    [39:0]    layer1_0;
reg    [39:0]    layer1_1;
reg    [39:0]    layer1_2;
reg    [39:0]    layer1_3;
reg    [39:0]    layer1_4;
reg    [39:0]    layer1_5;
reg    [39:0]    layer1_6;
reg    [39:0]    layer1_7;
reg    [39:0]    layer1_8;
reg    [39:0]    layer1_9;
reg    [39:0]    layer1_10;
reg    [39:0]    layer1_11;
reg    [39:0]    layer1_12;
reg    [39:0]    layer1_13;
reg    [39:0]    layer1_14;
reg    [39:0]    layer1_15;
reg    [39:0]    layer2_0;
reg    [39:0]    layer2_1;
reg    [39:0]    layer2_2;
reg    [39:0]    layer2_3;
reg    [39:0]    layer2_4;
reg    [39:0]    layer2_5;
reg    [39:0]    layer2_6;
reg    [39:0]    layer2_7;
reg    [39:0]    layer2_8;
reg    [39:0]    layer2_9;
reg    [39:0]    layer2_10;
reg    [39:0]    layer2_11;
reg    [39:0]    layer2_12;
reg    [39:0]    layer2_13;
reg    [39:0]    layer2_14;
reg    [39:0]    layer2_15;
reg    [39:0]    layer3_0;
reg    [39:0]    layer3_1;
reg    [39:0]    layer3_2;
reg    [39:0]    layer3_3;
reg    [39:0]    layer3_4;
reg    [39:0]    layer3_5;
reg    [39:0]    layer3_6;
reg    [39:0]    layer3_7;
reg    [39:0]    layer3_8;
reg    [39:0]    layer3_9;
reg    [39:0]    layer3_10;
reg    [39:0]    layer3_11;
reg    [39:0]    layer3_12;
reg    [39:0]    layer3_13;
reg    [39:0]    layer3_14;
reg    [39:0]    layer3_15;
reg    [39:0]    layer4_0;
reg    [39:0]    layer4_1;
reg    [39:0]    layer4_2;
reg    [39:0]    layer4_3;
reg    [39:0]    layer4_4;
reg    [39:0]    layer4_5;
reg    [39:0]    layer4_6;
reg    [39:0]    layer4_7;
reg    [39:0]    layer4_8;
reg    [39:0]    layer4_9;
reg    [39:0]    layer4_10;
reg    [39:0]    layer4_11;
reg    [39:0]    layer4_12;
reg    [39:0]    layer4_13;
reg    [39:0]    layer4_14;
reg    [39:0]    layer4_15;
always @(*) begin
  case(current_col)
    'd0: begin
        layer0_0[7:0] = 0;
        layer0_0[15:8] = 0;
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = 0;
        layer1_0[15:8] = 0;
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = 0;
        layer2_0[15:8] = 0;
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = 0;
        layer3_0[15:8] = 0;
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = 0;
        layer4_0[15:8] = 0;
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = 0;
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = 0;
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = 0;
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = 0;
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = 0;
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd1: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd2: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd3: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd4: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd5: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd6: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd7: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd8: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd9: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd10: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd11: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd12: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd13: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd14: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd15: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd16: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd17: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd18: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd19: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd20: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd21: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd22: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd23: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd24: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd25: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd26: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd27: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd28: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd29: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd30: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd31: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd32: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd33: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd34: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd35: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd36: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd37: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd38: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = buffer_data_4[159:152];
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = buffer_data_3[159:152];
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = buffer_data_2[159:152];
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = buffer_data_1[159:152];
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = buffer_data_0[159:152];
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = buffer_data_4[159:152];
        layer0_15[39:32] = buffer_data_4[167:160];
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = buffer_data_3[159:152];
        layer1_15[39:32] = buffer_data_3[167:160];
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = buffer_data_2[159:152];
        layer2_15[39:32] = buffer_data_2[167:160];
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = buffer_data_1[159:152];
        layer3_15[39:32] = buffer_data_1[167:160];
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = buffer_data_0[159:152];
        layer4_15[39:32] = buffer_data_0[167:160];
    end
    'd39: begin
        layer0_0[7:0] = buffer_data_4[15:8];
        layer0_0[15:8] = buffer_data_4[23:16];
        layer0_0[23:16] = buffer_data_4[31:24];
        layer0_0[31:24] = buffer_data_4[39:32];
        layer0_0[39:32] = buffer_data_4[47:40];
        layer1_0[7:0] = buffer_data_3[15:8];
        layer1_0[15:8] = buffer_data_3[23:16];
        layer1_0[23:16] = buffer_data_3[31:24];
        layer1_0[31:24] = buffer_data_3[39:32];
        layer1_0[39:32] = buffer_data_3[47:40];
        layer2_0[7:0] = buffer_data_2[15:8];
        layer2_0[15:8] = buffer_data_2[23:16];
        layer2_0[23:16] = buffer_data_2[31:24];
        layer2_0[31:24] = buffer_data_2[39:32];
        layer2_0[39:32] = buffer_data_2[47:40];
        layer3_0[7:0] = buffer_data_1[15:8];
        layer3_0[15:8] = buffer_data_1[23:16];
        layer3_0[23:16] = buffer_data_1[31:24];
        layer3_0[31:24] = buffer_data_1[39:32];
        layer3_0[39:32] = buffer_data_1[47:40];
        layer4_0[7:0] = buffer_data_0[15:8];
        layer4_0[15:8] = buffer_data_0[23:16];
        layer4_0[23:16] = buffer_data_0[31:24];
        layer4_0[31:24] = buffer_data_0[39:32];
        layer4_0[39:32] = buffer_data_0[47:40];
        layer0_1[7:0] = buffer_data_4[23:16];
        layer0_1[15:8] = buffer_data_4[31:24];
        layer0_1[23:16] = buffer_data_4[39:32];
        layer0_1[31:24] = buffer_data_4[47:40];
        layer0_1[39:32] = buffer_data_4[55:48];
        layer1_1[7:0] = buffer_data_3[23:16];
        layer1_1[15:8] = buffer_data_3[31:24];
        layer1_1[23:16] = buffer_data_3[39:32];
        layer1_1[31:24] = buffer_data_3[47:40];
        layer1_1[39:32] = buffer_data_3[55:48];
        layer2_1[7:0] = buffer_data_2[23:16];
        layer2_1[15:8] = buffer_data_2[31:24];
        layer2_1[23:16] = buffer_data_2[39:32];
        layer2_1[31:24] = buffer_data_2[47:40];
        layer2_1[39:32] = buffer_data_2[55:48];
        layer3_1[7:0] = buffer_data_1[23:16];
        layer3_1[15:8] = buffer_data_1[31:24];
        layer3_1[23:16] = buffer_data_1[39:32];
        layer3_1[31:24] = buffer_data_1[47:40];
        layer3_1[39:32] = buffer_data_1[55:48];
        layer4_1[7:0] = buffer_data_0[23:16];
        layer4_1[15:8] = buffer_data_0[31:24];
        layer4_1[23:16] = buffer_data_0[39:32];
        layer4_1[31:24] = buffer_data_0[47:40];
        layer4_1[39:32] = buffer_data_0[55:48];
        layer0_2[7:0] = buffer_data_4[31:24];
        layer0_2[15:8] = buffer_data_4[39:32];
        layer0_2[23:16] = buffer_data_4[47:40];
        layer0_2[31:24] = buffer_data_4[55:48];
        layer0_2[39:32] = buffer_data_4[63:56];
        layer1_2[7:0] = buffer_data_3[31:24];
        layer1_2[15:8] = buffer_data_3[39:32];
        layer1_2[23:16] = buffer_data_3[47:40];
        layer1_2[31:24] = buffer_data_3[55:48];
        layer1_2[39:32] = buffer_data_3[63:56];
        layer2_2[7:0] = buffer_data_2[31:24];
        layer2_2[15:8] = buffer_data_2[39:32];
        layer2_2[23:16] = buffer_data_2[47:40];
        layer2_2[31:24] = buffer_data_2[55:48];
        layer2_2[39:32] = buffer_data_2[63:56];
        layer3_2[7:0] = buffer_data_1[31:24];
        layer3_2[15:8] = buffer_data_1[39:32];
        layer3_2[23:16] = buffer_data_1[47:40];
        layer3_2[31:24] = buffer_data_1[55:48];
        layer3_2[39:32] = buffer_data_1[63:56];
        layer4_2[7:0] = buffer_data_0[31:24];
        layer4_2[15:8] = buffer_data_0[39:32];
        layer4_2[23:16] = buffer_data_0[47:40];
        layer4_2[31:24] = buffer_data_0[55:48];
        layer4_2[39:32] = buffer_data_0[63:56];
        layer0_3[7:0] = buffer_data_4[39:32];
        layer0_3[15:8] = buffer_data_4[47:40];
        layer0_3[23:16] = buffer_data_4[55:48];
        layer0_3[31:24] = buffer_data_4[63:56];
        layer0_3[39:32] = buffer_data_4[71:64];
        layer1_3[7:0] = buffer_data_3[39:32];
        layer1_3[15:8] = buffer_data_3[47:40];
        layer1_3[23:16] = buffer_data_3[55:48];
        layer1_3[31:24] = buffer_data_3[63:56];
        layer1_3[39:32] = buffer_data_3[71:64];
        layer2_3[7:0] = buffer_data_2[39:32];
        layer2_3[15:8] = buffer_data_2[47:40];
        layer2_3[23:16] = buffer_data_2[55:48];
        layer2_3[31:24] = buffer_data_2[63:56];
        layer2_3[39:32] = buffer_data_2[71:64];
        layer3_3[7:0] = buffer_data_1[39:32];
        layer3_3[15:8] = buffer_data_1[47:40];
        layer3_3[23:16] = buffer_data_1[55:48];
        layer3_3[31:24] = buffer_data_1[63:56];
        layer3_3[39:32] = buffer_data_1[71:64];
        layer4_3[7:0] = buffer_data_0[39:32];
        layer4_3[15:8] = buffer_data_0[47:40];
        layer4_3[23:16] = buffer_data_0[55:48];
        layer4_3[31:24] = buffer_data_0[63:56];
        layer4_3[39:32] = buffer_data_0[71:64];
        layer0_4[7:0] = buffer_data_4[47:40];
        layer0_4[15:8] = buffer_data_4[55:48];
        layer0_4[23:16] = buffer_data_4[63:56];
        layer0_4[31:24] = buffer_data_4[71:64];
        layer0_4[39:32] = buffer_data_4[79:72];
        layer1_4[7:0] = buffer_data_3[47:40];
        layer1_4[15:8] = buffer_data_3[55:48];
        layer1_4[23:16] = buffer_data_3[63:56];
        layer1_4[31:24] = buffer_data_3[71:64];
        layer1_4[39:32] = buffer_data_3[79:72];
        layer2_4[7:0] = buffer_data_2[47:40];
        layer2_4[15:8] = buffer_data_2[55:48];
        layer2_4[23:16] = buffer_data_2[63:56];
        layer2_4[31:24] = buffer_data_2[71:64];
        layer2_4[39:32] = buffer_data_2[79:72];
        layer3_4[7:0] = buffer_data_1[47:40];
        layer3_4[15:8] = buffer_data_1[55:48];
        layer3_4[23:16] = buffer_data_1[63:56];
        layer3_4[31:24] = buffer_data_1[71:64];
        layer3_4[39:32] = buffer_data_1[79:72];
        layer4_4[7:0] = buffer_data_0[47:40];
        layer4_4[15:8] = buffer_data_0[55:48];
        layer4_4[23:16] = buffer_data_0[63:56];
        layer4_4[31:24] = buffer_data_0[71:64];
        layer4_4[39:32] = buffer_data_0[79:72];
        layer0_5[7:0] = buffer_data_4[55:48];
        layer0_5[15:8] = buffer_data_4[63:56];
        layer0_5[23:16] = buffer_data_4[71:64];
        layer0_5[31:24] = buffer_data_4[79:72];
        layer0_5[39:32] = buffer_data_4[87:80];
        layer1_5[7:0] = buffer_data_3[55:48];
        layer1_5[15:8] = buffer_data_3[63:56];
        layer1_5[23:16] = buffer_data_3[71:64];
        layer1_5[31:24] = buffer_data_3[79:72];
        layer1_5[39:32] = buffer_data_3[87:80];
        layer2_5[7:0] = buffer_data_2[55:48];
        layer2_5[15:8] = buffer_data_2[63:56];
        layer2_5[23:16] = buffer_data_2[71:64];
        layer2_5[31:24] = buffer_data_2[79:72];
        layer2_5[39:32] = buffer_data_2[87:80];
        layer3_5[7:0] = buffer_data_1[55:48];
        layer3_5[15:8] = buffer_data_1[63:56];
        layer3_5[23:16] = buffer_data_1[71:64];
        layer3_5[31:24] = buffer_data_1[79:72];
        layer3_5[39:32] = buffer_data_1[87:80];
        layer4_5[7:0] = buffer_data_0[55:48];
        layer4_5[15:8] = buffer_data_0[63:56];
        layer4_5[23:16] = buffer_data_0[71:64];
        layer4_5[31:24] = buffer_data_0[79:72];
        layer4_5[39:32] = buffer_data_0[87:80];
        layer0_6[7:0] = buffer_data_4[63:56];
        layer0_6[15:8] = buffer_data_4[71:64];
        layer0_6[23:16] = buffer_data_4[79:72];
        layer0_6[31:24] = buffer_data_4[87:80];
        layer0_6[39:32] = buffer_data_4[95:88];
        layer1_6[7:0] = buffer_data_3[63:56];
        layer1_6[15:8] = buffer_data_3[71:64];
        layer1_6[23:16] = buffer_data_3[79:72];
        layer1_6[31:24] = buffer_data_3[87:80];
        layer1_6[39:32] = buffer_data_3[95:88];
        layer2_6[7:0] = buffer_data_2[63:56];
        layer2_6[15:8] = buffer_data_2[71:64];
        layer2_6[23:16] = buffer_data_2[79:72];
        layer2_6[31:24] = buffer_data_2[87:80];
        layer2_6[39:32] = buffer_data_2[95:88];
        layer3_6[7:0] = buffer_data_1[63:56];
        layer3_6[15:8] = buffer_data_1[71:64];
        layer3_6[23:16] = buffer_data_1[79:72];
        layer3_6[31:24] = buffer_data_1[87:80];
        layer3_6[39:32] = buffer_data_1[95:88];
        layer4_6[7:0] = buffer_data_0[63:56];
        layer4_6[15:8] = buffer_data_0[71:64];
        layer4_6[23:16] = buffer_data_0[79:72];
        layer4_6[31:24] = buffer_data_0[87:80];
        layer4_6[39:32] = buffer_data_0[95:88];
        layer0_7[7:0] = buffer_data_4[71:64];
        layer0_7[15:8] = buffer_data_4[79:72];
        layer0_7[23:16] = buffer_data_4[87:80];
        layer0_7[31:24] = buffer_data_4[95:88];
        layer0_7[39:32] = buffer_data_4[103:96];
        layer1_7[7:0] = buffer_data_3[71:64];
        layer1_7[15:8] = buffer_data_3[79:72];
        layer1_7[23:16] = buffer_data_3[87:80];
        layer1_7[31:24] = buffer_data_3[95:88];
        layer1_7[39:32] = buffer_data_3[103:96];
        layer2_7[7:0] = buffer_data_2[71:64];
        layer2_7[15:8] = buffer_data_2[79:72];
        layer2_7[23:16] = buffer_data_2[87:80];
        layer2_7[31:24] = buffer_data_2[95:88];
        layer2_7[39:32] = buffer_data_2[103:96];
        layer3_7[7:0] = buffer_data_1[71:64];
        layer3_7[15:8] = buffer_data_1[79:72];
        layer3_7[23:16] = buffer_data_1[87:80];
        layer3_7[31:24] = buffer_data_1[95:88];
        layer3_7[39:32] = buffer_data_1[103:96];
        layer4_7[7:0] = buffer_data_0[71:64];
        layer4_7[15:8] = buffer_data_0[79:72];
        layer4_7[23:16] = buffer_data_0[87:80];
        layer4_7[31:24] = buffer_data_0[95:88];
        layer4_7[39:32] = buffer_data_0[103:96];
        layer0_8[7:0] = buffer_data_4[79:72];
        layer0_8[15:8] = buffer_data_4[87:80];
        layer0_8[23:16] = buffer_data_4[95:88];
        layer0_8[31:24] = buffer_data_4[103:96];
        layer0_8[39:32] = buffer_data_4[111:104];
        layer1_8[7:0] = buffer_data_3[79:72];
        layer1_8[15:8] = buffer_data_3[87:80];
        layer1_8[23:16] = buffer_data_3[95:88];
        layer1_8[31:24] = buffer_data_3[103:96];
        layer1_8[39:32] = buffer_data_3[111:104];
        layer2_8[7:0] = buffer_data_2[79:72];
        layer2_8[15:8] = buffer_data_2[87:80];
        layer2_8[23:16] = buffer_data_2[95:88];
        layer2_8[31:24] = buffer_data_2[103:96];
        layer2_8[39:32] = buffer_data_2[111:104];
        layer3_8[7:0] = buffer_data_1[79:72];
        layer3_8[15:8] = buffer_data_1[87:80];
        layer3_8[23:16] = buffer_data_1[95:88];
        layer3_8[31:24] = buffer_data_1[103:96];
        layer3_8[39:32] = buffer_data_1[111:104];
        layer4_8[7:0] = buffer_data_0[79:72];
        layer4_8[15:8] = buffer_data_0[87:80];
        layer4_8[23:16] = buffer_data_0[95:88];
        layer4_8[31:24] = buffer_data_0[103:96];
        layer4_8[39:32] = buffer_data_0[111:104];
        layer0_9[7:0] = buffer_data_4[87:80];
        layer0_9[15:8] = buffer_data_4[95:88];
        layer0_9[23:16] = buffer_data_4[103:96];
        layer0_9[31:24] = buffer_data_4[111:104];
        layer0_9[39:32] = buffer_data_4[119:112];
        layer1_9[7:0] = buffer_data_3[87:80];
        layer1_9[15:8] = buffer_data_3[95:88];
        layer1_9[23:16] = buffer_data_3[103:96];
        layer1_9[31:24] = buffer_data_3[111:104];
        layer1_9[39:32] = buffer_data_3[119:112];
        layer2_9[7:0] = buffer_data_2[87:80];
        layer2_9[15:8] = buffer_data_2[95:88];
        layer2_9[23:16] = buffer_data_2[103:96];
        layer2_9[31:24] = buffer_data_2[111:104];
        layer2_9[39:32] = buffer_data_2[119:112];
        layer3_9[7:0] = buffer_data_1[87:80];
        layer3_9[15:8] = buffer_data_1[95:88];
        layer3_9[23:16] = buffer_data_1[103:96];
        layer3_9[31:24] = buffer_data_1[111:104];
        layer3_9[39:32] = buffer_data_1[119:112];
        layer4_9[7:0] = buffer_data_0[87:80];
        layer4_9[15:8] = buffer_data_0[95:88];
        layer4_9[23:16] = buffer_data_0[103:96];
        layer4_9[31:24] = buffer_data_0[111:104];
        layer4_9[39:32] = buffer_data_0[119:112];
        layer0_10[7:0] = buffer_data_4[95:88];
        layer0_10[15:8] = buffer_data_4[103:96];
        layer0_10[23:16] = buffer_data_4[111:104];
        layer0_10[31:24] = buffer_data_4[119:112];
        layer0_10[39:32] = buffer_data_4[127:120];
        layer1_10[7:0] = buffer_data_3[95:88];
        layer1_10[15:8] = buffer_data_3[103:96];
        layer1_10[23:16] = buffer_data_3[111:104];
        layer1_10[31:24] = buffer_data_3[119:112];
        layer1_10[39:32] = buffer_data_3[127:120];
        layer2_10[7:0] = buffer_data_2[95:88];
        layer2_10[15:8] = buffer_data_2[103:96];
        layer2_10[23:16] = buffer_data_2[111:104];
        layer2_10[31:24] = buffer_data_2[119:112];
        layer2_10[39:32] = buffer_data_2[127:120];
        layer3_10[7:0] = buffer_data_1[95:88];
        layer3_10[15:8] = buffer_data_1[103:96];
        layer3_10[23:16] = buffer_data_1[111:104];
        layer3_10[31:24] = buffer_data_1[119:112];
        layer3_10[39:32] = buffer_data_1[127:120];
        layer4_10[7:0] = buffer_data_0[95:88];
        layer4_10[15:8] = buffer_data_0[103:96];
        layer4_10[23:16] = buffer_data_0[111:104];
        layer4_10[31:24] = buffer_data_0[119:112];
        layer4_10[39:32] = buffer_data_0[127:120];
        layer0_11[7:0] = buffer_data_4[103:96];
        layer0_11[15:8] = buffer_data_4[111:104];
        layer0_11[23:16] = buffer_data_4[119:112];
        layer0_11[31:24] = buffer_data_4[127:120];
        layer0_11[39:32] = buffer_data_4[135:128];
        layer1_11[7:0] = buffer_data_3[103:96];
        layer1_11[15:8] = buffer_data_3[111:104];
        layer1_11[23:16] = buffer_data_3[119:112];
        layer1_11[31:24] = buffer_data_3[127:120];
        layer1_11[39:32] = buffer_data_3[135:128];
        layer2_11[7:0] = buffer_data_2[103:96];
        layer2_11[15:8] = buffer_data_2[111:104];
        layer2_11[23:16] = buffer_data_2[119:112];
        layer2_11[31:24] = buffer_data_2[127:120];
        layer2_11[39:32] = buffer_data_2[135:128];
        layer3_11[7:0] = buffer_data_1[103:96];
        layer3_11[15:8] = buffer_data_1[111:104];
        layer3_11[23:16] = buffer_data_1[119:112];
        layer3_11[31:24] = buffer_data_1[127:120];
        layer3_11[39:32] = buffer_data_1[135:128];
        layer4_11[7:0] = buffer_data_0[103:96];
        layer4_11[15:8] = buffer_data_0[111:104];
        layer4_11[23:16] = buffer_data_0[119:112];
        layer4_11[31:24] = buffer_data_0[127:120];
        layer4_11[39:32] = buffer_data_0[135:128];
        layer0_12[7:0] = buffer_data_4[111:104];
        layer0_12[15:8] = buffer_data_4[119:112];
        layer0_12[23:16] = buffer_data_4[127:120];
        layer0_12[31:24] = buffer_data_4[135:128];
        layer0_12[39:32] = buffer_data_4[143:136];
        layer1_12[7:0] = buffer_data_3[111:104];
        layer1_12[15:8] = buffer_data_3[119:112];
        layer1_12[23:16] = buffer_data_3[127:120];
        layer1_12[31:24] = buffer_data_3[135:128];
        layer1_12[39:32] = buffer_data_3[143:136];
        layer2_12[7:0] = buffer_data_2[111:104];
        layer2_12[15:8] = buffer_data_2[119:112];
        layer2_12[23:16] = buffer_data_2[127:120];
        layer2_12[31:24] = buffer_data_2[135:128];
        layer2_12[39:32] = buffer_data_2[143:136];
        layer3_12[7:0] = buffer_data_1[111:104];
        layer3_12[15:8] = buffer_data_1[119:112];
        layer3_12[23:16] = buffer_data_1[127:120];
        layer3_12[31:24] = buffer_data_1[135:128];
        layer3_12[39:32] = buffer_data_1[143:136];
        layer4_12[7:0] = buffer_data_0[111:104];
        layer4_12[15:8] = buffer_data_0[119:112];
        layer4_12[23:16] = buffer_data_0[127:120];
        layer4_12[31:24] = buffer_data_0[135:128];
        layer4_12[39:32] = buffer_data_0[143:136];
        layer0_13[7:0] = buffer_data_4[119:112];
        layer0_13[15:8] = buffer_data_4[127:120];
        layer0_13[23:16] = buffer_data_4[135:128];
        layer0_13[31:24] = buffer_data_4[143:136];
        layer0_13[39:32] = buffer_data_4[151:144];
        layer1_13[7:0] = buffer_data_3[119:112];
        layer1_13[15:8] = buffer_data_3[127:120];
        layer1_13[23:16] = buffer_data_3[135:128];
        layer1_13[31:24] = buffer_data_3[143:136];
        layer1_13[39:32] = buffer_data_3[151:144];
        layer2_13[7:0] = buffer_data_2[119:112];
        layer2_13[15:8] = buffer_data_2[127:120];
        layer2_13[23:16] = buffer_data_2[135:128];
        layer2_13[31:24] = buffer_data_2[143:136];
        layer2_13[39:32] = buffer_data_2[151:144];
        layer3_13[7:0] = buffer_data_1[119:112];
        layer3_13[15:8] = buffer_data_1[127:120];
        layer3_13[23:16] = buffer_data_1[135:128];
        layer3_13[31:24] = buffer_data_1[143:136];
        layer3_13[39:32] = buffer_data_1[151:144];
        layer4_13[7:0] = buffer_data_0[119:112];
        layer4_13[15:8] = buffer_data_0[127:120];
        layer4_13[23:16] = buffer_data_0[135:128];
        layer4_13[31:24] = buffer_data_0[143:136];
        layer4_13[39:32] = buffer_data_0[151:144];
        layer0_14[7:0] = buffer_data_4[127:120];
        layer0_14[15:8] = buffer_data_4[135:128];
        layer0_14[23:16] = buffer_data_4[143:136];
        layer0_14[31:24] = buffer_data_4[151:144];
        layer0_14[39:32] = 0;
        layer1_14[7:0] = buffer_data_3[127:120];
        layer1_14[15:8] = buffer_data_3[135:128];
        layer1_14[23:16] = buffer_data_3[143:136];
        layer1_14[31:24] = buffer_data_3[151:144];
        layer1_14[39:32] = 0;
        layer2_14[7:0] = buffer_data_2[127:120];
        layer2_14[15:8] = buffer_data_2[135:128];
        layer2_14[23:16] = buffer_data_2[143:136];
        layer2_14[31:24] = buffer_data_2[151:144];
        layer2_14[39:32] = 0;
        layer3_14[7:0] = buffer_data_1[127:120];
        layer3_14[15:8] = buffer_data_1[135:128];
        layer3_14[23:16] = buffer_data_1[143:136];
        layer3_14[31:24] = buffer_data_1[151:144];
        layer3_14[39:32] = 0;
        layer4_14[7:0] = buffer_data_0[127:120];
        layer4_14[15:8] = buffer_data_0[135:128];
        layer4_14[23:16] = buffer_data_0[143:136];
        layer4_14[31:24] = buffer_data_0[151:144];
        layer4_14[39:32] = 0;
        layer0_15[7:0] = buffer_data_4[135:128];
        layer0_15[15:8] = buffer_data_4[143:136];
        layer0_15[23:16] = buffer_data_4[151:144];
        layer0_15[31:24] = 0;
        layer0_15[39:32] = 0;
        layer1_15[7:0] = buffer_data_3[135:128];
        layer1_15[15:8] = buffer_data_3[143:136];
        layer1_15[23:16] = buffer_data_3[151:144];
        layer1_15[31:24] = 0;
        layer1_15[39:32] = 0;
        layer2_15[7:0] = buffer_data_2[135:128];
        layer2_15[15:8] = buffer_data_2[143:136];
        layer2_15[23:16] = buffer_data_2[151:144];
        layer2_15[31:24] = 0;
        layer2_15[39:32] = 0;
        layer3_15[7:0] = buffer_data_1[135:128];
        layer3_15[15:8] = buffer_data_1[143:136];
        layer3_15[23:16] = buffer_data_1[151:144];
        layer3_15[31:24] = 0;
        layer3_15[39:32] = 0;
        layer4_15[7:0] = buffer_data_0[135:128];
        layer4_15[15:8] = buffer_data_0[143:136];
        layer4_15[23:16] = buffer_data_0[151:144];
        layer4_15[31:24] = 0;
        layer4_15[39:32] = 0;
    end
    default: begin
        layer0_0[7:0] = 'd0;
        layer0_0[15:8] = 'd0;
        layer0_0[23:16] = 'd0;
        layer0_0[31:24] = 'd0;
        layer0_0[39:32] = 'd0;
        layer1_0[7:0] = 'd0;
        layer1_0[15:8] = 'd0;
        layer1_0[23:16] = 'd0;
        layer1_0[31:24] = 'd0;
        layer1_0[39:32] = 'd0;
        layer2_0[7:0] = 'd0;
        layer2_0[15:8] = 'd0;
        layer2_0[23:16] = 'd0;
        layer2_0[31:24] = 'd0;
        layer2_0[39:32] = 'd0;
        layer3_0[7:0] = 'd0;
        layer3_0[15:8] = 'd0;
        layer3_0[23:16] = 'd0;
        layer3_0[31:24] = 'd0;
        layer3_0[39:32] = 'd0;
        layer4_0[7:0] = 'd0;
        layer4_0[15:8] = 'd0;
        layer4_0[23:16] = 'd0;
        layer4_0[31:24] = 'd0;
        layer4_0[39:32] = 'd0;
        layer0_1[7:0] = 'd0;
        layer0_1[15:8] = 'd0;
        layer0_1[23:16] = 'd0;
        layer0_1[31:24] = 'd0;
        layer0_1[39:32] = 'd0;
        layer1_1[7:0] = 'd0;
        layer1_1[15:8] = 'd0;
        layer1_1[23:16] = 'd0;
        layer1_1[31:24] = 'd0;
        layer1_1[39:32] = 'd0;
        layer2_1[7:0] = 'd0;
        layer2_1[15:8] = 'd0;
        layer2_1[23:16] = 'd0;
        layer2_1[31:24] = 'd0;
        layer2_1[39:32] = 'd0;
        layer3_1[7:0] = 'd0;
        layer3_1[15:8] = 'd0;
        layer3_1[23:16] = 'd0;
        layer3_1[31:24] = 'd0;
        layer3_1[39:32] = 'd0;
        layer4_1[7:0] = 'd0;
        layer4_1[15:8] = 'd0;
        layer4_1[23:16] = 'd0;
        layer4_1[31:24] = 'd0;
        layer4_1[39:32] = 'd0;
        layer0_2[7:0] = 'd0;
        layer0_2[15:8] = 'd0;
        layer0_2[23:16] = 'd0;
        layer0_2[31:24] = 'd0;
        layer0_2[39:32] = 'd0;
        layer1_2[7:0] = 'd0;
        layer1_2[15:8] = 'd0;
        layer1_2[23:16] = 'd0;
        layer1_2[31:24] = 'd0;
        layer1_2[39:32] = 'd0;
        layer2_2[7:0] = 'd0;
        layer2_2[15:8] = 'd0;
        layer2_2[23:16] = 'd0;
        layer2_2[31:24] = 'd0;
        layer2_2[39:32] = 'd0;
        layer3_2[7:0] = 'd0;
        layer3_2[15:8] = 'd0;
        layer3_2[23:16] = 'd0;
        layer3_2[31:24] = 'd0;
        layer3_2[39:32] = 'd0;
        layer4_2[7:0] = 'd0;
        layer4_2[15:8] = 'd0;
        layer4_2[23:16] = 'd0;
        layer4_2[31:24] = 'd0;
        layer4_2[39:32] = 'd0;
        layer0_3[7:0] = 'd0;
        layer0_3[15:8] = 'd0;
        layer0_3[23:16] = 'd0;
        layer0_3[31:24] = 'd0;
        layer0_3[39:32] = 'd0;
        layer1_3[7:0] = 'd0;
        layer1_3[15:8] = 'd0;
        layer1_3[23:16] = 'd0;
        layer1_3[31:24] = 'd0;
        layer1_3[39:32] = 'd0;
        layer2_3[7:0] = 'd0;
        layer2_3[15:8] = 'd0;
        layer2_3[23:16] = 'd0;
        layer2_3[31:24] = 'd0;
        layer2_3[39:32] = 'd0;
        layer3_3[7:0] = 'd0;
        layer3_3[15:8] = 'd0;
        layer3_3[23:16] = 'd0;
        layer3_3[31:24] = 'd0;
        layer3_3[39:32] = 'd0;
        layer4_3[7:0] = 'd0;
        layer4_3[15:8] = 'd0;
        layer4_3[23:16] = 'd0;
        layer4_3[31:24] = 'd0;
        layer4_3[39:32] = 'd0;
        layer0_4[7:0] = 'd0;
        layer0_4[15:8] = 'd0;
        layer0_4[23:16] = 'd0;
        layer0_4[31:24] = 'd0;
        layer0_4[39:32] = 'd0;
        layer1_4[7:0] = 'd0;
        layer1_4[15:8] = 'd0;
        layer1_4[23:16] = 'd0;
        layer1_4[31:24] = 'd0;
        layer1_4[39:32] = 'd0;
        layer2_4[7:0] = 'd0;
        layer2_4[15:8] = 'd0;
        layer2_4[23:16] = 'd0;
        layer2_4[31:24] = 'd0;
        layer2_4[39:32] = 'd0;
        layer3_4[7:0] = 'd0;
        layer3_4[15:8] = 'd0;
        layer3_4[23:16] = 'd0;
        layer3_4[31:24] = 'd0;
        layer3_4[39:32] = 'd0;
        layer4_4[7:0] = 'd0;
        layer4_4[15:8] = 'd0;
        layer4_4[23:16] = 'd0;
        layer4_4[31:24] = 'd0;
        layer4_4[39:32] = 'd0;
        layer0_5[7:0] = 'd0;
        layer0_5[15:8] = 'd0;
        layer0_5[23:16] = 'd0;
        layer0_5[31:24] = 'd0;
        layer0_5[39:32] = 'd0;
        layer1_5[7:0] = 'd0;
        layer1_5[15:8] = 'd0;
        layer1_5[23:16] = 'd0;
        layer1_5[31:24] = 'd0;
        layer1_5[39:32] = 'd0;
        layer2_5[7:0] = 'd0;
        layer2_5[15:8] = 'd0;
        layer2_5[23:16] = 'd0;
        layer2_5[31:24] = 'd0;
        layer2_5[39:32] = 'd0;
        layer3_5[7:0] = 'd0;
        layer3_5[15:8] = 'd0;
        layer3_5[23:16] = 'd0;
        layer3_5[31:24] = 'd0;
        layer3_5[39:32] = 'd0;
        layer4_5[7:0] = 'd0;
        layer4_5[15:8] = 'd0;
        layer4_5[23:16] = 'd0;
        layer4_5[31:24] = 'd0;
        layer4_5[39:32] = 'd0;
        layer0_6[7:0] = 'd0;
        layer0_6[15:8] = 'd0;
        layer0_6[23:16] = 'd0;
        layer0_6[31:24] = 'd0;
        layer0_6[39:32] = 'd0;
        layer1_6[7:0] = 'd0;
        layer1_6[15:8] = 'd0;
        layer1_6[23:16] = 'd0;
        layer1_6[31:24] = 'd0;
        layer1_6[39:32] = 'd0;
        layer2_6[7:0] = 'd0;
        layer2_6[15:8] = 'd0;
        layer2_6[23:16] = 'd0;
        layer2_6[31:24] = 'd0;
        layer2_6[39:32] = 'd0;
        layer3_6[7:0] = 'd0;
        layer3_6[15:8] = 'd0;
        layer3_6[23:16] = 'd0;
        layer3_6[31:24] = 'd0;
        layer3_6[39:32] = 'd0;
        layer4_6[7:0] = 'd0;
        layer4_6[15:8] = 'd0;
        layer4_6[23:16] = 'd0;
        layer4_6[31:24] = 'd0;
        layer4_6[39:32] = 'd0;
        layer0_7[7:0] = 'd0;
        layer0_7[15:8] = 'd0;
        layer0_7[23:16] = 'd0;
        layer0_7[31:24] = 'd0;
        layer0_7[39:32] = 'd0;
        layer1_7[7:0] = 'd0;
        layer1_7[15:8] = 'd0;
        layer1_7[23:16] = 'd0;
        layer1_7[31:24] = 'd0;
        layer1_7[39:32] = 'd0;
        layer2_7[7:0] = 'd0;
        layer2_7[15:8] = 'd0;
        layer2_7[23:16] = 'd0;
        layer2_7[31:24] = 'd0;
        layer2_7[39:32] = 'd0;
        layer3_7[7:0] = 'd0;
        layer3_7[15:8] = 'd0;
        layer3_7[23:16] = 'd0;
        layer3_7[31:24] = 'd0;
        layer3_7[39:32] = 'd0;
        layer4_7[7:0] = 'd0;
        layer4_7[15:8] = 'd0;
        layer4_7[23:16] = 'd0;
        layer4_7[31:24] = 'd0;
        layer4_7[39:32] = 'd0;
        layer0_8[7:0] = 'd0;
        layer0_8[15:8] = 'd0;
        layer0_8[23:16] = 'd0;
        layer0_8[31:24] = 'd0;
        layer0_8[39:32] = 'd0;
        layer1_8[7:0] = 'd0;
        layer1_8[15:8] = 'd0;
        layer1_8[23:16] = 'd0;
        layer1_8[31:24] = 'd0;
        layer1_8[39:32] = 'd0;
        layer2_8[7:0] = 'd0;
        layer2_8[15:8] = 'd0;
        layer2_8[23:16] = 'd0;
        layer2_8[31:24] = 'd0;
        layer2_8[39:32] = 'd0;
        layer3_8[7:0] = 'd0;
        layer3_8[15:8] = 'd0;
        layer3_8[23:16] = 'd0;
        layer3_8[31:24] = 'd0;
        layer3_8[39:32] = 'd0;
        layer4_8[7:0] = 'd0;
        layer4_8[15:8] = 'd0;
        layer4_8[23:16] = 'd0;
        layer4_8[31:24] = 'd0;
        layer4_8[39:32] = 'd0;
        layer0_9[7:0] = 'd0;
        layer0_9[15:8] = 'd0;
        layer0_9[23:16] = 'd0;
        layer0_9[31:24] = 'd0;
        layer0_9[39:32] = 'd0;
        layer1_9[7:0] = 'd0;
        layer1_9[15:8] = 'd0;
        layer1_9[23:16] = 'd0;
        layer1_9[31:24] = 'd0;
        layer1_9[39:32] = 'd0;
        layer2_9[7:0] = 'd0;
        layer2_9[15:8] = 'd0;
        layer2_9[23:16] = 'd0;
        layer2_9[31:24] = 'd0;
        layer2_9[39:32] = 'd0;
        layer3_9[7:0] = 'd0;
        layer3_9[15:8] = 'd0;
        layer3_9[23:16] = 'd0;
        layer3_9[31:24] = 'd0;
        layer3_9[39:32] = 'd0;
        layer4_9[7:0] = 'd0;
        layer4_9[15:8] = 'd0;
        layer4_9[23:16] = 'd0;
        layer4_9[31:24] = 'd0;
        layer4_9[39:32] = 'd0;
        layer0_10[7:0] = 'd0;
        layer0_10[15:8] = 'd0;
        layer0_10[23:16] = 'd0;
        layer0_10[31:24] = 'd0;
        layer0_10[39:32] = 'd0;
        layer1_10[7:0] = 'd0;
        layer1_10[15:8] = 'd0;
        layer1_10[23:16] = 'd0;
        layer1_10[31:24] = 'd0;
        layer1_10[39:32] = 'd0;
        layer2_10[7:0] = 'd0;
        layer2_10[15:8] = 'd0;
        layer2_10[23:16] = 'd0;
        layer2_10[31:24] = 'd0;
        layer2_10[39:32] = 'd0;
        layer3_10[7:0] = 'd0;
        layer3_10[15:8] = 'd0;
        layer3_10[23:16] = 'd0;
        layer3_10[31:24] = 'd0;
        layer3_10[39:32] = 'd0;
        layer4_10[7:0] = 'd0;
        layer4_10[15:8] = 'd0;
        layer4_10[23:16] = 'd0;
        layer4_10[31:24] = 'd0;
        layer4_10[39:32] = 'd0;
        layer0_11[7:0] = 'd0;
        layer0_11[15:8] = 'd0;
        layer0_11[23:16] = 'd0;
        layer0_11[31:24] = 'd0;
        layer0_11[39:32] = 'd0;
        layer1_11[7:0] = 'd0;
        layer1_11[15:8] = 'd0;
        layer1_11[23:16] = 'd0;
        layer1_11[31:24] = 'd0;
        layer1_11[39:32] = 'd0;
        layer2_11[7:0] = 'd0;
        layer2_11[15:8] = 'd0;
        layer2_11[23:16] = 'd0;
        layer2_11[31:24] = 'd0;
        layer2_11[39:32] = 'd0;
        layer3_11[7:0] = 'd0;
        layer3_11[15:8] = 'd0;
        layer3_11[23:16] = 'd0;
        layer3_11[31:24] = 'd0;
        layer3_11[39:32] = 'd0;
        layer4_11[7:0] = 'd0;
        layer4_11[15:8] = 'd0;
        layer4_11[23:16] = 'd0;
        layer4_11[31:24] = 'd0;
        layer4_11[39:32] = 'd0;
        layer0_12[7:0] = 'd0;
        layer0_12[15:8] = 'd0;
        layer0_12[23:16] = 'd0;
        layer0_12[31:24] = 'd0;
        layer0_12[39:32] = 'd0;
        layer1_12[7:0] = 'd0;
        layer1_12[15:8] = 'd0;
        layer1_12[23:16] = 'd0;
        layer1_12[31:24] = 'd0;
        layer1_12[39:32] = 'd0;
        layer2_12[7:0] = 'd0;
        layer2_12[15:8] = 'd0;
        layer2_12[23:16] = 'd0;
        layer2_12[31:24] = 'd0;
        layer2_12[39:32] = 'd0;
        layer3_12[7:0] = 'd0;
        layer3_12[15:8] = 'd0;
        layer3_12[23:16] = 'd0;
        layer3_12[31:24] = 'd0;
        layer3_12[39:32] = 'd0;
        layer4_12[7:0] = 'd0;
        layer4_12[15:8] = 'd0;
        layer4_12[23:16] = 'd0;
        layer4_12[31:24] = 'd0;
        layer4_12[39:32] = 'd0;
        layer0_13[7:0] = 'd0;
        layer0_13[15:8] = 'd0;
        layer0_13[23:16] = 'd0;
        layer0_13[31:24] = 'd0;
        layer0_13[39:32] = 'd0;
        layer1_13[7:0] = 'd0;
        layer1_13[15:8] = 'd0;
        layer1_13[23:16] = 'd0;
        layer1_13[31:24] = 'd0;
        layer1_13[39:32] = 'd0;
        layer2_13[7:0] = 'd0;
        layer2_13[15:8] = 'd0;
        layer2_13[23:16] = 'd0;
        layer2_13[31:24] = 'd0;
        layer2_13[39:32] = 'd0;
        layer3_13[7:0] = 'd0;
        layer3_13[15:8] = 'd0;
        layer3_13[23:16] = 'd0;
        layer3_13[31:24] = 'd0;
        layer3_13[39:32] = 'd0;
        layer4_13[7:0] = 'd0;
        layer4_13[15:8] = 'd0;
        layer4_13[23:16] = 'd0;
        layer4_13[31:24] = 'd0;
        layer4_13[39:32] = 'd0;
        layer0_14[7:0] = 'd0;
        layer0_14[15:8] = 'd0;
        layer0_14[23:16] = 'd0;
        layer0_14[31:24] = 'd0;
        layer0_14[39:32] = 'd0;
        layer1_14[7:0] = 'd0;
        layer1_14[15:8] = 'd0;
        layer1_14[23:16] = 'd0;
        layer1_14[31:24] = 'd0;
        layer1_14[39:32] = 'd0;
        layer2_14[7:0] = 'd0;
        layer2_14[15:8] = 'd0;
        layer2_14[23:16] = 'd0;
        layer2_14[31:24] = 'd0;
        layer2_14[39:32] = 'd0;
        layer3_14[7:0] = 'd0;
        layer3_14[15:8] = 'd0;
        layer3_14[23:16] = 'd0;
        layer3_14[31:24] = 'd0;
        layer3_14[39:32] = 'd0;
        layer4_14[7:0] = 'd0;
        layer4_14[15:8] = 'd0;
        layer4_14[23:16] = 'd0;
        layer4_14[31:24] = 'd0;
        layer4_14[39:32] = 'd0;
        layer0_15[7:0] = 'd0;
        layer0_15[15:8] = 'd0;
        layer0_15[23:16] = 'd0;
        layer0_15[31:24] = 'd0;
        layer0_15[39:32] = 'd0;
        layer1_15[7:0] = 'd0;
        layer1_15[15:8] = 'd0;
        layer1_15[23:16] = 'd0;
        layer1_15[31:24] = 'd0;
        layer1_15[39:32] = 'd0;
        layer2_15[7:0] = 'd0;
        layer2_15[15:8] = 'd0;
        layer2_15[23:16] = 'd0;
        layer2_15[31:24] = 'd0;
        layer2_15[39:32] = 'd0;
        layer3_15[7:0] = 'd0;
        layer3_15[15:8] = 'd0;
        layer3_15[23:16] = 'd0;
        layer3_15[31:24] = 'd0;
        layer3_15[39:32] = 'd0;
        layer4_15[7:0] = 'd0;
        layer4_15[15:8] = 'd0;
        layer4_15[23:16] = 'd0;
        layer4_15[31:24] = 'd0;
        layer4_15[39:32] = 'd0;
    end
  endcase
end

reg    [39:0]    layer0_reg_0;
reg    [39:0]    layer0_reg_1;
reg    [39:0]    layer0_reg_2;
reg    [39:0]    layer0_reg_3;
reg    [39:0]    layer0_reg_4;
reg    [39:0]    layer0_reg_5;
reg    [39:0]    layer0_reg_6;
reg    [39:0]    layer0_reg_7;
reg    [39:0]    layer0_reg_8;
reg    [39:0]    layer0_reg_9;
reg    [39:0]    layer0_reg_10;
reg    [39:0]    layer0_reg_11;
reg    [39:0]    layer0_reg_12;
reg    [39:0]    layer0_reg_13;
reg    [39:0]    layer0_reg_14;
reg    [39:0]    layer0_reg_15;
reg    [39:0]    layer1_reg_0;
reg    [39:0]    layer1_reg_1;
reg    [39:0]    layer1_reg_2;
reg    [39:0]    layer1_reg_3;
reg    [39:0]    layer1_reg_4;
reg    [39:0]    layer1_reg_5;
reg    [39:0]    layer1_reg_6;
reg    [39:0]    layer1_reg_7;
reg    [39:0]    layer1_reg_8;
reg    [39:0]    layer1_reg_9;
reg    [39:0]    layer1_reg_10;
reg    [39:0]    layer1_reg_11;
reg    [39:0]    layer1_reg_12;
reg    [39:0]    layer1_reg_13;
reg    [39:0]    layer1_reg_14;
reg    [39:0]    layer1_reg_15;
reg    [39:0]    layer2_reg_0;
reg    [39:0]    layer2_reg_1;
reg    [39:0]    layer2_reg_2;
reg    [39:0]    layer2_reg_3;
reg    [39:0]    layer2_reg_4;
reg    [39:0]    layer2_reg_5;
reg    [39:0]    layer2_reg_6;
reg    [39:0]    layer2_reg_7;
reg    [39:0]    layer2_reg_8;
reg    [39:0]    layer2_reg_9;
reg    [39:0]    layer2_reg_10;
reg    [39:0]    layer2_reg_11;
reg    [39:0]    layer2_reg_12;
reg    [39:0]    layer2_reg_13;
reg    [39:0]    layer2_reg_14;
reg    [39:0]    layer2_reg_15;
reg    [39:0]    layer3_reg_0;
reg    [39:0]    layer3_reg_1;
reg    [39:0]    layer3_reg_2;
reg    [39:0]    layer3_reg_3;
reg    [39:0]    layer3_reg_4;
reg    [39:0]    layer3_reg_5;
reg    [39:0]    layer3_reg_6;
reg    [39:0]    layer3_reg_7;
reg    [39:0]    layer3_reg_8;
reg    [39:0]    layer3_reg_9;
reg    [39:0]    layer3_reg_10;
reg    [39:0]    layer3_reg_11;
reg    [39:0]    layer3_reg_12;
reg    [39:0]    layer3_reg_13;
reg    [39:0]    layer3_reg_14;
reg    [39:0]    layer3_reg_15;
reg    [39:0]    layer4_reg_0;
reg    [39:0]    layer4_reg_1;
reg    [39:0]    layer4_reg_2;
reg    [39:0]    layer4_reg_3;
reg    [39:0]    layer4_reg_4;
reg    [39:0]    layer4_reg_5;
reg    [39:0]    layer4_reg_6;
reg    [39:0]    layer4_reg_7;
reg    [39:0]    layer4_reg_8;
reg    [39:0]    layer4_reg_9;
reg    [39:0]    layer4_reg_10;
reg    [39:0]    layer4_reg_11;
reg    [39:0]    layer4_reg_12;
reg    [39:0]    layer4_reg_13;
reg    [39:0]    layer4_reg_14;
reg    [39:0]    layer4_reg_15;
always@(posedge clk) begin
  if(!rst_n) begin
    layer0_reg_0 <= 'd0;
    layer0_reg_1 <= 'd0;
    layer0_reg_2 <= 'd0;
    layer0_reg_3 <= 'd0;
    layer0_reg_4 <= 'd0;
    layer0_reg_5 <= 'd0;
    layer0_reg_6 <= 'd0;
    layer0_reg_7 <= 'd0;
    layer0_reg_8 <= 'd0;
    layer0_reg_9 <= 'd0;
    layer0_reg_10 <= 'd0;
    layer0_reg_11 <= 'd0;
    layer0_reg_12 <= 'd0;
    layer0_reg_13 <= 'd0;
    layer0_reg_14 <= 'd0;
    layer0_reg_15 <= 'd0;
    layer1_reg_0 <= 'd0;
    layer1_reg_1 <= 'd0;
    layer1_reg_2 <= 'd0;
    layer1_reg_3 <= 'd0;
    layer1_reg_4 <= 'd0;
    layer1_reg_5 <= 'd0;
    layer1_reg_6 <= 'd0;
    layer1_reg_7 <= 'd0;
    layer1_reg_8 <= 'd0;
    layer1_reg_9 <= 'd0;
    layer1_reg_10 <= 'd0;
    layer1_reg_11 <= 'd0;
    layer1_reg_12 <= 'd0;
    layer1_reg_13 <= 'd0;
    layer1_reg_14 <= 'd0;
    layer1_reg_15 <= 'd0;
    layer2_reg_0 <= 'd0;
    layer2_reg_1 <= 'd0;
    layer2_reg_2 <= 'd0;
    layer2_reg_3 <= 'd0;
    layer2_reg_4 <= 'd0;
    layer2_reg_5 <= 'd0;
    layer2_reg_6 <= 'd0;
    layer2_reg_7 <= 'd0;
    layer2_reg_8 <= 'd0;
    layer2_reg_9 <= 'd0;
    layer2_reg_10 <= 'd0;
    layer2_reg_11 <= 'd0;
    layer2_reg_12 <= 'd0;
    layer2_reg_13 <= 'd0;
    layer2_reg_14 <= 'd0;
    layer2_reg_15 <= 'd0;
    layer3_reg_0 <= 'd0;
    layer3_reg_1 <= 'd0;
    layer3_reg_2 <= 'd0;
    layer3_reg_3 <= 'd0;
    layer3_reg_4 <= 'd0;
    layer3_reg_5 <= 'd0;
    layer3_reg_6 <= 'd0;
    layer3_reg_7 <= 'd0;
    layer3_reg_8 <= 'd0;
    layer3_reg_9 <= 'd0;
    layer3_reg_10 <= 'd0;
    layer3_reg_11 <= 'd0;
    layer3_reg_12 <= 'd0;
    layer3_reg_13 <= 'd0;
    layer3_reg_14 <= 'd0;
    layer3_reg_15 <= 'd0;
    layer4_reg_0 <= 'd0;
    layer4_reg_1 <= 'd0;
    layer4_reg_2 <= 'd0;
    layer4_reg_3 <= 'd0;
    layer4_reg_4 <= 'd0;
    layer4_reg_5 <= 'd0;
    layer4_reg_6 <= 'd0;
    layer4_reg_7 <= 'd0;
    layer4_reg_8 <= 'd0;
    layer4_reg_9 <= 'd0;
    layer4_reg_10 <= 'd0;
    layer4_reg_11 <= 'd0;
    layer4_reg_12 <= 'd0;
    layer4_reg_13 <= 'd0;
    layer4_reg_14 <= 'd0;
    layer4_reg_15 <= 'd0;
  end
  else if(current_state==ST_MUX) begin
    layer0_reg_0 <= layer0_0;
    layer0_reg_1 <= layer0_1;
    layer0_reg_2 <= layer0_2;
    layer0_reg_3 <= layer0_3;
    layer0_reg_4 <= layer0_4;
    layer0_reg_5 <= layer0_5;
    layer0_reg_6 <= layer0_6;
    layer0_reg_7 <= layer0_7;
    layer0_reg_8 <= layer0_8;
    layer0_reg_9 <= layer0_9;
    layer0_reg_10 <= layer0_10;
    layer0_reg_11 <= layer0_11;
    layer0_reg_12 <= layer0_12;
    layer0_reg_13 <= layer0_13;
    layer0_reg_14 <= layer0_14;
    layer0_reg_15 <= layer0_15;
    layer1_reg_0 <= layer1_0;
    layer1_reg_1 <= layer1_1;
    layer1_reg_2 <= layer1_2;
    layer1_reg_3 <= layer1_3;
    layer1_reg_4 <= layer1_4;
    layer1_reg_5 <= layer1_5;
    layer1_reg_6 <= layer1_6;
    layer1_reg_7 <= layer1_7;
    layer1_reg_8 <= layer1_8;
    layer1_reg_9 <= layer1_9;
    layer1_reg_10 <= layer1_10;
    layer1_reg_11 <= layer1_11;
    layer1_reg_12 <= layer1_12;
    layer1_reg_13 <= layer1_13;
    layer1_reg_14 <= layer1_14;
    layer1_reg_15 <= layer1_15;
    layer2_reg_0 <= layer2_0;
    layer2_reg_1 <= layer2_1;
    layer2_reg_2 <= layer2_2;
    layer2_reg_3 <= layer2_3;
    layer2_reg_4 <= layer2_4;
    layer2_reg_5 <= layer2_5;
    layer2_reg_6 <= layer2_6;
    layer2_reg_7 <= layer2_7;
    layer2_reg_8 <= layer2_8;
    layer2_reg_9 <= layer2_9;
    layer2_reg_10 <= layer2_10;
    layer2_reg_11 <= layer2_11;
    layer2_reg_12 <= layer2_12;
    layer2_reg_13 <= layer2_13;
    layer2_reg_14 <= layer2_14;
    layer2_reg_15 <= layer2_15;
    layer3_reg_0 <= layer3_0;
    layer3_reg_1 <= layer3_1;
    layer3_reg_2 <= layer3_2;
    layer3_reg_3 <= layer3_3;
    layer3_reg_4 <= layer3_4;
    layer3_reg_5 <= layer3_5;
    layer3_reg_6 <= layer3_6;
    layer3_reg_7 <= layer3_7;
    layer3_reg_8 <= layer3_8;
    layer3_reg_9 <= layer3_9;
    layer3_reg_10 <= layer3_10;
    layer3_reg_11 <= layer3_11;
    layer3_reg_12 <= layer3_12;
    layer3_reg_13 <= layer3_13;
    layer3_reg_14 <= layer3_14;
    layer3_reg_15 <= layer3_15;
    layer4_reg_0 <= layer4_0;
    layer4_reg_1 <= layer4_1;
    layer4_reg_2 <= layer4_2;
    layer4_reg_3 <= layer4_3;
    layer4_reg_4 <= layer4_4;
    layer4_reg_5 <= layer4_5;
    layer4_reg_6 <= layer4_6;
    layer4_reg_7 <= layer4_7;
    layer4_reg_8 <= layer4_8;
    layer4_reg_9 <= layer4_9;
    layer4_reg_10 <= layer4_10;
    layer4_reg_11 <= layer4_11;
    layer4_reg_12 <= layer4_12;
    layer4_reg_13 <= layer4_13;
    layer4_reg_14 <= layer4_14;
    layer4_reg_15 <= layer4_15;
  end
end
reg  [15:0]  kernel_img_mul_0[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_0[0] <= 'd0;
    kernel_img_mul_0[1] <= 'd0;
    kernel_img_mul_0[2] <= 'd0;
    kernel_img_mul_0[3] <= 'd0;
    kernel_img_mul_0[4] <= 'd0;
    kernel_img_mul_0[5] <= 'd0;
    kernel_img_mul_0[6] <= 'd0;
    kernel_img_mul_0[7] <= 'd0;
    kernel_img_mul_0[8] <= 'd0;
    kernel_img_mul_0[9] <= 'd0;
    kernel_img_mul_0[10] <= 'd0;
    kernel_img_mul_0[11] <= 'd0;
    kernel_img_mul_0[12] <= 'd0;
    kernel_img_mul_0[13] <= 'd0;
    kernel_img_mul_0[14] <= 'd0;
    kernel_img_mul_0[15] <= 'd0;
    kernel_img_mul_0[16] <= 'd0;
    kernel_img_mul_0[17] <= 'd0;
    kernel_img_mul_0[18] <= 'd0;
    kernel_img_mul_0[19] <= 'd0;
    kernel_img_mul_0[20] <= 'd0;
    kernel_img_mul_0[21] <= 'd0;
    kernel_img_mul_0[22] <= 'd0;
    kernel_img_mul_0[23] <= 'd0;
    kernel_img_mul_0[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_0[0] <= { {8{1'b0}},layer0_reg_0[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_0[1] <= { {8{1'b0}},layer0_reg_0[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_0[2] <= { {8{1'b0}},layer0_reg_0[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_0[3] <= { {8{1'b0}},layer0_reg_0[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_0[4] <= { {8{1'b0}},layer0_reg_0[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_0[5] <= { {8{1'b0}},layer1_reg_0[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_0[6] <= { {8{1'b0}},layer1_reg_0[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_0[7] <= { {8{1'b0}},layer1_reg_0[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_0[8] <= { {8{1'b0}},layer1_reg_0[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_0[9] <= { {8{1'b0}},layer1_reg_0[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_0[10] <= { {8{1'b0}},layer2_reg_0[7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_0[11] <= { {8{1'b0}},layer2_reg_0[15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_0[12] <= { {8{1'b0}},layer2_reg_0[23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_0[13] <= { {8{1'b0}},layer2_reg_0[31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_0[14] <= { {8{1'b0}},layer2_reg_0[39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_0[15] <= { {8{1'b0}},layer3_reg_0[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_0[16] <= { {8{1'b0}},layer3_reg_0[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_0[17] <= { {8{1'b0}},layer3_reg_0[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_0[18] <= { {8{1'b0}},layer3_reg_0[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_0[19] <= { {8{1'b0}},layer3_reg_0[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_0[20] <= { {8{1'b0}},layer4_reg_0[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_0[21] <= { {8{1'b0}},layer4_reg_0[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_0[22] <= { {8{1'b0}},layer4_reg_0[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_0[23] <= { {8{1'b0}},layer4_reg_0[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_0[24] <= { {8{1'b0}},layer4_reg_0[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_0;
reg  [15:0]  kernel_img_sum_2_0;
reg  [15:0]  kernel_img_sum_3_0;
reg  [15:0]  kernel_img_sum_4_0;
reg  [15:0]  kernel_img_sum_5_0;
reg  [15:0]  kernel_img_sum_6_0;
reg  [15:0]  kernel_img_sum_7_0;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_0 <= kernel_img_mul_0[0] + kernel_img_mul_0[1] + kernel_img_mul_0[2] + kernel_img_mul_0[3] + kernel_img_mul_0[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_0 <= kernel_img_mul_0[5] + kernel_img_mul_0[6] + kernel_img_mul_0[7] + kernel_img_mul_0[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_0 <= kernel_img_mul_0[9] + kernel_img_mul_0[10] + kernel_img_mul_0[11] + kernel_img_mul_0[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_0 <= kernel_img_mul_0[13] + kernel_img_mul_0[14] + kernel_img_mul_0[15] + kernel_img_mul_0[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_0 <= kernel_img_mul_0[17] + kernel_img_mul_0[18] + kernel_img_mul_0[19] + kernel_img_mul_0[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_0 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_0 <= kernel_img_mul_0[21] + kernel_img_mul_0[22] + kernel_img_mul_0[23] + kernel_img_mul_0[24];
  end
end
always@(*) begin
  kernel_img_sum_7_0 = kernel_img_sum_1_0 + kernel_img_sum_2_0 + kernel_img_sum_3_0 + kernel_img_sum_4_0 + kernel_img_sum_5_0 + kernel_img_sum_6_0;
end
reg  [15:0]  kernel_img_mul_1[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_1[0] <= 'd0;
    kernel_img_mul_1[1] <= 'd0;
    kernel_img_mul_1[2] <= 'd0;
    kernel_img_mul_1[3] <= 'd0;
    kernel_img_mul_1[4] <= 'd0;
    kernel_img_mul_1[5] <= 'd0;
    kernel_img_mul_1[6] <= 'd0;
    kernel_img_mul_1[7] <= 'd0;
    kernel_img_mul_1[8] <= 'd0;
    kernel_img_mul_1[9] <= 'd0;
    kernel_img_mul_1[10] <= 'd0;
    kernel_img_mul_1[11] <= 'd0;
    kernel_img_mul_1[12] <= 'd0;
    kernel_img_mul_1[13] <= 'd0;
    kernel_img_mul_1[14] <= 'd0;
    kernel_img_mul_1[15] <= 'd0;
    kernel_img_mul_1[16] <= 'd0;
    kernel_img_mul_1[17] <= 'd0;
    kernel_img_mul_1[18] <= 'd0;
    kernel_img_mul_1[19] <= 'd0;
    kernel_img_mul_1[20] <= 'd0;
    kernel_img_mul_1[21] <= 'd0;
    kernel_img_mul_1[22] <= 'd0;
    kernel_img_mul_1[23] <= 'd0;
    kernel_img_mul_1[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_1[0] <= { {8{1'b0}},layer0_reg_1[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_1[1] <= { {8{1'b0}},layer0_reg_1[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_1[2] <= { {8{1'b0}},layer0_reg_1[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_1[3] <= { {8{1'b0}},layer0_reg_1[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_1[4] <= { {8{1'b0}},layer0_reg_1[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_1[5] <= { {8{1'b0}},layer1_reg_1[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_1[6] <= { {8{1'b0}},layer1_reg_1[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_1[7] <= { {8{1'b0}},layer1_reg_1[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_1[8] <= { {8{1'b0}},layer1_reg_1[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_1[9] <= { {8{1'b0}},layer1_reg_1[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_1[10] <= { {8{1'b0}},layer2_reg_1[7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_1[11] <= { {8{1'b0}},layer2_reg_1[15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_1[12] <= { {8{1'b0}},layer2_reg_1[23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_1[13] <= { {8{1'b0}},layer2_reg_1[31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_1[14] <= { {8{1'b0}},layer2_reg_1[39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_1[15] <= { {8{1'b0}},layer3_reg_1[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_1[16] <= { {8{1'b0}},layer3_reg_1[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_1[17] <= { {8{1'b0}},layer3_reg_1[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_1[18] <= { {8{1'b0}},layer3_reg_1[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_1[19] <= { {8{1'b0}},layer3_reg_1[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_1[20] <= { {8{1'b0}},layer4_reg_1[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_1[21] <= { {8{1'b0}},layer4_reg_1[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_1[22] <= { {8{1'b0}},layer4_reg_1[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_1[23] <= { {8{1'b0}},layer4_reg_1[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_1[24] <= { {8{1'b0}},layer4_reg_1[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_1;
reg  [15:0]  kernel_img_sum_2_1;
reg  [15:0]  kernel_img_sum_3_1;
reg  [15:0]  kernel_img_sum_4_1;
reg  [15:0]  kernel_img_sum_5_1;
reg  [15:0]  kernel_img_sum_6_1;
reg  [15:0]  kernel_img_sum_7_1;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_1 <= kernel_img_mul_1[0] + kernel_img_mul_1[1] + kernel_img_mul_1[2] + kernel_img_mul_1[3] + kernel_img_mul_1[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_1 <= kernel_img_mul_1[5] + kernel_img_mul_1[6] + kernel_img_mul_1[7] + kernel_img_mul_1[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_1 <= kernel_img_mul_1[9] + kernel_img_mul_1[10] + kernel_img_mul_1[11] + kernel_img_mul_1[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_1 <= kernel_img_mul_1[13] + kernel_img_mul_1[14] + kernel_img_mul_1[15] + kernel_img_mul_1[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_1 <= kernel_img_mul_1[17] + kernel_img_mul_1[18] + kernel_img_mul_1[19] + kernel_img_mul_1[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_1 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_1 <= kernel_img_mul_1[21] + kernel_img_mul_1[22] + kernel_img_mul_1[23] + kernel_img_mul_1[24];
  end
end
always@(*) begin
  kernel_img_sum_7_1 = kernel_img_sum_1_1 + kernel_img_sum_2_1 + kernel_img_sum_3_1 + kernel_img_sum_4_1 + kernel_img_sum_5_1 + kernel_img_sum_6_1;
end
reg  [15:0]  kernel_img_mul_2[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_2[0] <= 'd0;
    kernel_img_mul_2[1] <= 'd0;
    kernel_img_mul_2[2] <= 'd0;
    kernel_img_mul_2[3] <= 'd0;
    kernel_img_mul_2[4] <= 'd0;
    kernel_img_mul_2[5] <= 'd0;
    kernel_img_mul_2[6] <= 'd0;
    kernel_img_mul_2[7] <= 'd0;
    kernel_img_mul_2[8] <= 'd0;
    kernel_img_mul_2[9] <= 'd0;
    kernel_img_mul_2[10] <= 'd0;
    kernel_img_mul_2[11] <= 'd0;
    kernel_img_mul_2[12] <= 'd0;
    kernel_img_mul_2[13] <= 'd0;
    kernel_img_mul_2[14] <= 'd0;
    kernel_img_mul_2[15] <= 'd0;
    kernel_img_mul_2[16] <= 'd0;
    kernel_img_mul_2[17] <= 'd0;
    kernel_img_mul_2[18] <= 'd0;
    kernel_img_mul_2[19] <= 'd0;
    kernel_img_mul_2[20] <= 'd0;
    kernel_img_mul_2[21] <= 'd0;
    kernel_img_mul_2[22] <= 'd0;
    kernel_img_mul_2[23] <= 'd0;
    kernel_img_mul_2[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_2[0] <= { {8{1'b0}},layer0_reg_2[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_2[1] <= { {8{1'b0}},layer0_reg_2[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_2[2] <= { {8{1'b0}},layer0_reg_2[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_2[3] <= { {8{1'b0}},layer0_reg_2[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_2[4] <= { {8{1'b0}},layer0_reg_2[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_2[5] <= { {8{1'b0}},layer1_reg_2[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_2[6] <= { {8{1'b0}},layer1_reg_2[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_2[7] <= { {8{1'b0}},layer1_reg_2[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_2[8] <= { {8{1'b0}},layer1_reg_2[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_2[9] <= { {8{1'b0}},layer1_reg_2[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_2[10] <= { {8{1'b0}},layer2_reg_2[7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_2[11] <= { {8{1'b0}},layer2_reg_2[15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_2[12] <= { {8{1'b0}},layer2_reg_2[23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_2[13] <= { {8{1'b0}},layer2_reg_2[31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_2[14] <= { {8{1'b0}},layer2_reg_2[39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_2[15] <= { {8{1'b0}},layer3_reg_2[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_2[16] <= { {8{1'b0}},layer3_reg_2[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_2[17] <= { {8{1'b0}},layer3_reg_2[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_2[18] <= { {8{1'b0}},layer3_reg_2[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_2[19] <= { {8{1'b0}},layer3_reg_2[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_2[20] <= { {8{1'b0}},layer4_reg_2[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_2[21] <= { {8{1'b0}},layer4_reg_2[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_2[22] <= { {8{1'b0}},layer4_reg_2[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_2[23] <= { {8{1'b0}},layer4_reg_2[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_2[24] <= { {8{1'b0}},layer4_reg_2[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_2;
reg  [15:0]  kernel_img_sum_2_2;
reg  [15:0]  kernel_img_sum_3_2;
reg  [15:0]  kernel_img_sum_4_2;
reg  [15:0]  kernel_img_sum_5_2;
reg  [15:0]  kernel_img_sum_6_2;
reg  [15:0]  kernel_img_sum_7_2;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_2 <= kernel_img_mul_2[0] + kernel_img_mul_2[1] + kernel_img_mul_2[2] + kernel_img_mul_2[3] + kernel_img_mul_2[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_2 <= kernel_img_mul_2[5] + kernel_img_mul_2[6] + kernel_img_mul_2[7] + kernel_img_mul_2[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_2 <= kernel_img_mul_2[9] + kernel_img_mul_2[10] + kernel_img_mul_2[11] + kernel_img_mul_2[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_2 <= kernel_img_mul_2[13] + kernel_img_mul_2[14] + kernel_img_mul_2[15] + kernel_img_mul_2[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_2 <= kernel_img_mul_2[17] + kernel_img_mul_2[18] + kernel_img_mul_2[19] + kernel_img_mul_2[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_2 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_2 <= kernel_img_mul_2[21] + kernel_img_mul_2[22] + kernel_img_mul_2[23] + kernel_img_mul_2[24];
  end
end
always@(*) begin
  kernel_img_sum_7_2 = kernel_img_sum_1_2 + kernel_img_sum_2_2 + kernel_img_sum_3_2 + kernel_img_sum_4_2 + kernel_img_sum_5_2 + kernel_img_sum_6_2;
end
reg  [15:0]  kernel_img_mul_3[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_3[0] <= 'd0;
    kernel_img_mul_3[1] <= 'd0;
    kernel_img_mul_3[2] <= 'd0;
    kernel_img_mul_3[3] <= 'd0;
    kernel_img_mul_3[4] <= 'd0;
    kernel_img_mul_3[5] <= 'd0;
    kernel_img_mul_3[6] <= 'd0;
    kernel_img_mul_3[7] <= 'd0;
    kernel_img_mul_3[8] <= 'd0;
    kernel_img_mul_3[9] <= 'd0;
    kernel_img_mul_3[10] <= 'd0;
    kernel_img_mul_3[11] <= 'd0;
    kernel_img_mul_3[12] <= 'd0;
    kernel_img_mul_3[13] <= 'd0;
    kernel_img_mul_3[14] <= 'd0;
    kernel_img_mul_3[15] <= 'd0;
    kernel_img_mul_3[16] <= 'd0;
    kernel_img_mul_3[17] <= 'd0;
    kernel_img_mul_3[18] <= 'd0;
    kernel_img_mul_3[19] <= 'd0;
    kernel_img_mul_3[20] <= 'd0;
    kernel_img_mul_3[21] <= 'd0;
    kernel_img_mul_3[22] <= 'd0;
    kernel_img_mul_3[23] <= 'd0;
    kernel_img_mul_3[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_3[0] <= { {8{1'b0}},layer0_reg_3[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_3[1] <= { {8{1'b0}},layer0_reg_3[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_3[2] <= { {8{1'b0}},layer0_reg_3[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_3[3] <= { {8{1'b0}},layer0_reg_3[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_3[4] <= { {8{1'b0}},layer0_reg_3[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_3[5] <= { {8{1'b0}},layer1_reg_3[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_3[6] <= { {8{1'b0}},layer1_reg_3[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_3[7] <= { {8{1'b0}},layer1_reg_3[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_3[8] <= { {8{1'b0}},layer1_reg_3[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_3[9] <= { {8{1'b0}},layer1_reg_3[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_3[10] <= { {8{1'b0}},layer2_reg_3[7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_3[11] <= { {8{1'b0}},layer2_reg_3[15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_3[12] <= { {8{1'b0}},layer2_reg_3[23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_3[13] <= { {8{1'b0}},layer2_reg_3[31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_3[14] <= { {8{1'b0}},layer2_reg_3[39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_3[15] <= { {8{1'b0}},layer3_reg_3[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_3[16] <= { {8{1'b0}},layer3_reg_3[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_3[17] <= { {8{1'b0}},layer3_reg_3[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_3[18] <= { {8{1'b0}},layer3_reg_3[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_3[19] <= { {8{1'b0}},layer3_reg_3[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_3[20] <= { {8{1'b0}},layer4_reg_3[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_3[21] <= { {8{1'b0}},layer4_reg_3[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_3[22] <= { {8{1'b0}},layer4_reg_3[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_3[23] <= { {8{1'b0}},layer4_reg_3[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_3[24] <= { {8{1'b0}},layer4_reg_3[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_3;
reg  [15:0]  kernel_img_sum_2_3;
reg  [15:0]  kernel_img_sum_3_3;
reg  [15:0]  kernel_img_sum_4_3;
reg  [15:0]  kernel_img_sum_5_3;
reg  [15:0]  kernel_img_sum_6_3;
reg  [15:0]  kernel_img_sum_7_3;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_3 <= kernel_img_mul_3[0] + kernel_img_mul_3[1] + kernel_img_mul_3[2] + kernel_img_mul_3[3] + kernel_img_mul_3[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_3 <= kernel_img_mul_3[5] + kernel_img_mul_3[6] + kernel_img_mul_3[7] + kernel_img_mul_3[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_3 <= kernel_img_mul_3[9] + kernel_img_mul_3[10] + kernel_img_mul_3[11] + kernel_img_mul_3[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_3 <= kernel_img_mul_3[13] + kernel_img_mul_3[14] + kernel_img_mul_3[15] + kernel_img_mul_3[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_3 <= kernel_img_mul_3[17] + kernel_img_mul_3[18] + kernel_img_mul_3[19] + kernel_img_mul_3[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_3 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_3 <= kernel_img_mul_3[21] + kernel_img_mul_3[22] + kernel_img_mul_3[23] + kernel_img_mul_3[24];
  end
end
always@(*) begin
  kernel_img_sum_7_3 = kernel_img_sum_1_3 + kernel_img_sum_2_3 + kernel_img_sum_3_3 + kernel_img_sum_4_3 + kernel_img_sum_5_3 + kernel_img_sum_6_3;
end
reg  [15:0]  kernel_img_mul_4[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_4[0] <= 'd0;
    kernel_img_mul_4[1] <= 'd0;
    kernel_img_mul_4[2] <= 'd0;
    kernel_img_mul_4[3] <= 'd0;
    kernel_img_mul_4[4] <= 'd0;
    kernel_img_mul_4[5] <= 'd0;
    kernel_img_mul_4[6] <= 'd0;
    kernel_img_mul_4[7] <= 'd0;
    kernel_img_mul_4[8] <= 'd0;
    kernel_img_mul_4[9] <= 'd0;
    kernel_img_mul_4[10] <= 'd0;
    kernel_img_mul_4[11] <= 'd0;
    kernel_img_mul_4[12] <= 'd0;
    kernel_img_mul_4[13] <= 'd0;
    kernel_img_mul_4[14] <= 'd0;
    kernel_img_mul_4[15] <= 'd0;
    kernel_img_mul_4[16] <= 'd0;
    kernel_img_mul_4[17] <= 'd0;
    kernel_img_mul_4[18] <= 'd0;
    kernel_img_mul_4[19] <= 'd0;
    kernel_img_mul_4[20] <= 'd0;
    kernel_img_mul_4[21] <= 'd0;
    kernel_img_mul_4[22] <= 'd0;
    kernel_img_mul_4[23] <= 'd0;
    kernel_img_mul_4[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_4[0] <= { {8{1'b0}},layer0_reg_4[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_4[1] <= { {8{1'b0}},layer0_reg_4[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_4[2] <= { {8{1'b0}},layer0_reg_4[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_4[3] <= { {8{1'b0}},layer0_reg_4[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_4[4] <= { {8{1'b0}},layer0_reg_4[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_4[5] <= { {8{1'b0}},layer1_reg_4[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_4[6] <= { {8{1'b0}},layer1_reg_4[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_4[7] <= { {8{1'b0}},layer1_reg_4[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_4[8] <= { {8{1'b0}},layer1_reg_4[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_4[9] <= { {8{1'b0}},layer1_reg_4[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_4[10] <= { {8{1'b0}},layer2_reg_4[7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_4[11] <= { {8{1'b0}},layer2_reg_4[15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_4[12] <= { {8{1'b0}},layer2_reg_4[23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_4[13] <= { {8{1'b0}},layer2_reg_4[31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_4[14] <= { {8{1'b0}},layer2_reg_4[39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_4[15] <= { {8{1'b0}},layer3_reg_4[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_4[16] <= { {8{1'b0}},layer3_reg_4[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_4[17] <= { {8{1'b0}},layer3_reg_4[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_4[18] <= { {8{1'b0}},layer3_reg_4[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_4[19] <= { {8{1'b0}},layer3_reg_4[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_4[20] <= { {8{1'b0}},layer4_reg_4[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_4[21] <= { {8{1'b0}},layer4_reg_4[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_4[22] <= { {8{1'b0}},layer4_reg_4[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_4[23] <= { {8{1'b0}},layer4_reg_4[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_4[24] <= { {8{1'b0}},layer4_reg_4[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_4;
reg  [15:0]  kernel_img_sum_2_4;
reg  [15:0]  kernel_img_sum_3_4;
reg  [15:0]  kernel_img_sum_4_4;
reg  [15:0]  kernel_img_sum_5_4;
reg  [15:0]  kernel_img_sum_6_4;
reg  [15:0]  kernel_img_sum_7_4;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_4 <= kernel_img_mul_4[0] + kernel_img_mul_4[1] + kernel_img_mul_4[2] + kernel_img_mul_4[3] + kernel_img_mul_4[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_4 <= kernel_img_mul_4[5] + kernel_img_mul_4[6] + kernel_img_mul_4[7] + kernel_img_mul_4[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_4 <= kernel_img_mul_4[9] + kernel_img_mul_4[10] + kernel_img_mul_4[11] + kernel_img_mul_4[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_4 <= kernel_img_mul_4[13] + kernel_img_mul_4[14] + kernel_img_mul_4[15] + kernel_img_mul_4[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_4 <= kernel_img_mul_4[17] + kernel_img_mul_4[18] + kernel_img_mul_4[19] + kernel_img_mul_4[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_4 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_4 <= kernel_img_mul_4[21] + kernel_img_mul_4[22] + kernel_img_mul_4[23] + kernel_img_mul_4[24];
  end
end
always@(*) begin
  kernel_img_sum_7_4 = kernel_img_sum_1_4 + kernel_img_sum_2_4 + kernel_img_sum_3_4 + kernel_img_sum_4_4 + kernel_img_sum_5_4 + kernel_img_sum_6_4;
end
reg  [15:0]  kernel_img_mul_5[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_5[0] <= 'd0;
    kernel_img_mul_5[1] <= 'd0;
    kernel_img_mul_5[2] <= 'd0;
    kernel_img_mul_5[3] <= 'd0;
    kernel_img_mul_5[4] <= 'd0;
    kernel_img_mul_5[5] <= 'd0;
    kernel_img_mul_5[6] <= 'd0;
    kernel_img_mul_5[7] <= 'd0;
    kernel_img_mul_5[8] <= 'd0;
    kernel_img_mul_5[9] <= 'd0;
    kernel_img_mul_5[10] <= 'd0;
    kernel_img_mul_5[11] <= 'd0;
    kernel_img_mul_5[12] <= 'd0;
    kernel_img_mul_5[13] <= 'd0;
    kernel_img_mul_5[14] <= 'd0;
    kernel_img_mul_5[15] <= 'd0;
    kernel_img_mul_5[16] <= 'd0;
    kernel_img_mul_5[17] <= 'd0;
    kernel_img_mul_5[18] <= 'd0;
    kernel_img_mul_5[19] <= 'd0;
    kernel_img_mul_5[20] <= 'd0;
    kernel_img_mul_5[21] <= 'd0;
    kernel_img_mul_5[22] <= 'd0;
    kernel_img_mul_5[23] <= 'd0;
    kernel_img_mul_5[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_5[0] <= { {8{1'b0}},layer0_reg_5[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_5[1] <= { {8{1'b0}},layer0_reg_5[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_5[2] <= { {8{1'b0}},layer0_reg_5[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_5[3] <= { {8{1'b0}},layer0_reg_5[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_5[4] <= { {8{1'b0}},layer0_reg_5[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_5[5] <= { {8{1'b0}},layer1_reg_5[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_5[6] <= { {8{1'b0}},layer1_reg_5[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_5[7] <= { {8{1'b0}},layer1_reg_5[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_5[8] <= { {8{1'b0}},layer1_reg_5[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_5[9] <= { {8{1'b0}},layer1_reg_5[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_5[10] <= { {8{1'b0}},layer2_reg_5[7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_5[11] <= { {8{1'b0}},layer2_reg_5[15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_5[12] <= { {8{1'b0}},layer2_reg_5[23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_5[13] <= { {8{1'b0}},layer2_reg_5[31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_5[14] <= { {8{1'b0}},layer2_reg_5[39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_5[15] <= { {8{1'b0}},layer3_reg_5[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_5[16] <= { {8{1'b0}},layer3_reg_5[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_5[17] <= { {8{1'b0}},layer3_reg_5[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_5[18] <= { {8{1'b0}},layer3_reg_5[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_5[19] <= { {8{1'b0}},layer3_reg_5[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_5[20] <= { {8{1'b0}},layer4_reg_5[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_5[21] <= { {8{1'b0}},layer4_reg_5[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_5[22] <= { {8{1'b0}},layer4_reg_5[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_5[23] <= { {8{1'b0}},layer4_reg_5[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_5[24] <= { {8{1'b0}},layer4_reg_5[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_5;
reg  [15:0]  kernel_img_sum_2_5;
reg  [15:0]  kernel_img_sum_3_5;
reg  [15:0]  kernel_img_sum_4_5;
reg  [15:0]  kernel_img_sum_5_5;
reg  [15:0]  kernel_img_sum_6_5;
reg  [15:0]  kernel_img_sum_7_5;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_5 <= kernel_img_mul_5[0] + kernel_img_mul_5[1] + kernel_img_mul_5[2] + kernel_img_mul_5[3] + kernel_img_mul_5[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_5 <= kernel_img_mul_5[5] + kernel_img_mul_5[6] + kernel_img_mul_5[7] + kernel_img_mul_5[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_5 <= kernel_img_mul_5[9] + kernel_img_mul_5[10] + kernel_img_mul_5[11] + kernel_img_mul_5[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_5 <= kernel_img_mul_5[13] + kernel_img_mul_5[14] + kernel_img_mul_5[15] + kernel_img_mul_5[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_5 <= kernel_img_mul_5[17] + kernel_img_mul_5[18] + kernel_img_mul_5[19] + kernel_img_mul_5[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_5 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_5 <= kernel_img_mul_5[21] + kernel_img_mul_5[22] + kernel_img_mul_5[23] + kernel_img_mul_5[24];
  end
end
always@(*) begin
  kernel_img_sum_7_5 = kernel_img_sum_1_5 + kernel_img_sum_2_5 + kernel_img_sum_3_5 + kernel_img_sum_4_5 + kernel_img_sum_5_5 + kernel_img_sum_6_5;
end
reg  [15:0]  kernel_img_mul_6[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_6[0] <= 'd0;
    kernel_img_mul_6[1] <= 'd0;
    kernel_img_mul_6[2] <= 'd0;
    kernel_img_mul_6[3] <= 'd0;
    kernel_img_mul_6[4] <= 'd0;
    kernel_img_mul_6[5] <= 'd0;
    kernel_img_mul_6[6] <= 'd0;
    kernel_img_mul_6[7] <= 'd0;
    kernel_img_mul_6[8] <= 'd0;
    kernel_img_mul_6[9] <= 'd0;
    kernel_img_mul_6[10] <= 'd0;
    kernel_img_mul_6[11] <= 'd0;
    kernel_img_mul_6[12] <= 'd0;
    kernel_img_mul_6[13] <= 'd0;
    kernel_img_mul_6[14] <= 'd0;
    kernel_img_mul_6[15] <= 'd0;
    kernel_img_mul_6[16] <= 'd0;
    kernel_img_mul_6[17] <= 'd0;
    kernel_img_mul_6[18] <= 'd0;
    kernel_img_mul_6[19] <= 'd0;
    kernel_img_mul_6[20] <= 'd0;
    kernel_img_mul_6[21] <= 'd0;
    kernel_img_mul_6[22] <= 'd0;
    kernel_img_mul_6[23] <= 'd0;
    kernel_img_mul_6[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_6[0] <= { {8{1'b0}},layer0_reg_6[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_6[1] <= { {8{1'b0}},layer0_reg_6[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_6[2] <= { {8{1'b0}},layer0_reg_6[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_6[3] <= { {8{1'b0}},layer0_reg_6[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_6[4] <= { {8{1'b0}},layer0_reg_6[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_6[5] <= { {8{1'b0}},layer1_reg_6[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_6[6] <= { {8{1'b0}},layer1_reg_6[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_6[7] <= { {8{1'b0}},layer1_reg_6[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_6[8] <= { {8{1'b0}},layer1_reg_6[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_6[9] <= { {8{1'b0}},layer1_reg_6[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_6[10] <= { {8{1'b0}},layer2_reg_6[7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_6[11] <= { {8{1'b0}},layer2_reg_6[15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_6[12] <= { {8{1'b0}},layer2_reg_6[23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_6[13] <= { {8{1'b0}},layer2_reg_6[31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_6[14] <= { {8{1'b0}},layer2_reg_6[39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_6[15] <= { {8{1'b0}},layer3_reg_6[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_6[16] <= { {8{1'b0}},layer3_reg_6[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_6[17] <= { {8{1'b0}},layer3_reg_6[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_6[18] <= { {8{1'b0}},layer3_reg_6[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_6[19] <= { {8{1'b0}},layer3_reg_6[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_6[20] <= { {8{1'b0}},layer4_reg_6[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_6[21] <= { {8{1'b0}},layer4_reg_6[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_6[22] <= { {8{1'b0}},layer4_reg_6[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_6[23] <= { {8{1'b0}},layer4_reg_6[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_6[24] <= { {8{1'b0}},layer4_reg_6[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_6;
reg  [15:0]  kernel_img_sum_2_6;
reg  [15:0]  kernel_img_sum_3_6;
reg  [15:0]  kernel_img_sum_4_6;
reg  [15:0]  kernel_img_sum_5_6;
reg  [15:0]  kernel_img_sum_6_6;
reg  [15:0]  kernel_img_sum_7_6;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_6 <= kernel_img_mul_6[0] + kernel_img_mul_6[1] + kernel_img_mul_6[2] + kernel_img_mul_6[3] + kernel_img_mul_6[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_6 <= kernel_img_mul_6[5] + kernel_img_mul_6[6] + kernel_img_mul_6[7] + kernel_img_mul_6[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_6 <= kernel_img_mul_6[9] + kernel_img_mul_6[10] + kernel_img_mul_6[11] + kernel_img_mul_6[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_6 <= kernel_img_mul_6[13] + kernel_img_mul_6[14] + kernel_img_mul_6[15] + kernel_img_mul_6[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_6 <= kernel_img_mul_6[17] + kernel_img_mul_6[18] + kernel_img_mul_6[19] + kernel_img_mul_6[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_6 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_6 <= kernel_img_mul_6[21] + kernel_img_mul_6[22] + kernel_img_mul_6[23] + kernel_img_mul_6[24];
  end
end
always@(*) begin
  kernel_img_sum_7_6 = kernel_img_sum_1_6 + kernel_img_sum_2_6 + kernel_img_sum_3_6 + kernel_img_sum_4_6 + kernel_img_sum_5_6 + kernel_img_sum_6_6;
end
reg  [15:0]  kernel_img_mul_7[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_7[0] <= 'd0;
    kernel_img_mul_7[1] <= 'd0;
    kernel_img_mul_7[2] <= 'd0;
    kernel_img_mul_7[3] <= 'd0;
    kernel_img_mul_7[4] <= 'd0;
    kernel_img_mul_7[5] <= 'd0;
    kernel_img_mul_7[6] <= 'd0;
    kernel_img_mul_7[7] <= 'd0;
    kernel_img_mul_7[8] <= 'd0;
    kernel_img_mul_7[9] <= 'd0;
    kernel_img_mul_7[10] <= 'd0;
    kernel_img_mul_7[11] <= 'd0;
    kernel_img_mul_7[12] <= 'd0;
    kernel_img_mul_7[13] <= 'd0;
    kernel_img_mul_7[14] <= 'd0;
    kernel_img_mul_7[15] <= 'd0;
    kernel_img_mul_7[16] <= 'd0;
    kernel_img_mul_7[17] <= 'd0;
    kernel_img_mul_7[18] <= 'd0;
    kernel_img_mul_7[19] <= 'd0;
    kernel_img_mul_7[20] <= 'd0;
    kernel_img_mul_7[21] <= 'd0;
    kernel_img_mul_7[22] <= 'd0;
    kernel_img_mul_7[23] <= 'd0;
    kernel_img_mul_7[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_7[0] <= { {8{1'b0}},layer0_reg_7[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_7[1] <= { {8{1'b0}},layer0_reg_7[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_7[2] <= { {8{1'b0}},layer0_reg_7[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_7[3] <= { {8{1'b0}},layer0_reg_7[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_7[4] <= { {8{1'b0}},layer0_reg_7[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_7[5] <= { {8{1'b0}},layer1_reg_7[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_7[6] <= { {8{1'b0}},layer1_reg_7[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_7[7] <= { {8{1'b0}},layer1_reg_7[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_7[8] <= { {8{1'b0}},layer1_reg_7[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_7[9] <= { {8{1'b0}},layer1_reg_7[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_7[10] <= { {8{1'b0}},layer2_reg_7[7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_7[11] <= { {8{1'b0}},layer2_reg_7[15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_7[12] <= { {8{1'b0}},layer2_reg_7[23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_7[13] <= { {8{1'b0}},layer2_reg_7[31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_7[14] <= { {8{1'b0}},layer2_reg_7[39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_7[15] <= { {8{1'b0}},layer3_reg_7[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_7[16] <= { {8{1'b0}},layer3_reg_7[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_7[17] <= { {8{1'b0}},layer3_reg_7[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_7[18] <= { {8{1'b0}},layer3_reg_7[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_7[19] <= { {8{1'b0}},layer3_reg_7[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_7[20] <= { {8{1'b0}},layer4_reg_7[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_7[21] <= { {8{1'b0}},layer4_reg_7[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_7[22] <= { {8{1'b0}},layer4_reg_7[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_7[23] <= { {8{1'b0}},layer4_reg_7[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_7[24] <= { {8{1'b0}},layer4_reg_7[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_7;
reg  [15:0]  kernel_img_sum_2_7;
reg  [15:0]  kernel_img_sum_3_7;
reg  [15:0]  kernel_img_sum_4_7;
reg  [15:0]  kernel_img_sum_5_7;
reg  [15:0]  kernel_img_sum_6_7;
reg  [15:0]  kernel_img_sum_7_7;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_7 <= kernel_img_mul_7[0] + kernel_img_mul_7[1] + kernel_img_mul_7[2] + kernel_img_mul_7[3] + kernel_img_mul_7[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_7 <= kernel_img_mul_7[5] + kernel_img_mul_7[6] + kernel_img_mul_7[7] + kernel_img_mul_7[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_7 <= kernel_img_mul_7[9] + kernel_img_mul_7[10] + kernel_img_mul_7[11] + kernel_img_mul_7[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_7 <= kernel_img_mul_7[13] + kernel_img_mul_7[14] + kernel_img_mul_7[15] + kernel_img_mul_7[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_7 <= kernel_img_mul_7[17] + kernel_img_mul_7[18] + kernel_img_mul_7[19] + kernel_img_mul_7[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_7 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_7 <= kernel_img_mul_7[21] + kernel_img_mul_7[22] + kernel_img_mul_7[23] + kernel_img_mul_7[24];
  end
end
always@(*) begin
  kernel_img_sum_7_7 = kernel_img_sum_1_7 + kernel_img_sum_2_7 + kernel_img_sum_3_7 + kernel_img_sum_4_7 + kernel_img_sum_5_7 + kernel_img_sum_6_7;
end
reg  [15:0]  kernel_img_mul_8[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_8[0] <= 'd0;
    kernel_img_mul_8[1] <= 'd0;
    kernel_img_mul_8[2] <= 'd0;
    kernel_img_mul_8[3] <= 'd0;
    kernel_img_mul_8[4] <= 'd0;
    kernel_img_mul_8[5] <= 'd0;
    kernel_img_mul_8[6] <= 'd0;
    kernel_img_mul_8[7] <= 'd0;
    kernel_img_mul_8[8] <= 'd0;
    kernel_img_mul_8[9] <= 'd0;
    kernel_img_mul_8[10] <= 'd0;
    kernel_img_mul_8[11] <= 'd0;
    kernel_img_mul_8[12] <= 'd0;
    kernel_img_mul_8[13] <= 'd0;
    kernel_img_mul_8[14] <= 'd0;
    kernel_img_mul_8[15] <= 'd0;
    kernel_img_mul_8[16] <= 'd0;
    kernel_img_mul_8[17] <= 'd0;
    kernel_img_mul_8[18] <= 'd0;
    kernel_img_mul_8[19] <= 'd0;
    kernel_img_mul_8[20] <= 'd0;
    kernel_img_mul_8[21] <= 'd0;
    kernel_img_mul_8[22] <= 'd0;
    kernel_img_mul_8[23] <= 'd0;
    kernel_img_mul_8[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_8[0] <= { {8{1'b0}},layer0_reg_8[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_8[1] <= { {8{1'b0}},layer0_reg_8[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_8[2] <= { {8{1'b0}},layer0_reg_8[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_8[3] <= { {8{1'b0}},layer0_reg_8[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_8[4] <= { {8{1'b0}},layer0_reg_8[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_8[5] <= { {8{1'b0}},layer1_reg_8[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_8[6] <= { {8{1'b0}},layer1_reg_8[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_8[7] <= { {8{1'b0}},layer1_reg_8[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_8[8] <= { {8{1'b0}},layer1_reg_8[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_8[9] <= { {8{1'b0}},layer1_reg_8[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_8[10] <= { {8{1'b0}},layer2_reg_8[7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_8[11] <= { {8{1'b0}},layer2_reg_8[15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_8[12] <= { {8{1'b0}},layer2_reg_8[23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_8[13] <= { {8{1'b0}},layer2_reg_8[31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_8[14] <= { {8{1'b0}},layer2_reg_8[39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_8[15] <= { {8{1'b0}},layer3_reg_8[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_8[16] <= { {8{1'b0}},layer3_reg_8[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_8[17] <= { {8{1'b0}},layer3_reg_8[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_8[18] <= { {8{1'b0}},layer3_reg_8[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_8[19] <= { {8{1'b0}},layer3_reg_8[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_8[20] <= { {8{1'b0}},layer4_reg_8[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_8[21] <= { {8{1'b0}},layer4_reg_8[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_8[22] <= { {8{1'b0}},layer4_reg_8[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_8[23] <= { {8{1'b0}},layer4_reg_8[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_8[24] <= { {8{1'b0}},layer4_reg_8[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_8;
reg  [15:0]  kernel_img_sum_2_8;
reg  [15:0]  kernel_img_sum_3_8;
reg  [15:0]  kernel_img_sum_4_8;
reg  [15:0]  kernel_img_sum_5_8;
reg  [15:0]  kernel_img_sum_6_8;
reg  [15:0]  kernel_img_sum_7_8;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_8 <= kernel_img_mul_8[0] + kernel_img_mul_8[1] + kernel_img_mul_8[2] + kernel_img_mul_8[3] + kernel_img_mul_8[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_8 <= kernel_img_mul_8[5] + kernel_img_mul_8[6] + kernel_img_mul_8[7] + kernel_img_mul_8[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_8 <= kernel_img_mul_8[9] + kernel_img_mul_8[10] + kernel_img_mul_8[11] + kernel_img_mul_8[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_8 <= kernel_img_mul_8[13] + kernel_img_mul_8[14] + kernel_img_mul_8[15] + kernel_img_mul_8[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_8 <= kernel_img_mul_8[17] + kernel_img_mul_8[18] + kernel_img_mul_8[19] + kernel_img_mul_8[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_8 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_8 <= kernel_img_mul_8[21] + kernel_img_mul_8[22] + kernel_img_mul_8[23] + kernel_img_mul_8[24];
  end
end
always@(*) begin
  kernel_img_sum_7_8 = kernel_img_sum_1_8 + kernel_img_sum_2_8 + kernel_img_sum_3_8 + kernel_img_sum_4_8 + kernel_img_sum_5_8 + kernel_img_sum_6_8;
end
reg  [15:0]  kernel_img_mul_9[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_9[0] <= 'd0;
    kernel_img_mul_9[1] <= 'd0;
    kernel_img_mul_9[2] <= 'd0;
    kernel_img_mul_9[3] <= 'd0;
    kernel_img_mul_9[4] <= 'd0;
    kernel_img_mul_9[5] <= 'd0;
    kernel_img_mul_9[6] <= 'd0;
    kernel_img_mul_9[7] <= 'd0;
    kernel_img_mul_9[8] <= 'd0;
    kernel_img_mul_9[9] <= 'd0;
    kernel_img_mul_9[10] <= 'd0;
    kernel_img_mul_9[11] <= 'd0;
    kernel_img_mul_9[12] <= 'd0;
    kernel_img_mul_9[13] <= 'd0;
    kernel_img_mul_9[14] <= 'd0;
    kernel_img_mul_9[15] <= 'd0;
    kernel_img_mul_9[16] <= 'd0;
    kernel_img_mul_9[17] <= 'd0;
    kernel_img_mul_9[18] <= 'd0;
    kernel_img_mul_9[19] <= 'd0;
    kernel_img_mul_9[20] <= 'd0;
    kernel_img_mul_9[21] <= 'd0;
    kernel_img_mul_9[22] <= 'd0;
    kernel_img_mul_9[23] <= 'd0;
    kernel_img_mul_9[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_9[0] <= { {8{1'b0}},layer0_reg_9[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_9[1] <= { {8{1'b0}},layer0_reg_9[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_9[2] <= { {8{1'b0}},layer0_reg_9[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_9[3] <= { {8{1'b0}},layer0_reg_9[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_9[4] <= { {8{1'b0}},layer0_reg_9[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_9[5] <= { {8{1'b0}},layer1_reg_9[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_9[6] <= { {8{1'b0}},layer1_reg_9[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_9[7] <= { {8{1'b0}},layer1_reg_9[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_9[8] <= { {8{1'b0}},layer1_reg_9[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_9[9] <= { {8{1'b0}},layer1_reg_9[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_9[10] <= { {8{1'b0}},layer2_reg_9[7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_9[11] <= { {8{1'b0}},layer2_reg_9[15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_9[12] <= { {8{1'b0}},layer2_reg_9[23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_9[13] <= { {8{1'b0}},layer2_reg_9[31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_9[14] <= { {8{1'b0}},layer2_reg_9[39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_9[15] <= { {8{1'b0}},layer3_reg_9[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_9[16] <= { {8{1'b0}},layer3_reg_9[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_9[17] <= { {8{1'b0}},layer3_reg_9[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_9[18] <= { {8{1'b0}},layer3_reg_9[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_9[19] <= { {8{1'b0}},layer3_reg_9[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_9[20] <= { {8{1'b0}},layer4_reg_9[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_9[21] <= { {8{1'b0}},layer4_reg_9[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_9[22] <= { {8{1'b0}},layer4_reg_9[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_9[23] <= { {8{1'b0}},layer4_reg_9[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_9[24] <= { {8{1'b0}},layer4_reg_9[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_9;
reg  [15:0]  kernel_img_sum_2_9;
reg  [15:0]  kernel_img_sum_3_9;
reg  [15:0]  kernel_img_sum_4_9;
reg  [15:0]  kernel_img_sum_5_9;
reg  [15:0]  kernel_img_sum_6_9;
reg  [15:0]  kernel_img_sum_7_9;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_9 <= kernel_img_mul_9[0] + kernel_img_mul_9[1] + kernel_img_mul_9[2] + kernel_img_mul_9[3] + kernel_img_mul_9[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_9 <= kernel_img_mul_9[5] + kernel_img_mul_9[6] + kernel_img_mul_9[7] + kernel_img_mul_9[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_9 <= kernel_img_mul_9[9] + kernel_img_mul_9[10] + kernel_img_mul_9[11] + kernel_img_mul_9[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_9 <= kernel_img_mul_9[13] + kernel_img_mul_9[14] + kernel_img_mul_9[15] + kernel_img_mul_9[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_9 <= kernel_img_mul_9[17] + kernel_img_mul_9[18] + kernel_img_mul_9[19] + kernel_img_mul_9[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_9 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_9 <= kernel_img_mul_9[21] + kernel_img_mul_9[22] + kernel_img_mul_9[23] + kernel_img_mul_9[24];
  end
end
always@(*) begin
  kernel_img_sum_7_9 = kernel_img_sum_1_9 + kernel_img_sum_2_9 + kernel_img_sum_3_9 + kernel_img_sum_4_9 + kernel_img_sum_5_9 + kernel_img_sum_6_9;
end
reg  [15:0]  kernel_img_mul_10[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_10[0] <= 'd0;
    kernel_img_mul_10[1] <= 'd0;
    kernel_img_mul_10[2] <= 'd0;
    kernel_img_mul_10[3] <= 'd0;
    kernel_img_mul_10[4] <= 'd0;
    kernel_img_mul_10[5] <= 'd0;
    kernel_img_mul_10[6] <= 'd0;
    kernel_img_mul_10[7] <= 'd0;
    kernel_img_mul_10[8] <= 'd0;
    kernel_img_mul_10[9] <= 'd0;
    kernel_img_mul_10[10] <= 'd0;
    kernel_img_mul_10[11] <= 'd0;
    kernel_img_mul_10[12] <= 'd0;
    kernel_img_mul_10[13] <= 'd0;
    kernel_img_mul_10[14] <= 'd0;
    kernel_img_mul_10[15] <= 'd0;
    kernel_img_mul_10[16] <= 'd0;
    kernel_img_mul_10[17] <= 'd0;
    kernel_img_mul_10[18] <= 'd0;
    kernel_img_mul_10[19] <= 'd0;
    kernel_img_mul_10[20] <= 'd0;
    kernel_img_mul_10[21] <= 'd0;
    kernel_img_mul_10[22] <= 'd0;
    kernel_img_mul_10[23] <= 'd0;
    kernel_img_mul_10[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_10[0] <= { {8{1'b0}},layer0_reg_10[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_10[1] <= { {8{1'b0}},layer0_reg_10[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_10[2] <= { {8{1'b0}},layer0_reg_10[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_10[3] <= { {8{1'b0}},layer0_reg_10[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_10[4] <= { {8{1'b0}},layer0_reg_10[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_10[5] <= { {8{1'b0}},layer1_reg_10[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_10[6] <= { {8{1'b0}},layer1_reg_10[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_10[7] <= { {8{1'b0}},layer1_reg_10[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_10[8] <= { {8{1'b0}},layer1_reg_10[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_10[9] <= { {8{1'b0}},layer1_reg_10[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_10[10] <= { {8{1'b0}},layer2_reg_10[7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_10[11] <= { {8{1'b0}},layer2_reg_10[15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_10[12] <= { {8{1'b0}},layer2_reg_10[23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_10[13] <= { {8{1'b0}},layer2_reg_10[31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_10[14] <= { {8{1'b0}},layer2_reg_10[39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_10[15] <= { {8{1'b0}},layer3_reg_10[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_10[16] <= { {8{1'b0}},layer3_reg_10[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_10[17] <= { {8{1'b0}},layer3_reg_10[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_10[18] <= { {8{1'b0}},layer3_reg_10[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_10[19] <= { {8{1'b0}},layer3_reg_10[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_10[20] <= { {8{1'b0}},layer4_reg_10[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_10[21] <= { {8{1'b0}},layer4_reg_10[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_10[22] <= { {8{1'b0}},layer4_reg_10[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_10[23] <= { {8{1'b0}},layer4_reg_10[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_10[24] <= { {8{1'b0}},layer4_reg_10[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_10;
reg  [15:0]  kernel_img_sum_2_10;
reg  [15:0]  kernel_img_sum_3_10;
reg  [15:0]  kernel_img_sum_4_10;
reg  [15:0]  kernel_img_sum_5_10;
reg  [15:0]  kernel_img_sum_6_10;
reg  [15:0]  kernel_img_sum_7_10;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_10 <= kernel_img_mul_10[0] + kernel_img_mul_10[1] + kernel_img_mul_10[2] + kernel_img_mul_10[3] + kernel_img_mul_10[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_10 <= kernel_img_mul_10[5] + kernel_img_mul_10[6] + kernel_img_mul_10[7] + kernel_img_mul_10[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_10 <= kernel_img_mul_10[9] + kernel_img_mul_10[10] + kernel_img_mul_10[11] + kernel_img_mul_10[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_10 <= kernel_img_mul_10[13] + kernel_img_mul_10[14] + kernel_img_mul_10[15] + kernel_img_mul_10[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_10 <= kernel_img_mul_10[17] + kernel_img_mul_10[18] + kernel_img_mul_10[19] + kernel_img_mul_10[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_10 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_10 <= kernel_img_mul_10[21] + kernel_img_mul_10[22] + kernel_img_mul_10[23] + kernel_img_mul_10[24];
  end
end
always@(*) begin
  kernel_img_sum_7_10 = kernel_img_sum_1_10 + kernel_img_sum_2_10 + kernel_img_sum_3_10 + kernel_img_sum_4_10 + kernel_img_sum_5_10 + kernel_img_sum_6_10;
end
reg  [15:0]  kernel_img_mul_11[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_11[0] <= 'd0;
    kernel_img_mul_11[1] <= 'd0;
    kernel_img_mul_11[2] <= 'd0;
    kernel_img_mul_11[3] <= 'd0;
    kernel_img_mul_11[4] <= 'd0;
    kernel_img_mul_11[5] <= 'd0;
    kernel_img_mul_11[6] <= 'd0;
    kernel_img_mul_11[7] <= 'd0;
    kernel_img_mul_11[8] <= 'd0;
    kernel_img_mul_11[9] <= 'd0;
    kernel_img_mul_11[10] <= 'd0;
    kernel_img_mul_11[11] <= 'd0;
    kernel_img_mul_11[12] <= 'd0;
    kernel_img_mul_11[13] <= 'd0;
    kernel_img_mul_11[14] <= 'd0;
    kernel_img_mul_11[15] <= 'd0;
    kernel_img_mul_11[16] <= 'd0;
    kernel_img_mul_11[17] <= 'd0;
    kernel_img_mul_11[18] <= 'd0;
    kernel_img_mul_11[19] <= 'd0;
    kernel_img_mul_11[20] <= 'd0;
    kernel_img_mul_11[21] <= 'd0;
    kernel_img_mul_11[22] <= 'd0;
    kernel_img_mul_11[23] <= 'd0;
    kernel_img_mul_11[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_11[0] <= { {8{1'b0}},layer0_reg_11[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_11[1] <= { {8{1'b0}},layer0_reg_11[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_11[2] <= { {8{1'b0}},layer0_reg_11[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_11[3] <= { {8{1'b0}},layer0_reg_11[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_11[4] <= { {8{1'b0}},layer0_reg_11[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_11[5] <= { {8{1'b0}},layer1_reg_11[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_11[6] <= { {8{1'b0}},layer1_reg_11[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_11[7] <= { {8{1'b0}},layer1_reg_11[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_11[8] <= { {8{1'b0}},layer1_reg_11[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_11[9] <= { {8{1'b0}},layer1_reg_11[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_11[10] <= { {8{1'b0}},layer2_reg_11[7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_11[11] <= { {8{1'b0}},layer2_reg_11[15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_11[12] <= { {8{1'b0}},layer2_reg_11[23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_11[13] <= { {8{1'b0}},layer2_reg_11[31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_11[14] <= { {8{1'b0}},layer2_reg_11[39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_11[15] <= { {8{1'b0}},layer3_reg_11[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_11[16] <= { {8{1'b0}},layer3_reg_11[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_11[17] <= { {8{1'b0}},layer3_reg_11[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_11[18] <= { {8{1'b0}},layer3_reg_11[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_11[19] <= { {8{1'b0}},layer3_reg_11[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_11[20] <= { {8{1'b0}},layer4_reg_11[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_11[21] <= { {8{1'b0}},layer4_reg_11[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_11[22] <= { {8{1'b0}},layer4_reg_11[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_11[23] <= { {8{1'b0}},layer4_reg_11[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_11[24] <= { {8{1'b0}},layer4_reg_11[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_11;
reg  [15:0]  kernel_img_sum_2_11;
reg  [15:0]  kernel_img_sum_3_11;
reg  [15:0]  kernel_img_sum_4_11;
reg  [15:0]  kernel_img_sum_5_11;
reg  [15:0]  kernel_img_sum_6_11;
reg  [15:0]  kernel_img_sum_7_11;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_11 <= kernel_img_mul_11[0] + kernel_img_mul_11[1] + kernel_img_mul_11[2] + kernel_img_mul_11[3] + kernel_img_mul_11[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_11 <= kernel_img_mul_11[5] + kernel_img_mul_11[6] + kernel_img_mul_11[7] + kernel_img_mul_11[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_11 <= kernel_img_mul_11[9] + kernel_img_mul_11[10] + kernel_img_mul_11[11] + kernel_img_mul_11[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_11 <= kernel_img_mul_11[13] + kernel_img_mul_11[14] + kernel_img_mul_11[15] + kernel_img_mul_11[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_11 <= kernel_img_mul_11[17] + kernel_img_mul_11[18] + kernel_img_mul_11[19] + kernel_img_mul_11[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_11 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_11 <= kernel_img_mul_11[21] + kernel_img_mul_11[22] + kernel_img_mul_11[23] + kernel_img_mul_11[24];
  end
end
always@(*) begin
  kernel_img_sum_7_11 = kernel_img_sum_1_11 + kernel_img_sum_2_11 + kernel_img_sum_3_11 + kernel_img_sum_4_11 + kernel_img_sum_5_11 + kernel_img_sum_6_11;
end
reg  [15:0]  kernel_img_mul_12[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_12[0] <= 'd0;
    kernel_img_mul_12[1] <= 'd0;
    kernel_img_mul_12[2] <= 'd0;
    kernel_img_mul_12[3] <= 'd0;
    kernel_img_mul_12[4] <= 'd0;
    kernel_img_mul_12[5] <= 'd0;
    kernel_img_mul_12[6] <= 'd0;
    kernel_img_mul_12[7] <= 'd0;
    kernel_img_mul_12[8] <= 'd0;
    kernel_img_mul_12[9] <= 'd0;
    kernel_img_mul_12[10] <= 'd0;
    kernel_img_mul_12[11] <= 'd0;
    kernel_img_mul_12[12] <= 'd0;
    kernel_img_mul_12[13] <= 'd0;
    kernel_img_mul_12[14] <= 'd0;
    kernel_img_mul_12[15] <= 'd0;
    kernel_img_mul_12[16] <= 'd0;
    kernel_img_mul_12[17] <= 'd0;
    kernel_img_mul_12[18] <= 'd0;
    kernel_img_mul_12[19] <= 'd0;
    kernel_img_mul_12[20] <= 'd0;
    kernel_img_mul_12[21] <= 'd0;
    kernel_img_mul_12[22] <= 'd0;
    kernel_img_mul_12[23] <= 'd0;
    kernel_img_mul_12[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_12[0] <= { {8{1'b0}},layer0_reg_12[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_12[1] <= { {8{1'b0}},layer0_reg_12[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_12[2] <= { {8{1'b0}},layer0_reg_12[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_12[3] <= { {8{1'b0}},layer0_reg_12[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_12[4] <= { {8{1'b0}},layer0_reg_12[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_12[5] <= { {8{1'b0}},layer1_reg_12[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_12[6] <= { {8{1'b0}},layer1_reg_12[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_12[7] <= { {8{1'b0}},layer1_reg_12[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_12[8] <= { {8{1'b0}},layer1_reg_12[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_12[9] <= { {8{1'b0}},layer1_reg_12[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_12[10] <= { {8{1'b0}},layer2_reg_12[7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_12[11] <= { {8{1'b0}},layer2_reg_12[15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_12[12] <= { {8{1'b0}},layer2_reg_12[23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_12[13] <= { {8{1'b0}},layer2_reg_12[31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_12[14] <= { {8{1'b0}},layer2_reg_12[39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_12[15] <= { {8{1'b0}},layer3_reg_12[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_12[16] <= { {8{1'b0}},layer3_reg_12[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_12[17] <= { {8{1'b0}},layer3_reg_12[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_12[18] <= { {8{1'b0}},layer3_reg_12[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_12[19] <= { {8{1'b0}},layer3_reg_12[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_12[20] <= { {8{1'b0}},layer4_reg_12[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_12[21] <= { {8{1'b0}},layer4_reg_12[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_12[22] <= { {8{1'b0}},layer4_reg_12[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_12[23] <= { {8{1'b0}},layer4_reg_12[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_12[24] <= { {8{1'b0}},layer4_reg_12[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_12;
reg  [15:0]  kernel_img_sum_2_12;
reg  [15:0]  kernel_img_sum_3_12;
reg  [15:0]  kernel_img_sum_4_12;
reg  [15:0]  kernel_img_sum_5_12;
reg  [15:0]  kernel_img_sum_6_12;
reg  [15:0]  kernel_img_sum_7_12;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_12 <= kernel_img_mul_12[0] + kernel_img_mul_12[1] + kernel_img_mul_12[2] + kernel_img_mul_12[3] + kernel_img_mul_12[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_12 <= kernel_img_mul_12[5] + kernel_img_mul_12[6] + kernel_img_mul_12[7] + kernel_img_mul_12[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_12 <= kernel_img_mul_12[9] + kernel_img_mul_12[10] + kernel_img_mul_12[11] + kernel_img_mul_12[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_12 <= kernel_img_mul_12[13] + kernel_img_mul_12[14] + kernel_img_mul_12[15] + kernel_img_mul_12[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_12 <= kernel_img_mul_12[17] + kernel_img_mul_12[18] + kernel_img_mul_12[19] + kernel_img_mul_12[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_12 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_12 <= kernel_img_mul_12[21] + kernel_img_mul_12[22] + kernel_img_mul_12[23] + kernel_img_mul_12[24];
  end
end
always@(*) begin
  kernel_img_sum_7_12 = kernel_img_sum_1_12 + kernel_img_sum_2_12 + kernel_img_sum_3_12 + kernel_img_sum_4_12 + kernel_img_sum_5_12 + kernel_img_sum_6_12;
end
reg  [15:0]  kernel_img_mul_13[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_13[0] <= 'd0;
    kernel_img_mul_13[1] <= 'd0;
    kernel_img_mul_13[2] <= 'd0;
    kernel_img_mul_13[3] <= 'd0;
    kernel_img_mul_13[4] <= 'd0;
    kernel_img_mul_13[5] <= 'd0;
    kernel_img_mul_13[6] <= 'd0;
    kernel_img_mul_13[7] <= 'd0;
    kernel_img_mul_13[8] <= 'd0;
    kernel_img_mul_13[9] <= 'd0;
    kernel_img_mul_13[10] <= 'd0;
    kernel_img_mul_13[11] <= 'd0;
    kernel_img_mul_13[12] <= 'd0;
    kernel_img_mul_13[13] <= 'd0;
    kernel_img_mul_13[14] <= 'd0;
    kernel_img_mul_13[15] <= 'd0;
    kernel_img_mul_13[16] <= 'd0;
    kernel_img_mul_13[17] <= 'd0;
    kernel_img_mul_13[18] <= 'd0;
    kernel_img_mul_13[19] <= 'd0;
    kernel_img_mul_13[20] <= 'd0;
    kernel_img_mul_13[21] <= 'd0;
    kernel_img_mul_13[22] <= 'd0;
    kernel_img_mul_13[23] <= 'd0;
    kernel_img_mul_13[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_13[0] <= { {8{1'b0}},layer0_reg_13[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_13[1] <= { {8{1'b0}},layer0_reg_13[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_13[2] <= { {8{1'b0}},layer0_reg_13[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_13[3] <= { {8{1'b0}},layer0_reg_13[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_13[4] <= { {8{1'b0}},layer0_reg_13[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_13[5] <= { {8{1'b0}},layer1_reg_13[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_13[6] <= { {8{1'b0}},layer1_reg_13[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_13[7] <= { {8{1'b0}},layer1_reg_13[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_13[8] <= { {8{1'b0}},layer1_reg_13[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_13[9] <= { {8{1'b0}},layer1_reg_13[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_13[10] <= { {8{1'b0}},layer2_reg_13[7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_13[11] <= { {8{1'b0}},layer2_reg_13[15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_13[12] <= { {8{1'b0}},layer2_reg_13[23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_13[13] <= { {8{1'b0}},layer2_reg_13[31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_13[14] <= { {8{1'b0}},layer2_reg_13[39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_13[15] <= { {8{1'b0}},layer3_reg_13[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_13[16] <= { {8{1'b0}},layer3_reg_13[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_13[17] <= { {8{1'b0}},layer3_reg_13[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_13[18] <= { {8{1'b0}},layer3_reg_13[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_13[19] <= { {8{1'b0}},layer3_reg_13[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_13[20] <= { {8{1'b0}},layer4_reg_13[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_13[21] <= { {8{1'b0}},layer4_reg_13[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_13[22] <= { {8{1'b0}},layer4_reg_13[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_13[23] <= { {8{1'b0}},layer4_reg_13[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_13[24] <= { {8{1'b0}},layer4_reg_13[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_13;
reg  [15:0]  kernel_img_sum_2_13;
reg  [15:0]  kernel_img_sum_3_13;
reg  [15:0]  kernel_img_sum_4_13;
reg  [15:0]  kernel_img_sum_5_13;
reg  [15:0]  kernel_img_sum_6_13;
reg  [15:0]  kernel_img_sum_7_13;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_13 <= kernel_img_mul_13[0] + kernel_img_mul_13[1] + kernel_img_mul_13[2] + kernel_img_mul_13[3] + kernel_img_mul_13[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_13 <= kernel_img_mul_13[5] + kernel_img_mul_13[6] + kernel_img_mul_13[7] + kernel_img_mul_13[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_13 <= kernel_img_mul_13[9] + kernel_img_mul_13[10] + kernel_img_mul_13[11] + kernel_img_mul_13[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_13 <= kernel_img_mul_13[13] + kernel_img_mul_13[14] + kernel_img_mul_13[15] + kernel_img_mul_13[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_13 <= kernel_img_mul_13[17] + kernel_img_mul_13[18] + kernel_img_mul_13[19] + kernel_img_mul_13[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_13 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_13 <= kernel_img_mul_13[21] + kernel_img_mul_13[22] + kernel_img_mul_13[23] + kernel_img_mul_13[24];
  end
end
always@(*) begin
  kernel_img_sum_7_13 = kernel_img_sum_1_13 + kernel_img_sum_2_13 + kernel_img_sum_3_13 + kernel_img_sum_4_13 + kernel_img_sum_5_13 + kernel_img_sum_6_13;
end
reg  [15:0]  kernel_img_mul_14[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_14[0] <= 'd0;
    kernel_img_mul_14[1] <= 'd0;
    kernel_img_mul_14[2] <= 'd0;
    kernel_img_mul_14[3] <= 'd0;
    kernel_img_mul_14[4] <= 'd0;
    kernel_img_mul_14[5] <= 'd0;
    kernel_img_mul_14[6] <= 'd0;
    kernel_img_mul_14[7] <= 'd0;
    kernel_img_mul_14[8] <= 'd0;
    kernel_img_mul_14[9] <= 'd0;
    kernel_img_mul_14[10] <= 'd0;
    kernel_img_mul_14[11] <= 'd0;
    kernel_img_mul_14[12] <= 'd0;
    kernel_img_mul_14[13] <= 'd0;
    kernel_img_mul_14[14] <= 'd0;
    kernel_img_mul_14[15] <= 'd0;
    kernel_img_mul_14[16] <= 'd0;
    kernel_img_mul_14[17] <= 'd0;
    kernel_img_mul_14[18] <= 'd0;
    kernel_img_mul_14[19] <= 'd0;
    kernel_img_mul_14[20] <= 'd0;
    kernel_img_mul_14[21] <= 'd0;
    kernel_img_mul_14[22] <= 'd0;
    kernel_img_mul_14[23] <= 'd0;
    kernel_img_mul_14[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_14[0] <= { {8{1'b0}},layer0_reg_14[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_14[1] <= { {8{1'b0}},layer0_reg_14[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_14[2] <= { {8{1'b0}},layer0_reg_14[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_14[3] <= { {8{1'b0}},layer0_reg_14[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_14[4] <= { {8{1'b0}},layer0_reg_14[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_14[5] <= { {8{1'b0}},layer1_reg_14[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_14[6] <= { {8{1'b0}},layer1_reg_14[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_14[7] <= { {8{1'b0}},layer1_reg_14[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_14[8] <= { {8{1'b0}},layer1_reg_14[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_14[9] <= { {8{1'b0}},layer1_reg_14[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_14[10] <= { {8{1'b0}},layer2_reg_14[7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_14[11] <= { {8{1'b0}},layer2_reg_14[15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_14[12] <= { {8{1'b0}},layer2_reg_14[23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_14[13] <= { {8{1'b0}},layer2_reg_14[31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_14[14] <= { {8{1'b0}},layer2_reg_14[39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_14[15] <= { {8{1'b0}},layer3_reg_14[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_14[16] <= { {8{1'b0}},layer3_reg_14[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_14[17] <= { {8{1'b0}},layer3_reg_14[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_14[18] <= { {8{1'b0}},layer3_reg_14[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_14[19] <= { {8{1'b0}},layer3_reg_14[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_14[20] <= { {8{1'b0}},layer4_reg_14[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_14[21] <= { {8{1'b0}},layer4_reg_14[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_14[22] <= { {8{1'b0}},layer4_reg_14[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_14[23] <= { {8{1'b0}},layer4_reg_14[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_14[24] <= { {8{1'b0}},layer4_reg_14[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_14;
reg  [15:0]  kernel_img_sum_2_14;
reg  [15:0]  kernel_img_sum_3_14;
reg  [15:0]  kernel_img_sum_4_14;
reg  [15:0]  kernel_img_sum_5_14;
reg  [15:0]  kernel_img_sum_6_14;
reg  [15:0]  kernel_img_sum_7_14;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_14 <= kernel_img_mul_14[0] + kernel_img_mul_14[1] + kernel_img_mul_14[2] + kernel_img_mul_14[3] + kernel_img_mul_14[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_14 <= kernel_img_mul_14[5] + kernel_img_mul_14[6] + kernel_img_mul_14[7] + kernel_img_mul_14[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_14 <= kernel_img_mul_14[9] + kernel_img_mul_14[10] + kernel_img_mul_14[11] + kernel_img_mul_14[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_14 <= kernel_img_mul_14[13] + kernel_img_mul_14[14] + kernel_img_mul_14[15] + kernel_img_mul_14[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_14 <= kernel_img_mul_14[17] + kernel_img_mul_14[18] + kernel_img_mul_14[19] + kernel_img_mul_14[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_14 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_14 <= kernel_img_mul_14[21] + kernel_img_mul_14[22] + kernel_img_mul_14[23] + kernel_img_mul_14[24];
  end
end
always@(*) begin
  kernel_img_sum_7_14 = kernel_img_sum_1_14 + kernel_img_sum_2_14 + kernel_img_sum_3_14 + kernel_img_sum_4_14 + kernel_img_sum_5_14 + kernel_img_sum_6_14;
end
reg  [15:0]  kernel_img_mul_15[0:24];
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_mul_15[0] <= 'd0;
    kernel_img_mul_15[1] <= 'd0;
    kernel_img_mul_15[2] <= 'd0;
    kernel_img_mul_15[3] <= 'd0;
    kernel_img_mul_15[4] <= 'd0;
    kernel_img_mul_15[5] <= 'd0;
    kernel_img_mul_15[6] <= 'd0;
    kernel_img_mul_15[7] <= 'd0;
    kernel_img_mul_15[8] <= 'd0;
    kernel_img_mul_15[9] <= 'd0;
    kernel_img_mul_15[10] <= 'd0;
    kernel_img_mul_15[11] <= 'd0;
    kernel_img_mul_15[12] <= 'd0;
    kernel_img_mul_15[13] <= 'd0;
    kernel_img_mul_15[14] <= 'd0;
    kernel_img_mul_15[15] <= 'd0;
    kernel_img_mul_15[16] <= 'd0;
    kernel_img_mul_15[17] <= 'd0;
    kernel_img_mul_15[18] <= 'd0;
    kernel_img_mul_15[19] <= 'd0;
    kernel_img_mul_15[20] <= 'd0;
    kernel_img_mul_15[21] <= 'd0;
    kernel_img_mul_15[22] <= 'd0;
    kernel_img_mul_15[23] <= 'd0;
    kernel_img_mul_15[24] <= 'd0;
  end
  else if(current_state==ST_MUL) begin
    kernel_img_mul_15[0] <= { {8{1'b0}},layer0_reg_15[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_15[1] <= { {8{1'b0}},layer0_reg_15[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_15[2] <= { {8{1'b0}},layer0_reg_15[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_15[3] <= { {8{1'b0}},layer0_reg_15[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_15[4] <= { {8{1'b0}},layer0_reg_15[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
    kernel_img_mul_15[5] <= { {8{1'b0}},layer1_reg_15[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_15[6] <= { {8{1'b0}},layer1_reg_15[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_15[7] <= { {8{1'b0}},layer1_reg_15[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_15[8] <= { {8{1'b0}},layer1_reg_15[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_15[9] <= { {8{1'b0}},layer1_reg_15[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_15[10] <= { {8{1'b0}},layer2_reg_15[7:0]} * { {8{1'b0}}, G_Kernel_5x5_2[7:0]};
    kernel_img_mul_15[11] <= { {8{1'b0}},layer2_reg_15[15:8]} * { {8{1'b0}}, G_Kernel_5x5_2[15:8]};
    kernel_img_mul_15[12] <= { {8{1'b0}},layer2_reg_15[23:16]} * { {8{1'b0}}, G_Kernel_5x5_2[23:16]};
    kernel_img_mul_15[13] <= { {8{1'b0}},layer2_reg_15[31:24]} * { {8{1'b0}}, G_Kernel_5x5_2[31:24]};
    kernel_img_mul_15[14] <= { {8{1'b0}},layer2_reg_15[39:32]} * { {8{1'b0}}, G_Kernel_5x5_2[39:32]};
    kernel_img_mul_15[15] <= { {8{1'b0}},layer3_reg_15[7:0]} * { {8{1'b0}}, G_Kernel_5x5_1[7:0]};
    kernel_img_mul_15[16] <= { {8{1'b0}},layer3_reg_15[15:8]} * { {8{1'b0}}, G_Kernel_5x5_1[15:8]};
    kernel_img_mul_15[17] <= { {8{1'b0}},layer3_reg_15[23:16]} * { {8{1'b0}}, G_Kernel_5x5_1[23:16]};
    kernel_img_mul_15[18] <= { {8{1'b0}},layer3_reg_15[31:24]} * { {8{1'b0}}, G_Kernel_5x5_1[31:24]};
    kernel_img_mul_15[19] <= { {8{1'b0}},layer3_reg_15[39:32]} * { {8{1'b0}}, G_Kernel_5x5_1[39:32]};
    kernel_img_mul_15[20] <= { {8{1'b0}},layer4_reg_15[7:0]} * { {8{1'b0}}, G_Kernel_5x5_0[7:0]};
    kernel_img_mul_15[21] <= { {8{1'b0}},layer4_reg_15[15:8]} * { {8{1'b0}}, G_Kernel_5x5_0[15:8]};
    kernel_img_mul_15[22] <= { {8{1'b0}},layer4_reg_15[23:16]} * { {8{1'b0}}, G_Kernel_5x5_0[23:16]};
    kernel_img_mul_15[23] <= { {8{1'b0}},layer4_reg_15[31:24]} * { {8{1'b0}}, G_Kernel_5x5_0[31:24]};
    kernel_img_mul_15[24] <= { {8{1'b0}},layer4_reg_15[39:32]} * { {8{1'b0}}, G_Kernel_5x5_0[39:32]};
  end
end
reg  [15:0]  kernel_img_sum_1_15;
reg  [15:0]  kernel_img_sum_2_15;
reg  [15:0]  kernel_img_sum_3_15;
reg  [15:0]  kernel_img_sum_4_15;
reg  [15:0]  kernel_img_sum_5_15;
reg  [15:0]  kernel_img_sum_6_15;
reg  [15:0]  kernel_img_sum_7_15;
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_1_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_1_15 <= kernel_img_mul_15[0] + kernel_img_mul_15[1] + kernel_img_mul_15[2] + kernel_img_mul_15[3] + kernel_img_mul_15[4];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_2_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_2_15 <= kernel_img_mul_15[5] + kernel_img_mul_15[6] + kernel_img_mul_15[7] + kernel_img_mul_15[8];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_3_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_3_15 <= kernel_img_mul_15[9] + kernel_img_mul_15[10] + kernel_img_mul_15[11] + kernel_img_mul_15[12];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_4_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_4_15 <= kernel_img_mul_15[13] + kernel_img_mul_15[14] + kernel_img_mul_15[15] + kernel_img_mul_15[16];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_5_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_5_15 <= kernel_img_mul_15[17] + kernel_img_mul_15[18] + kernel_img_mul_15[19] + kernel_img_mul_15[20];
  end
end
always@(posedge clk) begin
  if(!rst_n) begin
    kernel_img_sum_6_15 <= 'd0;
  end
  else if(current_state==ST_ADD) begin
    kernel_img_sum_6_15 <= kernel_img_mul_15[21] + kernel_img_mul_15[22] + kernel_img_mul_15[23] + kernel_img_mul_15[24];
  end
end
always@(*) begin
  kernel_img_sum_7_15 = kernel_img_sum_1_15 + kernel_img_sum_2_15 + kernel_img_sum_3_15 + kernel_img_sum_4_15 + kernel_img_sum_5_15 + kernel_img_sum_6_15;
end
always @(posedge clk) begin
  if(!rst_n) begin
    blur_out[7:0] <= 'd0;
    blur_out[15:8] <= 'd0;
    blur_out[23:16] <= 'd0;
    blur_out[31:24] <= 'd0;
    blur_out[39:32] <= 'd0;
    blur_out[47:40] <= 'd0;
    blur_out[55:48] <= 'd0;
    blur_out[63:56] <= 'd0;
    blur_out[71:64] <= 'd0;
    blur_out[79:72] <= 'd0;
    blur_out[87:80] <= 'd0;
    blur_out[95:88] <= 'd0;
    blur_out[103:96] <= 'd0;
    blur_out[111:104] <= 'd0;
    blur_out[119:112] <= 'd0;
    blur_out[127:120] <= 'd0;
  end
  else if(current_state==ST_UPDATE) begin
    blur_out[7:0] <= kernel_img_sum_7_0[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[15:8] <= kernel_img_sum_7_1[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[23:16] <= kernel_img_sum_7_2[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[31:24] <= kernel_img_sum_7_3[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[39:32] <= kernel_img_sum_7_4[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[47:40] <= kernel_img_sum_7_5[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[55:48] <= kernel_img_sum_7_6[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[63:56] <= kernel_img_sum_7_7[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[71:64] <= kernel_img_sum_7_8[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[79:72] <= kernel_img_sum_7_9[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[87:80] <= kernel_img_sum_7_10[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[95:88] <= kernel_img_sum_7_11[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[103:96] <= kernel_img_sum_7_12[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[111:104] <= kernel_img_sum_7_13[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[119:112] <= kernel_img_sum_7_14[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
    blur_out[127:120] <= kernel_img_sum_7_15[15:8];/*Q8.8 -> Q8.0 Q8.32 -> Q8.0*/
  end
end

/*
 *  FSM
 *
 */
always @(posedge clk) begin
  if (!rst_n) begin
    current_state <= ST_MUX;    
  end
  else begin
    current_state <= next_state;
  end
end
always @(*) begin
  case(current_state)
    ST_MUX: begin
      if(start)
        next_state = ST_MUL;
      else
        next_state = ST_MUX;
    end
    ST_MUL: begin
      if(current_state==ST_MUL)
        next_state = ST_ADD;
      else 
        next_state = ST_MUL;
    end
    ST_ADD: begin
      if(current_state==ST_ADD)
        next_state = ST_UPDATE;
      else 
        next_state = ST_ADD;
    end
    ST_UPDATE: begin
      if(current_state==ST_UPDATE)
        next_state = ST_MUX;
      else 
        next_state = ST_UPDATE;
    end
    default:
      next_state = ST_MUX;
  endcase
end

endmodule