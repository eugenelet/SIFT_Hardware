module prepare_filter(
  clk,
  rst_n,
  current_state,
  img_addr,
  filter_input_0_0,
  filter_input_0_1,
  filter_input_0_2,
  filter_input_1_0,
  filter_input_1_1,
  filter_input_1_2,
  buffer_data_2,
  buffer_data_3,
  buffer_data_4,
  buffer_data_5,
  blur3x3_dout,
  blur5x5_1_dout,
  no_keypoint,
  is_keypoint_0,
  is_keypoint_1,
  current_RowCol_0
  current_RowCol_1
);

input      clk,
           rst_n;

input  [2:0]       current_state;
input  [8:0]       img_addr;
input  [5119:0]    buffer_data_2,
                   buffer_data_3,
                   buffer_data_4,
                   buffer_data_5,
                   blur3x3_dout,
                   blur5x5_1_dout;
input  [637:0]     is_keypoint_0;
input  [637:0]     is_keypoint_1;
output [23:0]      filter_input_0_0;
output [23:0]      filter_input_0_1;
output [23:0]      filter_input_0_2;
output [23:0]      filter_input_1_0;
output [23:0]      filter_input_1_1;
output [23:0]      filter_input_1_2;
output [1:0]       no_keypoint;
output [18:0]      current_RowCol_0;
output [18:0]      current_RowCol_1;

/*Module FSM*/
parameter ST_IDLE   = 0,
          ST_READY  = 1,/*Idle 1 state for SRAM to get READY*/
          ST_DETECT = 2,
          ST_FILTER = 3,
          ST_UPDATE = 4,/*Grants a cycle to update MEM addr*/
          ST_BUFFER = 5;/*Grants buffer a cycle to update*/

reg   [637:0] detected_keypoint[0:1];
always @(posedge clk) begin
  if (!rst_n)
    detected_keypoint[0] <= 'd0;
  else if (current_state==ST_DETECT)
    detected_keypoint[0] <= is_keypoint_0;
  else if (current_state==ST_FILTER && detected_keypoint[0][0])
    detected_keypoint[0][0] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][1])
    detected_keypoint[0][1] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][2])
    detected_keypoint[0][2] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][3])
    detected_keypoint[0][3] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][4])
    detected_keypoint[0][4] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][5])
    detected_keypoint[0][5] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][6])
    detected_keypoint[0][6] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][7])
    detected_keypoint[0][7] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][8])
    detected_keypoint[0][8] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][9])
    detected_keypoint[0][9] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][10])
    detected_keypoint[0][10] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][11])
    detected_keypoint[0][11] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][12])
    detected_keypoint[0][12] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][13])
    detected_keypoint[0][13] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][14])
    detected_keypoint[0][14] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][15])
    detected_keypoint[0][15] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][16])
    detected_keypoint[0][16] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][17])
    detected_keypoint[0][17] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][18])
    detected_keypoint[0][18] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][19])
    detected_keypoint[0][19] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][20])
    detected_keypoint[0][20] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][21])
    detected_keypoint[0][21] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][22])
    detected_keypoint[0][22] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][23])
    detected_keypoint[0][23] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][24])
    detected_keypoint[0][24] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][25])
    detected_keypoint[0][25] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][26])
    detected_keypoint[0][26] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][27])
    detected_keypoint[0][27] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][28])
    detected_keypoint[0][28] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][29])
    detected_keypoint[0][29] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][30])
    detected_keypoint[0][30] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][31])
    detected_keypoint[0][31] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][32])
    detected_keypoint[0][32] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][33])
    detected_keypoint[0][33] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][34])
    detected_keypoint[0][34] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][35])
    detected_keypoint[0][35] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][36])
    detected_keypoint[0][36] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][37])
    detected_keypoint[0][37] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][38])
    detected_keypoint[0][38] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][39])
    detected_keypoint[0][39] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][40])
    detected_keypoint[0][40] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][41])
    detected_keypoint[0][41] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][42])
    detected_keypoint[0][42] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][43])
    detected_keypoint[0][43] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][44])
    detected_keypoint[0][44] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][45])
    detected_keypoint[0][45] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][46])
    detected_keypoint[0][46] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][47])
    detected_keypoint[0][47] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][48])
    detected_keypoint[0][48] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][49])
    detected_keypoint[0][49] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][50])
    detected_keypoint[0][50] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][51])
    detected_keypoint[0][51] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][52])
    detected_keypoint[0][52] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][53])
    detected_keypoint[0][53] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][54])
    detected_keypoint[0][54] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][55])
    detected_keypoint[0][55] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][56])
    detected_keypoint[0][56] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][57])
    detected_keypoint[0][57] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][58])
    detected_keypoint[0][58] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][59])
    detected_keypoint[0][59] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][60])
    detected_keypoint[0][60] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][61])
    detected_keypoint[0][61] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][62])
    detected_keypoint[0][62] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][63])
    detected_keypoint[0][63] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][64])
    detected_keypoint[0][64] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][65])
    detected_keypoint[0][65] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][66])
    detected_keypoint[0][66] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][67])
    detected_keypoint[0][67] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][68])
    detected_keypoint[0][68] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][69])
    detected_keypoint[0][69] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][70])
    detected_keypoint[0][70] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][71])
    detected_keypoint[0][71] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][72])
    detected_keypoint[0][72] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][73])
    detected_keypoint[0][73] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][74])
    detected_keypoint[0][74] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][75])
    detected_keypoint[0][75] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][76])
    detected_keypoint[0][76] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][77])
    detected_keypoint[0][77] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][78])
    detected_keypoint[0][78] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][79])
    detected_keypoint[0][79] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][80])
    detected_keypoint[0][80] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][81])
    detected_keypoint[0][81] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][82])
    detected_keypoint[0][82] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][83])
    detected_keypoint[0][83] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][84])
    detected_keypoint[0][84] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][85])
    detected_keypoint[0][85] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][86])
    detected_keypoint[0][86] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][87])
    detected_keypoint[0][87] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][88])
    detected_keypoint[0][88] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][89])
    detected_keypoint[0][89] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][90])
    detected_keypoint[0][90] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][91])
    detected_keypoint[0][91] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][92])
    detected_keypoint[0][92] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][93])
    detected_keypoint[0][93] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][94])
    detected_keypoint[0][94] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][95])
    detected_keypoint[0][95] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][96])
    detected_keypoint[0][96] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][97])
    detected_keypoint[0][97] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][98])
    detected_keypoint[0][98] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][99])
    detected_keypoint[0][99] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][100])
    detected_keypoint[0][100] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][101])
    detected_keypoint[0][101] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][102])
    detected_keypoint[0][102] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][103])
    detected_keypoint[0][103] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][104])
    detected_keypoint[0][104] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][105])
    detected_keypoint[0][105] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][106])
    detected_keypoint[0][106] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][107])
    detected_keypoint[0][107] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][108])
    detected_keypoint[0][108] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][109])
    detected_keypoint[0][109] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][110])
    detected_keypoint[0][110] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][111])
    detected_keypoint[0][111] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][112])
    detected_keypoint[0][112] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][113])
    detected_keypoint[0][113] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][114])
    detected_keypoint[0][114] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][115])
    detected_keypoint[0][115] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][116])
    detected_keypoint[0][116] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][117])
    detected_keypoint[0][117] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][118])
    detected_keypoint[0][118] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][119])
    detected_keypoint[0][119] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][120])
    detected_keypoint[0][120] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][121])
    detected_keypoint[0][121] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][122])
    detected_keypoint[0][122] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][123])
    detected_keypoint[0][123] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][124])
    detected_keypoint[0][124] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][125])
    detected_keypoint[0][125] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][126])
    detected_keypoint[0][126] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][127])
    detected_keypoint[0][127] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][128])
    detected_keypoint[0][128] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][129])
    detected_keypoint[0][129] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][130])
    detected_keypoint[0][130] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][131])
    detected_keypoint[0][131] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][132])
    detected_keypoint[0][132] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][133])
    detected_keypoint[0][133] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][134])
    detected_keypoint[0][134] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][135])
    detected_keypoint[0][135] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][136])
    detected_keypoint[0][136] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][137])
    detected_keypoint[0][137] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][138])
    detected_keypoint[0][138] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][139])
    detected_keypoint[0][139] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][140])
    detected_keypoint[0][140] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][141])
    detected_keypoint[0][141] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][142])
    detected_keypoint[0][142] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][143])
    detected_keypoint[0][143] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][144])
    detected_keypoint[0][144] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][145])
    detected_keypoint[0][145] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][146])
    detected_keypoint[0][146] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][147])
    detected_keypoint[0][147] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][148])
    detected_keypoint[0][148] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][149])
    detected_keypoint[0][149] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][150])
    detected_keypoint[0][150] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][151])
    detected_keypoint[0][151] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][152])
    detected_keypoint[0][152] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][153])
    detected_keypoint[0][153] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][154])
    detected_keypoint[0][154] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][155])
    detected_keypoint[0][155] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][156])
    detected_keypoint[0][156] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][157])
    detected_keypoint[0][157] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][158])
    detected_keypoint[0][158] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][159])
    detected_keypoint[0][159] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][160])
    detected_keypoint[0][160] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][161])
    detected_keypoint[0][161] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][162])
    detected_keypoint[0][162] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][163])
    detected_keypoint[0][163] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][164])
    detected_keypoint[0][164] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][165])
    detected_keypoint[0][165] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][166])
    detected_keypoint[0][166] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][167])
    detected_keypoint[0][167] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][168])
    detected_keypoint[0][168] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][169])
    detected_keypoint[0][169] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][170])
    detected_keypoint[0][170] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][171])
    detected_keypoint[0][171] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][172])
    detected_keypoint[0][172] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][173])
    detected_keypoint[0][173] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][174])
    detected_keypoint[0][174] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][175])
    detected_keypoint[0][175] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][176])
    detected_keypoint[0][176] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][177])
    detected_keypoint[0][177] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][178])
    detected_keypoint[0][178] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][179])
    detected_keypoint[0][179] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][180])
    detected_keypoint[0][180] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][181])
    detected_keypoint[0][181] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][182])
    detected_keypoint[0][182] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][183])
    detected_keypoint[0][183] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][184])
    detected_keypoint[0][184] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][185])
    detected_keypoint[0][185] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][186])
    detected_keypoint[0][186] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][187])
    detected_keypoint[0][187] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][188])
    detected_keypoint[0][188] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][189])
    detected_keypoint[0][189] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][190])
    detected_keypoint[0][190] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][191])
    detected_keypoint[0][191] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][192])
    detected_keypoint[0][192] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][193])
    detected_keypoint[0][193] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][194])
    detected_keypoint[0][194] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][195])
    detected_keypoint[0][195] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][196])
    detected_keypoint[0][196] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][197])
    detected_keypoint[0][197] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][198])
    detected_keypoint[0][198] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][199])
    detected_keypoint[0][199] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][200])
    detected_keypoint[0][200] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][201])
    detected_keypoint[0][201] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][202])
    detected_keypoint[0][202] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][203])
    detected_keypoint[0][203] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][204])
    detected_keypoint[0][204] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][205])
    detected_keypoint[0][205] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][206])
    detected_keypoint[0][206] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][207])
    detected_keypoint[0][207] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][208])
    detected_keypoint[0][208] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][209])
    detected_keypoint[0][209] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][210])
    detected_keypoint[0][210] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][211])
    detected_keypoint[0][211] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][212])
    detected_keypoint[0][212] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][213])
    detected_keypoint[0][213] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][214])
    detected_keypoint[0][214] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][215])
    detected_keypoint[0][215] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][216])
    detected_keypoint[0][216] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][217])
    detected_keypoint[0][217] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][218])
    detected_keypoint[0][218] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][219])
    detected_keypoint[0][219] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][220])
    detected_keypoint[0][220] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][221])
    detected_keypoint[0][221] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][222])
    detected_keypoint[0][222] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][223])
    detected_keypoint[0][223] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][224])
    detected_keypoint[0][224] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][225])
    detected_keypoint[0][225] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][226])
    detected_keypoint[0][226] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][227])
    detected_keypoint[0][227] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][228])
    detected_keypoint[0][228] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][229])
    detected_keypoint[0][229] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][230])
    detected_keypoint[0][230] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][231])
    detected_keypoint[0][231] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][232])
    detected_keypoint[0][232] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][233])
    detected_keypoint[0][233] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][234])
    detected_keypoint[0][234] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][235])
    detected_keypoint[0][235] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][236])
    detected_keypoint[0][236] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][237])
    detected_keypoint[0][237] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][238])
    detected_keypoint[0][238] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][239])
    detected_keypoint[0][239] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][240])
    detected_keypoint[0][240] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][241])
    detected_keypoint[0][241] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][242])
    detected_keypoint[0][242] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][243])
    detected_keypoint[0][243] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][244])
    detected_keypoint[0][244] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][245])
    detected_keypoint[0][245] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][246])
    detected_keypoint[0][246] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][247])
    detected_keypoint[0][247] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][248])
    detected_keypoint[0][248] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][249])
    detected_keypoint[0][249] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][250])
    detected_keypoint[0][250] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][251])
    detected_keypoint[0][251] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][252])
    detected_keypoint[0][252] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][253])
    detected_keypoint[0][253] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][254])
    detected_keypoint[0][254] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][255])
    detected_keypoint[0][255] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][256])
    detected_keypoint[0][256] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][257])
    detected_keypoint[0][257] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][258])
    detected_keypoint[0][258] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][259])
    detected_keypoint[0][259] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][260])
    detected_keypoint[0][260] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][261])
    detected_keypoint[0][261] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][262])
    detected_keypoint[0][262] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][263])
    detected_keypoint[0][263] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][264])
    detected_keypoint[0][264] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][265])
    detected_keypoint[0][265] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][266])
    detected_keypoint[0][266] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][267])
    detected_keypoint[0][267] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][268])
    detected_keypoint[0][268] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][269])
    detected_keypoint[0][269] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][270])
    detected_keypoint[0][270] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][271])
    detected_keypoint[0][271] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][272])
    detected_keypoint[0][272] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][273])
    detected_keypoint[0][273] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][274])
    detected_keypoint[0][274] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][275])
    detected_keypoint[0][275] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][276])
    detected_keypoint[0][276] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][277])
    detected_keypoint[0][277] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][278])
    detected_keypoint[0][278] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][279])
    detected_keypoint[0][279] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][280])
    detected_keypoint[0][280] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][281])
    detected_keypoint[0][281] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][282])
    detected_keypoint[0][282] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][283])
    detected_keypoint[0][283] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][284])
    detected_keypoint[0][284] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][285])
    detected_keypoint[0][285] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][286])
    detected_keypoint[0][286] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][287])
    detected_keypoint[0][287] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][288])
    detected_keypoint[0][288] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][289])
    detected_keypoint[0][289] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][290])
    detected_keypoint[0][290] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][291])
    detected_keypoint[0][291] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][292])
    detected_keypoint[0][292] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][293])
    detected_keypoint[0][293] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][294])
    detected_keypoint[0][294] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][295])
    detected_keypoint[0][295] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][296])
    detected_keypoint[0][296] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][297])
    detected_keypoint[0][297] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][298])
    detected_keypoint[0][298] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][299])
    detected_keypoint[0][299] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][300])
    detected_keypoint[0][300] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][301])
    detected_keypoint[0][301] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][302])
    detected_keypoint[0][302] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][303])
    detected_keypoint[0][303] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][304])
    detected_keypoint[0][304] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][305])
    detected_keypoint[0][305] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][306])
    detected_keypoint[0][306] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][307])
    detected_keypoint[0][307] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][308])
    detected_keypoint[0][308] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][309])
    detected_keypoint[0][309] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][310])
    detected_keypoint[0][310] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][311])
    detected_keypoint[0][311] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][312])
    detected_keypoint[0][312] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][313])
    detected_keypoint[0][313] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][314])
    detected_keypoint[0][314] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][315])
    detected_keypoint[0][315] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][316])
    detected_keypoint[0][316] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][317])
    detected_keypoint[0][317] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][318])
    detected_keypoint[0][318] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][319])
    detected_keypoint[0][319] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][320])
    detected_keypoint[0][320] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][321])
    detected_keypoint[0][321] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][322])
    detected_keypoint[0][322] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][323])
    detected_keypoint[0][323] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][324])
    detected_keypoint[0][324] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][325])
    detected_keypoint[0][325] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][326])
    detected_keypoint[0][326] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][327])
    detected_keypoint[0][327] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][328])
    detected_keypoint[0][328] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][329])
    detected_keypoint[0][329] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][330])
    detected_keypoint[0][330] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][331])
    detected_keypoint[0][331] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][332])
    detected_keypoint[0][332] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][333])
    detected_keypoint[0][333] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][334])
    detected_keypoint[0][334] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][335])
    detected_keypoint[0][335] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][336])
    detected_keypoint[0][336] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][337])
    detected_keypoint[0][337] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][338])
    detected_keypoint[0][338] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][339])
    detected_keypoint[0][339] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][340])
    detected_keypoint[0][340] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][341])
    detected_keypoint[0][341] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][342])
    detected_keypoint[0][342] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][343])
    detected_keypoint[0][343] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][344])
    detected_keypoint[0][344] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][345])
    detected_keypoint[0][345] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][346])
    detected_keypoint[0][346] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][347])
    detected_keypoint[0][347] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][348])
    detected_keypoint[0][348] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][349])
    detected_keypoint[0][349] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][350])
    detected_keypoint[0][350] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][351])
    detected_keypoint[0][351] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][352])
    detected_keypoint[0][352] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][353])
    detected_keypoint[0][353] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][354])
    detected_keypoint[0][354] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][355])
    detected_keypoint[0][355] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][356])
    detected_keypoint[0][356] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][357])
    detected_keypoint[0][357] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][358])
    detected_keypoint[0][358] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][359])
    detected_keypoint[0][359] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][360])
    detected_keypoint[0][360] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][361])
    detected_keypoint[0][361] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][362])
    detected_keypoint[0][362] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][363])
    detected_keypoint[0][363] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][364])
    detected_keypoint[0][364] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][365])
    detected_keypoint[0][365] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][366])
    detected_keypoint[0][366] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][367])
    detected_keypoint[0][367] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][368])
    detected_keypoint[0][368] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][369])
    detected_keypoint[0][369] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][370])
    detected_keypoint[0][370] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][371])
    detected_keypoint[0][371] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][372])
    detected_keypoint[0][372] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][373])
    detected_keypoint[0][373] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][374])
    detected_keypoint[0][374] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][375])
    detected_keypoint[0][375] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][376])
    detected_keypoint[0][376] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][377])
    detected_keypoint[0][377] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][378])
    detected_keypoint[0][378] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][379])
    detected_keypoint[0][379] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][380])
    detected_keypoint[0][380] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][381])
    detected_keypoint[0][381] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][382])
    detected_keypoint[0][382] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][383])
    detected_keypoint[0][383] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][384])
    detected_keypoint[0][384] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][385])
    detected_keypoint[0][385] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][386])
    detected_keypoint[0][386] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][387])
    detected_keypoint[0][387] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][388])
    detected_keypoint[0][388] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][389])
    detected_keypoint[0][389] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][390])
    detected_keypoint[0][390] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][391])
    detected_keypoint[0][391] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][392])
    detected_keypoint[0][392] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][393])
    detected_keypoint[0][393] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][394])
    detected_keypoint[0][394] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][395])
    detected_keypoint[0][395] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][396])
    detected_keypoint[0][396] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][397])
    detected_keypoint[0][397] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][398])
    detected_keypoint[0][398] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][399])
    detected_keypoint[0][399] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][400])
    detected_keypoint[0][400] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][401])
    detected_keypoint[0][401] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][402])
    detected_keypoint[0][402] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][403])
    detected_keypoint[0][403] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][404])
    detected_keypoint[0][404] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][405])
    detected_keypoint[0][405] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][406])
    detected_keypoint[0][406] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][407])
    detected_keypoint[0][407] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][408])
    detected_keypoint[0][408] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][409])
    detected_keypoint[0][409] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][410])
    detected_keypoint[0][410] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][411])
    detected_keypoint[0][411] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][412])
    detected_keypoint[0][412] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][413])
    detected_keypoint[0][413] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][414])
    detected_keypoint[0][414] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][415])
    detected_keypoint[0][415] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][416])
    detected_keypoint[0][416] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][417])
    detected_keypoint[0][417] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][418])
    detected_keypoint[0][418] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][419])
    detected_keypoint[0][419] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][420])
    detected_keypoint[0][420] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][421])
    detected_keypoint[0][421] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][422])
    detected_keypoint[0][422] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][423])
    detected_keypoint[0][423] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][424])
    detected_keypoint[0][424] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][425])
    detected_keypoint[0][425] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][426])
    detected_keypoint[0][426] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][427])
    detected_keypoint[0][427] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][428])
    detected_keypoint[0][428] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][429])
    detected_keypoint[0][429] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][430])
    detected_keypoint[0][430] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][431])
    detected_keypoint[0][431] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][432])
    detected_keypoint[0][432] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][433])
    detected_keypoint[0][433] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][434])
    detected_keypoint[0][434] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][435])
    detected_keypoint[0][435] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][436])
    detected_keypoint[0][436] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][437])
    detected_keypoint[0][437] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][438])
    detected_keypoint[0][438] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][439])
    detected_keypoint[0][439] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][440])
    detected_keypoint[0][440] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][441])
    detected_keypoint[0][441] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][442])
    detected_keypoint[0][442] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][443])
    detected_keypoint[0][443] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][444])
    detected_keypoint[0][444] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][445])
    detected_keypoint[0][445] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][446])
    detected_keypoint[0][446] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][447])
    detected_keypoint[0][447] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][448])
    detected_keypoint[0][448] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][449])
    detected_keypoint[0][449] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][450])
    detected_keypoint[0][450] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][451])
    detected_keypoint[0][451] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][452])
    detected_keypoint[0][452] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][453])
    detected_keypoint[0][453] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][454])
    detected_keypoint[0][454] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][455])
    detected_keypoint[0][455] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][456])
    detected_keypoint[0][456] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][457])
    detected_keypoint[0][457] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][458])
    detected_keypoint[0][458] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][459])
    detected_keypoint[0][459] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][460])
    detected_keypoint[0][460] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][461])
    detected_keypoint[0][461] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][462])
    detected_keypoint[0][462] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][463])
    detected_keypoint[0][463] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][464])
    detected_keypoint[0][464] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][465])
    detected_keypoint[0][465] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][466])
    detected_keypoint[0][466] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][467])
    detected_keypoint[0][467] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][468])
    detected_keypoint[0][468] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][469])
    detected_keypoint[0][469] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][470])
    detected_keypoint[0][470] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][471])
    detected_keypoint[0][471] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][472])
    detected_keypoint[0][472] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][473])
    detected_keypoint[0][473] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][474])
    detected_keypoint[0][474] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][475])
    detected_keypoint[0][475] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][476])
    detected_keypoint[0][476] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][477])
    detected_keypoint[0][477] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][478])
    detected_keypoint[0][478] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][479])
    detected_keypoint[0][479] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][480])
    detected_keypoint[0][480] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][481])
    detected_keypoint[0][481] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][482])
    detected_keypoint[0][482] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][483])
    detected_keypoint[0][483] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][484])
    detected_keypoint[0][484] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][485])
    detected_keypoint[0][485] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][486])
    detected_keypoint[0][486] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][487])
    detected_keypoint[0][487] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][488])
    detected_keypoint[0][488] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][489])
    detected_keypoint[0][489] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][490])
    detected_keypoint[0][490] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][491])
    detected_keypoint[0][491] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][492])
    detected_keypoint[0][492] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][493])
    detected_keypoint[0][493] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][494])
    detected_keypoint[0][494] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][495])
    detected_keypoint[0][495] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][496])
    detected_keypoint[0][496] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][497])
    detected_keypoint[0][497] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][498])
    detected_keypoint[0][498] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][499])
    detected_keypoint[0][499] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][500])
    detected_keypoint[0][500] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][501])
    detected_keypoint[0][501] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][502])
    detected_keypoint[0][502] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][503])
    detected_keypoint[0][503] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][504])
    detected_keypoint[0][504] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][505])
    detected_keypoint[0][505] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][506])
    detected_keypoint[0][506] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][507])
    detected_keypoint[0][507] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][508])
    detected_keypoint[0][508] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][509])
    detected_keypoint[0][509] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][510])
    detected_keypoint[0][510] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][511])
    detected_keypoint[0][511] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][512])
    detected_keypoint[0][512] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][513])
    detected_keypoint[0][513] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][514])
    detected_keypoint[0][514] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][515])
    detected_keypoint[0][515] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][516])
    detected_keypoint[0][516] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][517])
    detected_keypoint[0][517] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][518])
    detected_keypoint[0][518] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][519])
    detected_keypoint[0][519] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][520])
    detected_keypoint[0][520] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][521])
    detected_keypoint[0][521] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][522])
    detected_keypoint[0][522] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][523])
    detected_keypoint[0][523] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][524])
    detected_keypoint[0][524] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][525])
    detected_keypoint[0][525] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][526])
    detected_keypoint[0][526] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][527])
    detected_keypoint[0][527] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][528])
    detected_keypoint[0][528] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][529])
    detected_keypoint[0][529] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][530])
    detected_keypoint[0][530] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][531])
    detected_keypoint[0][531] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][532])
    detected_keypoint[0][532] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][533])
    detected_keypoint[0][533] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][534])
    detected_keypoint[0][534] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][535])
    detected_keypoint[0][535] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][536])
    detected_keypoint[0][536] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][537])
    detected_keypoint[0][537] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][538])
    detected_keypoint[0][538] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][539])
    detected_keypoint[0][539] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][540])
    detected_keypoint[0][540] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][541])
    detected_keypoint[0][541] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][542])
    detected_keypoint[0][542] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][543])
    detected_keypoint[0][543] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][544])
    detected_keypoint[0][544] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][545])
    detected_keypoint[0][545] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][546])
    detected_keypoint[0][546] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][547])
    detected_keypoint[0][547] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][548])
    detected_keypoint[0][548] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][549])
    detected_keypoint[0][549] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][550])
    detected_keypoint[0][550] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][551])
    detected_keypoint[0][551] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][552])
    detected_keypoint[0][552] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][553])
    detected_keypoint[0][553] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][554])
    detected_keypoint[0][554] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][555])
    detected_keypoint[0][555] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][556])
    detected_keypoint[0][556] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][557])
    detected_keypoint[0][557] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][558])
    detected_keypoint[0][558] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][559])
    detected_keypoint[0][559] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][560])
    detected_keypoint[0][560] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][561])
    detected_keypoint[0][561] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][562])
    detected_keypoint[0][562] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][563])
    detected_keypoint[0][563] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][564])
    detected_keypoint[0][564] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][565])
    detected_keypoint[0][565] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][566])
    detected_keypoint[0][566] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][567])
    detected_keypoint[0][567] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][568])
    detected_keypoint[0][568] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][569])
    detected_keypoint[0][569] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][570])
    detected_keypoint[0][570] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][571])
    detected_keypoint[0][571] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][572])
    detected_keypoint[0][572] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][573])
    detected_keypoint[0][573] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][574])
    detected_keypoint[0][574] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][575])
    detected_keypoint[0][575] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][576])
    detected_keypoint[0][576] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][577])
    detected_keypoint[0][577] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][578])
    detected_keypoint[0][578] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][579])
    detected_keypoint[0][579] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][580])
    detected_keypoint[0][580] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][581])
    detected_keypoint[0][581] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][582])
    detected_keypoint[0][582] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][583])
    detected_keypoint[0][583] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][584])
    detected_keypoint[0][584] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][585])
    detected_keypoint[0][585] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][586])
    detected_keypoint[0][586] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][587])
    detected_keypoint[0][587] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][588])
    detected_keypoint[0][588] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][589])
    detected_keypoint[0][589] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][590])
    detected_keypoint[0][590] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][591])
    detected_keypoint[0][591] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][592])
    detected_keypoint[0][592] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][593])
    detected_keypoint[0][593] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][594])
    detected_keypoint[0][594] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][595])
    detected_keypoint[0][595] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][596])
    detected_keypoint[0][596] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][597])
    detected_keypoint[0][597] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][598])
    detected_keypoint[0][598] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][599])
    detected_keypoint[0][599] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][600])
    detected_keypoint[0][600] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][601])
    detected_keypoint[0][601] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][602])
    detected_keypoint[0][602] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][603])
    detected_keypoint[0][603] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][604])
    detected_keypoint[0][604] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][605])
    detected_keypoint[0][605] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][606])
    detected_keypoint[0][606] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][607])
    detected_keypoint[0][607] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][608])
    detected_keypoint[0][608] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][609])
    detected_keypoint[0][609] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][610])
    detected_keypoint[0][610] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][611])
    detected_keypoint[0][611] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][612])
    detected_keypoint[0][612] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][613])
    detected_keypoint[0][613] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][614])
    detected_keypoint[0][614] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][615])
    detected_keypoint[0][615] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][616])
    detected_keypoint[0][616] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][617])
    detected_keypoint[0][617] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][618])
    detected_keypoint[0][618] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][619])
    detected_keypoint[0][619] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][620])
    detected_keypoint[0][620] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][621])
    detected_keypoint[0][621] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][622])
    detected_keypoint[0][622] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][623])
    detected_keypoint[0][623] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][624])
    detected_keypoint[0][624] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][625])
    detected_keypoint[0][625] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][626])
    detected_keypoint[0][626] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][627])
    detected_keypoint[0][627] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][628])
    detected_keypoint[0][628] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][629])
    detected_keypoint[0][629] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][630])
    detected_keypoint[0][630] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][631])
    detected_keypoint[0][631] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][632])
    detected_keypoint[0][632] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][633])
    detected_keypoint[0][633] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][634])
    detected_keypoint[0][634] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][635])
    detected_keypoint[0][635] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][636])
    detected_keypoint[0][636] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[0][637])
    detected_keypoint[0][637] <= 1'b0;
  else
    detected_keypoint[0] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    detected_keypoint[1] <= 'd0;
  else if (current_state==ST_DETECT)
    detected_keypoint[1] <= is_keypoint_1;
  else if (current_state==ST_FILTER && detected_keypoint[1][0])
    detected_keypoint[1][0] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][1])
    detected_keypoint[1][1] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][2])
    detected_keypoint[1][2] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][3])
    detected_keypoint[1][3] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][4])
    detected_keypoint[1][4] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][5])
    detected_keypoint[1][5] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][6])
    detected_keypoint[1][6] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][7])
    detected_keypoint[1][7] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][8])
    detected_keypoint[1][8] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][9])
    detected_keypoint[1][9] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][10])
    detected_keypoint[1][10] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][11])
    detected_keypoint[1][11] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][12])
    detected_keypoint[1][12] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][13])
    detected_keypoint[1][13] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][14])
    detected_keypoint[1][14] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][15])
    detected_keypoint[1][15] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][16])
    detected_keypoint[1][16] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][17])
    detected_keypoint[1][17] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][18])
    detected_keypoint[1][18] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][19])
    detected_keypoint[1][19] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][20])
    detected_keypoint[1][20] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][21])
    detected_keypoint[1][21] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][22])
    detected_keypoint[1][22] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][23])
    detected_keypoint[1][23] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][24])
    detected_keypoint[1][24] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][25])
    detected_keypoint[1][25] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][26])
    detected_keypoint[1][26] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][27])
    detected_keypoint[1][27] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][28])
    detected_keypoint[1][28] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][29])
    detected_keypoint[1][29] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][30])
    detected_keypoint[1][30] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][31])
    detected_keypoint[1][31] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][32])
    detected_keypoint[1][32] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][33])
    detected_keypoint[1][33] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][34])
    detected_keypoint[1][34] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][35])
    detected_keypoint[1][35] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][36])
    detected_keypoint[1][36] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][37])
    detected_keypoint[1][37] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][38])
    detected_keypoint[1][38] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][39])
    detected_keypoint[1][39] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][40])
    detected_keypoint[1][40] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][41])
    detected_keypoint[1][41] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][42])
    detected_keypoint[1][42] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][43])
    detected_keypoint[1][43] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][44])
    detected_keypoint[1][44] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][45])
    detected_keypoint[1][45] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][46])
    detected_keypoint[1][46] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][47])
    detected_keypoint[1][47] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][48])
    detected_keypoint[1][48] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][49])
    detected_keypoint[1][49] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][50])
    detected_keypoint[1][50] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][51])
    detected_keypoint[1][51] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][52])
    detected_keypoint[1][52] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][53])
    detected_keypoint[1][53] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][54])
    detected_keypoint[1][54] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][55])
    detected_keypoint[1][55] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][56])
    detected_keypoint[1][56] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][57])
    detected_keypoint[1][57] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][58])
    detected_keypoint[1][58] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][59])
    detected_keypoint[1][59] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][60])
    detected_keypoint[1][60] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][61])
    detected_keypoint[1][61] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][62])
    detected_keypoint[1][62] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][63])
    detected_keypoint[1][63] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][64])
    detected_keypoint[1][64] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][65])
    detected_keypoint[1][65] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][66])
    detected_keypoint[1][66] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][67])
    detected_keypoint[1][67] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][68])
    detected_keypoint[1][68] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][69])
    detected_keypoint[1][69] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][70])
    detected_keypoint[1][70] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][71])
    detected_keypoint[1][71] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][72])
    detected_keypoint[1][72] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][73])
    detected_keypoint[1][73] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][74])
    detected_keypoint[1][74] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][75])
    detected_keypoint[1][75] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][76])
    detected_keypoint[1][76] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][77])
    detected_keypoint[1][77] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][78])
    detected_keypoint[1][78] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][79])
    detected_keypoint[1][79] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][80])
    detected_keypoint[1][80] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][81])
    detected_keypoint[1][81] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][82])
    detected_keypoint[1][82] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][83])
    detected_keypoint[1][83] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][84])
    detected_keypoint[1][84] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][85])
    detected_keypoint[1][85] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][86])
    detected_keypoint[1][86] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][87])
    detected_keypoint[1][87] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][88])
    detected_keypoint[1][88] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][89])
    detected_keypoint[1][89] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][90])
    detected_keypoint[1][90] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][91])
    detected_keypoint[1][91] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][92])
    detected_keypoint[1][92] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][93])
    detected_keypoint[1][93] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][94])
    detected_keypoint[1][94] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][95])
    detected_keypoint[1][95] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][96])
    detected_keypoint[1][96] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][97])
    detected_keypoint[1][97] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][98])
    detected_keypoint[1][98] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][99])
    detected_keypoint[1][99] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][100])
    detected_keypoint[1][100] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][101])
    detected_keypoint[1][101] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][102])
    detected_keypoint[1][102] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][103])
    detected_keypoint[1][103] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][104])
    detected_keypoint[1][104] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][105])
    detected_keypoint[1][105] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][106])
    detected_keypoint[1][106] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][107])
    detected_keypoint[1][107] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][108])
    detected_keypoint[1][108] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][109])
    detected_keypoint[1][109] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][110])
    detected_keypoint[1][110] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][111])
    detected_keypoint[1][111] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][112])
    detected_keypoint[1][112] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][113])
    detected_keypoint[1][113] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][114])
    detected_keypoint[1][114] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][115])
    detected_keypoint[1][115] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][116])
    detected_keypoint[1][116] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][117])
    detected_keypoint[1][117] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][118])
    detected_keypoint[1][118] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][119])
    detected_keypoint[1][119] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][120])
    detected_keypoint[1][120] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][121])
    detected_keypoint[1][121] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][122])
    detected_keypoint[1][122] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][123])
    detected_keypoint[1][123] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][124])
    detected_keypoint[1][124] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][125])
    detected_keypoint[1][125] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][126])
    detected_keypoint[1][126] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][127])
    detected_keypoint[1][127] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][128])
    detected_keypoint[1][128] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][129])
    detected_keypoint[1][129] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][130])
    detected_keypoint[1][130] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][131])
    detected_keypoint[1][131] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][132])
    detected_keypoint[1][132] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][133])
    detected_keypoint[1][133] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][134])
    detected_keypoint[1][134] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][135])
    detected_keypoint[1][135] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][136])
    detected_keypoint[1][136] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][137])
    detected_keypoint[1][137] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][138])
    detected_keypoint[1][138] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][139])
    detected_keypoint[1][139] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][140])
    detected_keypoint[1][140] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][141])
    detected_keypoint[1][141] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][142])
    detected_keypoint[1][142] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][143])
    detected_keypoint[1][143] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][144])
    detected_keypoint[1][144] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][145])
    detected_keypoint[1][145] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][146])
    detected_keypoint[1][146] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][147])
    detected_keypoint[1][147] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][148])
    detected_keypoint[1][148] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][149])
    detected_keypoint[1][149] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][150])
    detected_keypoint[1][150] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][151])
    detected_keypoint[1][151] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][152])
    detected_keypoint[1][152] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][153])
    detected_keypoint[1][153] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][154])
    detected_keypoint[1][154] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][155])
    detected_keypoint[1][155] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][156])
    detected_keypoint[1][156] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][157])
    detected_keypoint[1][157] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][158])
    detected_keypoint[1][158] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][159])
    detected_keypoint[1][159] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][160])
    detected_keypoint[1][160] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][161])
    detected_keypoint[1][161] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][162])
    detected_keypoint[1][162] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][163])
    detected_keypoint[1][163] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][164])
    detected_keypoint[1][164] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][165])
    detected_keypoint[1][165] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][166])
    detected_keypoint[1][166] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][167])
    detected_keypoint[1][167] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][168])
    detected_keypoint[1][168] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][169])
    detected_keypoint[1][169] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][170])
    detected_keypoint[1][170] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][171])
    detected_keypoint[1][171] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][172])
    detected_keypoint[1][172] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][173])
    detected_keypoint[1][173] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][174])
    detected_keypoint[1][174] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][175])
    detected_keypoint[1][175] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][176])
    detected_keypoint[1][176] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][177])
    detected_keypoint[1][177] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][178])
    detected_keypoint[1][178] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][179])
    detected_keypoint[1][179] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][180])
    detected_keypoint[1][180] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][181])
    detected_keypoint[1][181] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][182])
    detected_keypoint[1][182] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][183])
    detected_keypoint[1][183] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][184])
    detected_keypoint[1][184] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][185])
    detected_keypoint[1][185] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][186])
    detected_keypoint[1][186] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][187])
    detected_keypoint[1][187] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][188])
    detected_keypoint[1][188] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][189])
    detected_keypoint[1][189] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][190])
    detected_keypoint[1][190] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][191])
    detected_keypoint[1][191] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][192])
    detected_keypoint[1][192] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][193])
    detected_keypoint[1][193] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][194])
    detected_keypoint[1][194] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][195])
    detected_keypoint[1][195] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][196])
    detected_keypoint[1][196] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][197])
    detected_keypoint[1][197] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][198])
    detected_keypoint[1][198] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][199])
    detected_keypoint[1][199] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][200])
    detected_keypoint[1][200] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][201])
    detected_keypoint[1][201] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][202])
    detected_keypoint[1][202] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][203])
    detected_keypoint[1][203] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][204])
    detected_keypoint[1][204] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][205])
    detected_keypoint[1][205] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][206])
    detected_keypoint[1][206] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][207])
    detected_keypoint[1][207] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][208])
    detected_keypoint[1][208] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][209])
    detected_keypoint[1][209] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][210])
    detected_keypoint[1][210] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][211])
    detected_keypoint[1][211] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][212])
    detected_keypoint[1][212] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][213])
    detected_keypoint[1][213] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][214])
    detected_keypoint[1][214] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][215])
    detected_keypoint[1][215] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][216])
    detected_keypoint[1][216] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][217])
    detected_keypoint[1][217] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][218])
    detected_keypoint[1][218] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][219])
    detected_keypoint[1][219] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][220])
    detected_keypoint[1][220] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][221])
    detected_keypoint[1][221] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][222])
    detected_keypoint[1][222] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][223])
    detected_keypoint[1][223] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][224])
    detected_keypoint[1][224] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][225])
    detected_keypoint[1][225] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][226])
    detected_keypoint[1][226] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][227])
    detected_keypoint[1][227] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][228])
    detected_keypoint[1][228] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][229])
    detected_keypoint[1][229] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][230])
    detected_keypoint[1][230] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][231])
    detected_keypoint[1][231] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][232])
    detected_keypoint[1][232] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][233])
    detected_keypoint[1][233] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][234])
    detected_keypoint[1][234] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][235])
    detected_keypoint[1][235] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][236])
    detected_keypoint[1][236] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][237])
    detected_keypoint[1][237] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][238])
    detected_keypoint[1][238] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][239])
    detected_keypoint[1][239] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][240])
    detected_keypoint[1][240] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][241])
    detected_keypoint[1][241] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][242])
    detected_keypoint[1][242] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][243])
    detected_keypoint[1][243] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][244])
    detected_keypoint[1][244] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][245])
    detected_keypoint[1][245] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][246])
    detected_keypoint[1][246] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][247])
    detected_keypoint[1][247] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][248])
    detected_keypoint[1][248] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][249])
    detected_keypoint[1][249] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][250])
    detected_keypoint[1][250] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][251])
    detected_keypoint[1][251] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][252])
    detected_keypoint[1][252] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][253])
    detected_keypoint[1][253] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][254])
    detected_keypoint[1][254] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][255])
    detected_keypoint[1][255] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][256])
    detected_keypoint[1][256] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][257])
    detected_keypoint[1][257] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][258])
    detected_keypoint[1][258] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][259])
    detected_keypoint[1][259] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][260])
    detected_keypoint[1][260] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][261])
    detected_keypoint[1][261] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][262])
    detected_keypoint[1][262] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][263])
    detected_keypoint[1][263] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][264])
    detected_keypoint[1][264] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][265])
    detected_keypoint[1][265] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][266])
    detected_keypoint[1][266] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][267])
    detected_keypoint[1][267] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][268])
    detected_keypoint[1][268] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][269])
    detected_keypoint[1][269] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][270])
    detected_keypoint[1][270] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][271])
    detected_keypoint[1][271] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][272])
    detected_keypoint[1][272] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][273])
    detected_keypoint[1][273] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][274])
    detected_keypoint[1][274] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][275])
    detected_keypoint[1][275] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][276])
    detected_keypoint[1][276] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][277])
    detected_keypoint[1][277] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][278])
    detected_keypoint[1][278] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][279])
    detected_keypoint[1][279] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][280])
    detected_keypoint[1][280] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][281])
    detected_keypoint[1][281] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][282])
    detected_keypoint[1][282] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][283])
    detected_keypoint[1][283] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][284])
    detected_keypoint[1][284] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][285])
    detected_keypoint[1][285] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][286])
    detected_keypoint[1][286] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][287])
    detected_keypoint[1][287] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][288])
    detected_keypoint[1][288] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][289])
    detected_keypoint[1][289] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][290])
    detected_keypoint[1][290] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][291])
    detected_keypoint[1][291] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][292])
    detected_keypoint[1][292] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][293])
    detected_keypoint[1][293] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][294])
    detected_keypoint[1][294] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][295])
    detected_keypoint[1][295] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][296])
    detected_keypoint[1][296] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][297])
    detected_keypoint[1][297] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][298])
    detected_keypoint[1][298] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][299])
    detected_keypoint[1][299] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][300])
    detected_keypoint[1][300] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][301])
    detected_keypoint[1][301] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][302])
    detected_keypoint[1][302] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][303])
    detected_keypoint[1][303] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][304])
    detected_keypoint[1][304] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][305])
    detected_keypoint[1][305] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][306])
    detected_keypoint[1][306] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][307])
    detected_keypoint[1][307] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][308])
    detected_keypoint[1][308] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][309])
    detected_keypoint[1][309] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][310])
    detected_keypoint[1][310] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][311])
    detected_keypoint[1][311] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][312])
    detected_keypoint[1][312] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][313])
    detected_keypoint[1][313] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][314])
    detected_keypoint[1][314] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][315])
    detected_keypoint[1][315] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][316])
    detected_keypoint[1][316] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][317])
    detected_keypoint[1][317] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][318])
    detected_keypoint[1][318] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][319])
    detected_keypoint[1][319] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][320])
    detected_keypoint[1][320] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][321])
    detected_keypoint[1][321] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][322])
    detected_keypoint[1][322] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][323])
    detected_keypoint[1][323] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][324])
    detected_keypoint[1][324] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][325])
    detected_keypoint[1][325] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][326])
    detected_keypoint[1][326] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][327])
    detected_keypoint[1][327] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][328])
    detected_keypoint[1][328] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][329])
    detected_keypoint[1][329] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][330])
    detected_keypoint[1][330] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][331])
    detected_keypoint[1][331] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][332])
    detected_keypoint[1][332] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][333])
    detected_keypoint[1][333] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][334])
    detected_keypoint[1][334] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][335])
    detected_keypoint[1][335] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][336])
    detected_keypoint[1][336] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][337])
    detected_keypoint[1][337] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][338])
    detected_keypoint[1][338] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][339])
    detected_keypoint[1][339] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][340])
    detected_keypoint[1][340] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][341])
    detected_keypoint[1][341] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][342])
    detected_keypoint[1][342] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][343])
    detected_keypoint[1][343] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][344])
    detected_keypoint[1][344] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][345])
    detected_keypoint[1][345] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][346])
    detected_keypoint[1][346] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][347])
    detected_keypoint[1][347] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][348])
    detected_keypoint[1][348] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][349])
    detected_keypoint[1][349] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][350])
    detected_keypoint[1][350] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][351])
    detected_keypoint[1][351] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][352])
    detected_keypoint[1][352] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][353])
    detected_keypoint[1][353] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][354])
    detected_keypoint[1][354] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][355])
    detected_keypoint[1][355] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][356])
    detected_keypoint[1][356] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][357])
    detected_keypoint[1][357] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][358])
    detected_keypoint[1][358] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][359])
    detected_keypoint[1][359] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][360])
    detected_keypoint[1][360] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][361])
    detected_keypoint[1][361] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][362])
    detected_keypoint[1][362] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][363])
    detected_keypoint[1][363] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][364])
    detected_keypoint[1][364] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][365])
    detected_keypoint[1][365] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][366])
    detected_keypoint[1][366] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][367])
    detected_keypoint[1][367] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][368])
    detected_keypoint[1][368] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][369])
    detected_keypoint[1][369] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][370])
    detected_keypoint[1][370] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][371])
    detected_keypoint[1][371] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][372])
    detected_keypoint[1][372] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][373])
    detected_keypoint[1][373] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][374])
    detected_keypoint[1][374] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][375])
    detected_keypoint[1][375] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][376])
    detected_keypoint[1][376] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][377])
    detected_keypoint[1][377] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][378])
    detected_keypoint[1][378] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][379])
    detected_keypoint[1][379] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][380])
    detected_keypoint[1][380] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][381])
    detected_keypoint[1][381] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][382])
    detected_keypoint[1][382] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][383])
    detected_keypoint[1][383] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][384])
    detected_keypoint[1][384] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][385])
    detected_keypoint[1][385] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][386])
    detected_keypoint[1][386] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][387])
    detected_keypoint[1][387] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][388])
    detected_keypoint[1][388] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][389])
    detected_keypoint[1][389] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][390])
    detected_keypoint[1][390] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][391])
    detected_keypoint[1][391] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][392])
    detected_keypoint[1][392] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][393])
    detected_keypoint[1][393] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][394])
    detected_keypoint[1][394] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][395])
    detected_keypoint[1][395] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][396])
    detected_keypoint[1][396] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][397])
    detected_keypoint[1][397] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][398])
    detected_keypoint[1][398] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][399])
    detected_keypoint[1][399] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][400])
    detected_keypoint[1][400] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][401])
    detected_keypoint[1][401] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][402])
    detected_keypoint[1][402] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][403])
    detected_keypoint[1][403] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][404])
    detected_keypoint[1][404] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][405])
    detected_keypoint[1][405] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][406])
    detected_keypoint[1][406] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][407])
    detected_keypoint[1][407] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][408])
    detected_keypoint[1][408] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][409])
    detected_keypoint[1][409] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][410])
    detected_keypoint[1][410] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][411])
    detected_keypoint[1][411] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][412])
    detected_keypoint[1][412] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][413])
    detected_keypoint[1][413] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][414])
    detected_keypoint[1][414] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][415])
    detected_keypoint[1][415] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][416])
    detected_keypoint[1][416] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][417])
    detected_keypoint[1][417] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][418])
    detected_keypoint[1][418] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][419])
    detected_keypoint[1][419] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][420])
    detected_keypoint[1][420] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][421])
    detected_keypoint[1][421] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][422])
    detected_keypoint[1][422] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][423])
    detected_keypoint[1][423] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][424])
    detected_keypoint[1][424] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][425])
    detected_keypoint[1][425] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][426])
    detected_keypoint[1][426] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][427])
    detected_keypoint[1][427] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][428])
    detected_keypoint[1][428] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][429])
    detected_keypoint[1][429] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][430])
    detected_keypoint[1][430] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][431])
    detected_keypoint[1][431] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][432])
    detected_keypoint[1][432] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][433])
    detected_keypoint[1][433] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][434])
    detected_keypoint[1][434] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][435])
    detected_keypoint[1][435] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][436])
    detected_keypoint[1][436] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][437])
    detected_keypoint[1][437] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][438])
    detected_keypoint[1][438] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][439])
    detected_keypoint[1][439] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][440])
    detected_keypoint[1][440] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][441])
    detected_keypoint[1][441] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][442])
    detected_keypoint[1][442] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][443])
    detected_keypoint[1][443] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][444])
    detected_keypoint[1][444] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][445])
    detected_keypoint[1][445] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][446])
    detected_keypoint[1][446] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][447])
    detected_keypoint[1][447] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][448])
    detected_keypoint[1][448] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][449])
    detected_keypoint[1][449] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][450])
    detected_keypoint[1][450] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][451])
    detected_keypoint[1][451] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][452])
    detected_keypoint[1][452] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][453])
    detected_keypoint[1][453] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][454])
    detected_keypoint[1][454] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][455])
    detected_keypoint[1][455] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][456])
    detected_keypoint[1][456] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][457])
    detected_keypoint[1][457] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][458])
    detected_keypoint[1][458] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][459])
    detected_keypoint[1][459] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][460])
    detected_keypoint[1][460] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][461])
    detected_keypoint[1][461] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][462])
    detected_keypoint[1][462] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][463])
    detected_keypoint[1][463] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][464])
    detected_keypoint[1][464] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][465])
    detected_keypoint[1][465] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][466])
    detected_keypoint[1][466] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][467])
    detected_keypoint[1][467] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][468])
    detected_keypoint[1][468] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][469])
    detected_keypoint[1][469] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][470])
    detected_keypoint[1][470] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][471])
    detected_keypoint[1][471] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][472])
    detected_keypoint[1][472] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][473])
    detected_keypoint[1][473] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][474])
    detected_keypoint[1][474] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][475])
    detected_keypoint[1][475] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][476])
    detected_keypoint[1][476] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][477])
    detected_keypoint[1][477] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][478])
    detected_keypoint[1][478] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][479])
    detected_keypoint[1][479] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][480])
    detected_keypoint[1][480] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][481])
    detected_keypoint[1][481] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][482])
    detected_keypoint[1][482] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][483])
    detected_keypoint[1][483] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][484])
    detected_keypoint[1][484] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][485])
    detected_keypoint[1][485] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][486])
    detected_keypoint[1][486] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][487])
    detected_keypoint[1][487] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][488])
    detected_keypoint[1][488] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][489])
    detected_keypoint[1][489] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][490])
    detected_keypoint[1][490] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][491])
    detected_keypoint[1][491] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][492])
    detected_keypoint[1][492] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][493])
    detected_keypoint[1][493] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][494])
    detected_keypoint[1][494] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][495])
    detected_keypoint[1][495] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][496])
    detected_keypoint[1][496] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][497])
    detected_keypoint[1][497] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][498])
    detected_keypoint[1][498] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][499])
    detected_keypoint[1][499] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][500])
    detected_keypoint[1][500] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][501])
    detected_keypoint[1][501] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][502])
    detected_keypoint[1][502] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][503])
    detected_keypoint[1][503] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][504])
    detected_keypoint[1][504] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][505])
    detected_keypoint[1][505] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][506])
    detected_keypoint[1][506] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][507])
    detected_keypoint[1][507] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][508])
    detected_keypoint[1][508] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][509])
    detected_keypoint[1][509] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][510])
    detected_keypoint[1][510] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][511])
    detected_keypoint[1][511] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][512])
    detected_keypoint[1][512] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][513])
    detected_keypoint[1][513] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][514])
    detected_keypoint[1][514] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][515])
    detected_keypoint[1][515] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][516])
    detected_keypoint[1][516] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][517])
    detected_keypoint[1][517] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][518])
    detected_keypoint[1][518] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][519])
    detected_keypoint[1][519] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][520])
    detected_keypoint[1][520] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][521])
    detected_keypoint[1][521] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][522])
    detected_keypoint[1][522] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][523])
    detected_keypoint[1][523] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][524])
    detected_keypoint[1][524] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][525])
    detected_keypoint[1][525] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][526])
    detected_keypoint[1][526] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][527])
    detected_keypoint[1][527] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][528])
    detected_keypoint[1][528] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][529])
    detected_keypoint[1][529] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][530])
    detected_keypoint[1][530] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][531])
    detected_keypoint[1][531] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][532])
    detected_keypoint[1][532] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][533])
    detected_keypoint[1][533] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][534])
    detected_keypoint[1][534] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][535])
    detected_keypoint[1][535] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][536])
    detected_keypoint[1][536] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][537])
    detected_keypoint[1][537] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][538])
    detected_keypoint[1][538] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][539])
    detected_keypoint[1][539] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][540])
    detected_keypoint[1][540] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][541])
    detected_keypoint[1][541] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][542])
    detected_keypoint[1][542] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][543])
    detected_keypoint[1][543] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][544])
    detected_keypoint[1][544] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][545])
    detected_keypoint[1][545] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][546])
    detected_keypoint[1][546] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][547])
    detected_keypoint[1][547] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][548])
    detected_keypoint[1][548] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][549])
    detected_keypoint[1][549] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][550])
    detected_keypoint[1][550] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][551])
    detected_keypoint[1][551] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][552])
    detected_keypoint[1][552] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][553])
    detected_keypoint[1][553] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][554])
    detected_keypoint[1][554] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][555])
    detected_keypoint[1][555] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][556])
    detected_keypoint[1][556] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][557])
    detected_keypoint[1][557] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][558])
    detected_keypoint[1][558] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][559])
    detected_keypoint[1][559] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][560])
    detected_keypoint[1][560] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][561])
    detected_keypoint[1][561] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][562])
    detected_keypoint[1][562] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][563])
    detected_keypoint[1][563] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][564])
    detected_keypoint[1][564] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][565])
    detected_keypoint[1][565] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][566])
    detected_keypoint[1][566] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][567])
    detected_keypoint[1][567] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][568])
    detected_keypoint[1][568] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][569])
    detected_keypoint[1][569] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][570])
    detected_keypoint[1][570] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][571])
    detected_keypoint[1][571] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][572])
    detected_keypoint[1][572] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][573])
    detected_keypoint[1][573] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][574])
    detected_keypoint[1][574] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][575])
    detected_keypoint[1][575] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][576])
    detected_keypoint[1][576] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][577])
    detected_keypoint[1][577] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][578])
    detected_keypoint[1][578] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][579])
    detected_keypoint[1][579] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][580])
    detected_keypoint[1][580] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][581])
    detected_keypoint[1][581] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][582])
    detected_keypoint[1][582] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][583])
    detected_keypoint[1][583] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][584])
    detected_keypoint[1][584] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][585])
    detected_keypoint[1][585] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][586])
    detected_keypoint[1][586] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][587])
    detected_keypoint[1][587] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][588])
    detected_keypoint[1][588] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][589])
    detected_keypoint[1][589] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][590])
    detected_keypoint[1][590] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][591])
    detected_keypoint[1][591] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][592])
    detected_keypoint[1][592] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][593])
    detected_keypoint[1][593] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][594])
    detected_keypoint[1][594] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][595])
    detected_keypoint[1][595] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][596])
    detected_keypoint[1][596] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][597])
    detected_keypoint[1][597] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][598])
    detected_keypoint[1][598] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][599])
    detected_keypoint[1][599] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][600])
    detected_keypoint[1][600] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][601])
    detected_keypoint[1][601] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][602])
    detected_keypoint[1][602] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][603])
    detected_keypoint[1][603] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][604])
    detected_keypoint[1][604] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][605])
    detected_keypoint[1][605] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][606])
    detected_keypoint[1][606] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][607])
    detected_keypoint[1][607] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][608])
    detected_keypoint[1][608] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][609])
    detected_keypoint[1][609] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][610])
    detected_keypoint[1][610] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][611])
    detected_keypoint[1][611] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][612])
    detected_keypoint[1][612] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][613])
    detected_keypoint[1][613] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][614])
    detected_keypoint[1][614] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][615])
    detected_keypoint[1][615] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][616])
    detected_keypoint[1][616] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][617])
    detected_keypoint[1][617] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][618])
    detected_keypoint[1][618] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][619])
    detected_keypoint[1][619] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][620])
    detected_keypoint[1][620] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][621])
    detected_keypoint[1][621] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][622])
    detected_keypoint[1][622] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][623])
    detected_keypoint[1][623] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][624])
    detected_keypoint[1][624] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][625])
    detected_keypoint[1][625] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][626])
    detected_keypoint[1][626] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][627])
    detected_keypoint[1][627] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][628])
    detected_keypoint[1][628] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][629])
    detected_keypoint[1][629] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][630])
    detected_keypoint[1][630] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][631])
    detected_keypoint[1][631] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][632])
    detected_keypoint[1][632] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][633])
    detected_keypoint[1][633] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][634])
    detected_keypoint[1][634] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][635])
    detected_keypoint[1][635] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][636])
    detected_keypoint[1][636] <= 1'b0;
  else if (current_state==ST_FILTER && detected_keypoint[1][637])
    detected_keypoint[1][637] <= 1'b0;
  else
    detected_keypoint[1] <= 'd0;
end

assign no_keypoint[0] = (|detected_keypoint[0]) ? 0 : 1
assign no_keypoint[1] = (|detected_keypoint[1]) ? 0 : 1

always @(*) begin
  if (detected_keypoint[0][0]) begin
    filter_input_0_0 = buffer_data_3[23:0];
    filter_input_0_1 = buffer_data_2[23:0];
    filter_input_0_2 = blur3x3_dout[23:0];
    current_RowCol_0 = {img_addr, 10'd1};
  end
  else if (detected_keypoint[0][1]) begin
    filter_input_0_0 = buffer_data_3[31:8];
    filter_input_0_1 = buffer_data_2[31:8];
    filter_input_0_2 = blur3x3_dout[31:8];
    current_RowCol_0 = {img_addr, 10'd2};
  end
  else if (detected_keypoint[0][2]) begin
    filter_input_0_0 = buffer_data_3[39:16];
    filter_input_0_1 = buffer_data_2[39:16];
    filter_input_0_2 = blur3x3_dout[39:16];
    current_RowCol_0 = {img_addr, 10'd3};
  end
  else if (detected_keypoint[0][3]) begin
    filter_input_0_0 = buffer_data_3[47:24];
    filter_input_0_1 = buffer_data_2[47:24];
    filter_input_0_2 = blur3x3_dout[47:24];
    current_RowCol_0 = {img_addr, 10'd4};
  end
  else if (detected_keypoint[0][4]) begin
    filter_input_0_0 = buffer_data_3[55:32];
    filter_input_0_1 = buffer_data_2[55:32];
    filter_input_0_2 = blur3x3_dout[55:32];
    current_RowCol_0 = {img_addr, 10'd5};
  end
  else if (detected_keypoint[0][5]) begin
    filter_input_0_0 = buffer_data_3[63:40];
    filter_input_0_1 = buffer_data_2[63:40];
    filter_input_0_2 = blur3x3_dout[63:40];
    current_RowCol_0 = {img_addr, 10'd6};
  end
  else if (detected_keypoint[0][6]) begin
    filter_input_0_0 = buffer_data_3[71:48];
    filter_input_0_1 = buffer_data_2[71:48];
    filter_input_0_2 = blur3x3_dout[71:48];
    current_RowCol_0 = {img_addr, 10'd7};
  end
  else if (detected_keypoint[0][7]) begin
    filter_input_0_0 = buffer_data_3[79:56];
    filter_input_0_1 = buffer_data_2[79:56];
    filter_input_0_2 = blur3x3_dout[79:56];
    current_RowCol_0 = {img_addr, 10'd8};
  end
  else if (detected_keypoint[0][8]) begin
    filter_input_0_0 = buffer_data_3[87:64];
    filter_input_0_1 = buffer_data_2[87:64];
    filter_input_0_2 = blur3x3_dout[87:64];
    current_RowCol_0 = {img_addr, 10'd9};
  end
  else if (detected_keypoint[0][9]) begin
    filter_input_0_0 = buffer_data_3[95:72];
    filter_input_0_1 = buffer_data_2[95:72];
    filter_input_0_2 = blur3x3_dout[95:72];
    current_RowCol_0 = {img_addr, 10'd10};
  end
  else if (detected_keypoint[0][10]) begin
    filter_input_0_0 = buffer_data_3[103:80];
    filter_input_0_1 = buffer_data_2[103:80];
    filter_input_0_2 = blur3x3_dout[103:80];
    current_RowCol_0 = {img_addr, 10'd11};
  end
  else if (detected_keypoint[0][11]) begin
    filter_input_0_0 = buffer_data_3[111:88];
    filter_input_0_1 = buffer_data_2[111:88];
    filter_input_0_2 = blur3x3_dout[111:88];
    current_RowCol_0 = {img_addr, 10'd12};
  end
  else if (detected_keypoint[0][12]) begin
    filter_input_0_0 = buffer_data_3[119:96];
    filter_input_0_1 = buffer_data_2[119:96];
    filter_input_0_2 = blur3x3_dout[119:96];
    current_RowCol_0 = {img_addr, 10'd13};
  end
  else if (detected_keypoint[0][13]) begin
    filter_input_0_0 = buffer_data_3[127:104];
    filter_input_0_1 = buffer_data_2[127:104];
    filter_input_0_2 = blur3x3_dout[127:104];
    current_RowCol_0 = {img_addr, 10'd14};
  end
  else if (detected_keypoint[0][14]) begin
    filter_input_0_0 = buffer_data_3[135:112];
    filter_input_0_1 = buffer_data_2[135:112];
    filter_input_0_2 = blur3x3_dout[135:112];
    current_RowCol_0 = {img_addr, 10'd15};
  end
  else if (detected_keypoint[0][15]) begin
    filter_input_0_0 = buffer_data_3[143:120];
    filter_input_0_1 = buffer_data_2[143:120];
    filter_input_0_2 = blur3x3_dout[143:120];
    current_RowCol_0 = {img_addr, 10'd16};
  end
  else if (detected_keypoint[0][16]) begin
    filter_input_0_0 = buffer_data_3[151:128];
    filter_input_0_1 = buffer_data_2[151:128];
    filter_input_0_2 = blur3x3_dout[151:128];
    current_RowCol_0 = {img_addr, 10'd17};
  end
  else if (detected_keypoint[0][17]) begin
    filter_input_0_0 = buffer_data_3[159:136];
    filter_input_0_1 = buffer_data_2[159:136];
    filter_input_0_2 = blur3x3_dout[159:136];
    current_RowCol_0 = {img_addr, 10'd18};
  end
  else if (detected_keypoint[0][18]) begin
    filter_input_0_0 = buffer_data_3[167:144];
    filter_input_0_1 = buffer_data_2[167:144];
    filter_input_0_2 = blur3x3_dout[167:144];
    current_RowCol_0 = {img_addr, 10'd19};
  end
  else if (detected_keypoint[0][19]) begin
    filter_input_0_0 = buffer_data_3[175:152];
    filter_input_0_1 = buffer_data_2[175:152];
    filter_input_0_2 = blur3x3_dout[175:152];
    current_RowCol_0 = {img_addr, 10'd20};
  end
  else if (detected_keypoint[0][20]) begin
    filter_input_0_0 = buffer_data_3[183:160];
    filter_input_0_1 = buffer_data_2[183:160];
    filter_input_0_2 = blur3x3_dout[183:160];
    current_RowCol_0 = {img_addr, 10'd21};
  end
  else if (detected_keypoint[0][21]) begin
    filter_input_0_0 = buffer_data_3[191:168];
    filter_input_0_1 = buffer_data_2[191:168];
    filter_input_0_2 = blur3x3_dout[191:168];
    current_RowCol_0 = {img_addr, 10'd22};
  end
  else if (detected_keypoint[0][22]) begin
    filter_input_0_0 = buffer_data_3[199:176];
    filter_input_0_1 = buffer_data_2[199:176];
    filter_input_0_2 = blur3x3_dout[199:176];
    current_RowCol_0 = {img_addr, 10'd23};
  end
  else if (detected_keypoint[0][23]) begin
    filter_input_0_0 = buffer_data_3[207:184];
    filter_input_0_1 = buffer_data_2[207:184];
    filter_input_0_2 = blur3x3_dout[207:184];
    current_RowCol_0 = {img_addr, 10'd24};
  end
  else if (detected_keypoint[0][24]) begin
    filter_input_0_0 = buffer_data_3[215:192];
    filter_input_0_1 = buffer_data_2[215:192];
    filter_input_0_2 = blur3x3_dout[215:192];
    current_RowCol_0 = {img_addr, 10'd25};
  end
  else if (detected_keypoint[0][25]) begin
    filter_input_0_0 = buffer_data_3[223:200];
    filter_input_0_1 = buffer_data_2[223:200];
    filter_input_0_2 = blur3x3_dout[223:200];
    current_RowCol_0 = {img_addr, 10'd26};
  end
  else if (detected_keypoint[0][26]) begin
    filter_input_0_0 = buffer_data_3[231:208];
    filter_input_0_1 = buffer_data_2[231:208];
    filter_input_0_2 = blur3x3_dout[231:208];
    current_RowCol_0 = {img_addr, 10'd27};
  end
  else if (detected_keypoint[0][27]) begin
    filter_input_0_0 = buffer_data_3[239:216];
    filter_input_0_1 = buffer_data_2[239:216];
    filter_input_0_2 = blur3x3_dout[239:216];
    current_RowCol_0 = {img_addr, 10'd28};
  end
  else if (detected_keypoint[0][28]) begin
    filter_input_0_0 = buffer_data_3[247:224];
    filter_input_0_1 = buffer_data_2[247:224];
    filter_input_0_2 = blur3x3_dout[247:224];
    current_RowCol_0 = {img_addr, 10'd29};
  end
  else if (detected_keypoint[0][29]) begin
    filter_input_0_0 = buffer_data_3[255:232];
    filter_input_0_1 = buffer_data_2[255:232];
    filter_input_0_2 = blur3x3_dout[255:232];
    current_RowCol_0 = {img_addr, 10'd30};
  end
  else if (detected_keypoint[0][30]) begin
    filter_input_0_0 = buffer_data_3[263:240];
    filter_input_0_1 = buffer_data_2[263:240];
    filter_input_0_2 = blur3x3_dout[263:240];
    current_RowCol_0 = {img_addr, 10'd31};
  end
  else if (detected_keypoint[0][31]) begin
    filter_input_0_0 = buffer_data_3[271:248];
    filter_input_0_1 = buffer_data_2[271:248];
    filter_input_0_2 = blur3x3_dout[271:248];
    current_RowCol_0 = {img_addr, 10'd32};
  end
  else if (detected_keypoint[0][32]) begin
    filter_input_0_0 = buffer_data_3[279:256];
    filter_input_0_1 = buffer_data_2[279:256];
    filter_input_0_2 = blur3x3_dout[279:256];
    current_RowCol_0 = {img_addr, 10'd33};
  end
  else if (detected_keypoint[0][33]) begin
    filter_input_0_0 = buffer_data_3[287:264];
    filter_input_0_1 = buffer_data_2[287:264];
    filter_input_0_2 = blur3x3_dout[287:264];
    current_RowCol_0 = {img_addr, 10'd34};
  end
  else if (detected_keypoint[0][34]) begin
    filter_input_0_0 = buffer_data_3[295:272];
    filter_input_0_1 = buffer_data_2[295:272];
    filter_input_0_2 = blur3x3_dout[295:272];
    current_RowCol_0 = {img_addr, 10'd35};
  end
  else if (detected_keypoint[0][35]) begin
    filter_input_0_0 = buffer_data_3[303:280];
    filter_input_0_1 = buffer_data_2[303:280];
    filter_input_0_2 = blur3x3_dout[303:280];
    current_RowCol_0 = {img_addr, 10'd36};
  end
  else if (detected_keypoint[0][36]) begin
    filter_input_0_0 = buffer_data_3[311:288];
    filter_input_0_1 = buffer_data_2[311:288];
    filter_input_0_2 = blur3x3_dout[311:288];
    current_RowCol_0 = {img_addr, 10'd37};
  end
  else if (detected_keypoint[0][37]) begin
    filter_input_0_0 = buffer_data_3[319:296];
    filter_input_0_1 = buffer_data_2[319:296];
    filter_input_0_2 = blur3x3_dout[319:296];
    current_RowCol_0 = {img_addr, 10'd38};
  end
  else if (detected_keypoint[0][38]) begin
    filter_input_0_0 = buffer_data_3[327:304];
    filter_input_0_1 = buffer_data_2[327:304];
    filter_input_0_2 = blur3x3_dout[327:304];
    current_RowCol_0 = {img_addr, 10'd39};
  end
  else if (detected_keypoint[0][39]) begin
    filter_input_0_0 = buffer_data_3[335:312];
    filter_input_0_1 = buffer_data_2[335:312];
    filter_input_0_2 = blur3x3_dout[335:312];
    current_RowCol_0 = {img_addr, 10'd40};
  end
  else if (detected_keypoint[0][40]) begin
    filter_input_0_0 = buffer_data_3[343:320];
    filter_input_0_1 = buffer_data_2[343:320];
    filter_input_0_2 = blur3x3_dout[343:320];
    current_RowCol_0 = {img_addr, 10'd41};
  end
  else if (detected_keypoint[0][41]) begin
    filter_input_0_0 = buffer_data_3[351:328];
    filter_input_0_1 = buffer_data_2[351:328];
    filter_input_0_2 = blur3x3_dout[351:328];
    current_RowCol_0 = {img_addr, 10'd42};
  end
  else if (detected_keypoint[0][42]) begin
    filter_input_0_0 = buffer_data_3[359:336];
    filter_input_0_1 = buffer_data_2[359:336];
    filter_input_0_2 = blur3x3_dout[359:336];
    current_RowCol_0 = {img_addr, 10'd43};
  end
  else if (detected_keypoint[0][43]) begin
    filter_input_0_0 = buffer_data_3[367:344];
    filter_input_0_1 = buffer_data_2[367:344];
    filter_input_0_2 = blur3x3_dout[367:344];
    current_RowCol_0 = {img_addr, 10'd44};
  end
  else if (detected_keypoint[0][44]) begin
    filter_input_0_0 = buffer_data_3[375:352];
    filter_input_0_1 = buffer_data_2[375:352];
    filter_input_0_2 = blur3x3_dout[375:352];
    current_RowCol_0 = {img_addr, 10'd45};
  end
  else if (detected_keypoint[0][45]) begin
    filter_input_0_0 = buffer_data_3[383:360];
    filter_input_0_1 = buffer_data_2[383:360];
    filter_input_0_2 = blur3x3_dout[383:360];
    current_RowCol_0 = {img_addr, 10'd46};
  end
  else if (detected_keypoint[0][46]) begin
    filter_input_0_0 = buffer_data_3[391:368];
    filter_input_0_1 = buffer_data_2[391:368];
    filter_input_0_2 = blur3x3_dout[391:368];
    current_RowCol_0 = {img_addr, 10'd47};
  end
  else if (detected_keypoint[0][47]) begin
    filter_input_0_0 = buffer_data_3[399:376];
    filter_input_0_1 = buffer_data_2[399:376];
    filter_input_0_2 = blur3x3_dout[399:376];
    current_RowCol_0 = {img_addr, 10'd48};
  end
  else if (detected_keypoint[0][48]) begin
    filter_input_0_0 = buffer_data_3[407:384];
    filter_input_0_1 = buffer_data_2[407:384];
    filter_input_0_2 = blur3x3_dout[407:384];
    current_RowCol_0 = {img_addr, 10'd49};
  end
  else if (detected_keypoint[0][49]) begin
    filter_input_0_0 = buffer_data_3[415:392];
    filter_input_0_1 = buffer_data_2[415:392];
    filter_input_0_2 = blur3x3_dout[415:392];
    current_RowCol_0 = {img_addr, 10'd50};
  end
  else if (detected_keypoint[0][50]) begin
    filter_input_0_0 = buffer_data_3[423:400];
    filter_input_0_1 = buffer_data_2[423:400];
    filter_input_0_2 = blur3x3_dout[423:400];
    current_RowCol_0 = {img_addr, 10'd51};
  end
  else if (detected_keypoint[0][51]) begin
    filter_input_0_0 = buffer_data_3[431:408];
    filter_input_0_1 = buffer_data_2[431:408];
    filter_input_0_2 = blur3x3_dout[431:408];
    current_RowCol_0 = {img_addr, 10'd52};
  end
  else if (detected_keypoint[0][52]) begin
    filter_input_0_0 = buffer_data_3[439:416];
    filter_input_0_1 = buffer_data_2[439:416];
    filter_input_0_2 = blur3x3_dout[439:416];
    current_RowCol_0 = {img_addr, 10'd53};
  end
  else if (detected_keypoint[0][53]) begin
    filter_input_0_0 = buffer_data_3[447:424];
    filter_input_0_1 = buffer_data_2[447:424];
    filter_input_0_2 = blur3x3_dout[447:424];
    current_RowCol_0 = {img_addr, 10'd54};
  end
  else if (detected_keypoint[0][54]) begin
    filter_input_0_0 = buffer_data_3[455:432];
    filter_input_0_1 = buffer_data_2[455:432];
    filter_input_0_2 = blur3x3_dout[455:432];
    current_RowCol_0 = {img_addr, 10'd55};
  end
  else if (detected_keypoint[0][55]) begin
    filter_input_0_0 = buffer_data_3[463:440];
    filter_input_0_1 = buffer_data_2[463:440];
    filter_input_0_2 = blur3x3_dout[463:440];
    current_RowCol_0 = {img_addr, 10'd56};
  end
  else if (detected_keypoint[0][56]) begin
    filter_input_0_0 = buffer_data_3[471:448];
    filter_input_0_1 = buffer_data_2[471:448];
    filter_input_0_2 = blur3x3_dout[471:448];
    current_RowCol_0 = {img_addr, 10'd57};
  end
  else if (detected_keypoint[0][57]) begin
    filter_input_0_0 = buffer_data_3[479:456];
    filter_input_0_1 = buffer_data_2[479:456];
    filter_input_0_2 = blur3x3_dout[479:456];
    current_RowCol_0 = {img_addr, 10'd58};
  end
  else if (detected_keypoint[0][58]) begin
    filter_input_0_0 = buffer_data_3[487:464];
    filter_input_0_1 = buffer_data_2[487:464];
    filter_input_0_2 = blur3x3_dout[487:464];
    current_RowCol_0 = {img_addr, 10'd59};
  end
  else if (detected_keypoint[0][59]) begin
    filter_input_0_0 = buffer_data_3[495:472];
    filter_input_0_1 = buffer_data_2[495:472];
    filter_input_0_2 = blur3x3_dout[495:472];
    current_RowCol_0 = {img_addr, 10'd60};
  end
  else if (detected_keypoint[0][60]) begin
    filter_input_0_0 = buffer_data_3[503:480];
    filter_input_0_1 = buffer_data_2[503:480];
    filter_input_0_2 = blur3x3_dout[503:480];
    current_RowCol_0 = {img_addr, 10'd61};
  end
  else if (detected_keypoint[0][61]) begin
    filter_input_0_0 = buffer_data_3[511:488];
    filter_input_0_1 = buffer_data_2[511:488];
    filter_input_0_2 = blur3x3_dout[511:488];
    current_RowCol_0 = {img_addr, 10'd62};
  end
  else if (detected_keypoint[0][62]) begin
    filter_input_0_0 = buffer_data_3[519:496];
    filter_input_0_1 = buffer_data_2[519:496];
    filter_input_0_2 = blur3x3_dout[519:496];
    current_RowCol_0 = {img_addr, 10'd63};
  end
  else if (detected_keypoint[0][63]) begin
    filter_input_0_0 = buffer_data_3[527:504];
    filter_input_0_1 = buffer_data_2[527:504];
    filter_input_0_2 = blur3x3_dout[527:504];
    current_RowCol_0 = {img_addr, 10'd64};
  end
  else if (detected_keypoint[0][64]) begin
    filter_input_0_0 = buffer_data_3[535:512];
    filter_input_0_1 = buffer_data_2[535:512];
    filter_input_0_2 = blur3x3_dout[535:512];
    current_RowCol_0 = {img_addr, 10'd65};
  end
  else if (detected_keypoint[0][65]) begin
    filter_input_0_0 = buffer_data_3[543:520];
    filter_input_0_1 = buffer_data_2[543:520];
    filter_input_0_2 = blur3x3_dout[543:520];
    current_RowCol_0 = {img_addr, 10'd66};
  end
  else if (detected_keypoint[0][66]) begin
    filter_input_0_0 = buffer_data_3[551:528];
    filter_input_0_1 = buffer_data_2[551:528];
    filter_input_0_2 = blur3x3_dout[551:528];
    current_RowCol_0 = {img_addr, 10'd67};
  end
  else if (detected_keypoint[0][67]) begin
    filter_input_0_0 = buffer_data_3[559:536];
    filter_input_0_1 = buffer_data_2[559:536];
    filter_input_0_2 = blur3x3_dout[559:536];
    current_RowCol_0 = {img_addr, 10'd68};
  end
  else if (detected_keypoint[0][68]) begin
    filter_input_0_0 = buffer_data_3[567:544];
    filter_input_0_1 = buffer_data_2[567:544];
    filter_input_0_2 = blur3x3_dout[567:544];
    current_RowCol_0 = {img_addr, 10'd69};
  end
  else if (detected_keypoint[0][69]) begin
    filter_input_0_0 = buffer_data_3[575:552];
    filter_input_0_1 = buffer_data_2[575:552];
    filter_input_0_2 = blur3x3_dout[575:552];
    current_RowCol_0 = {img_addr, 10'd70};
  end
  else if (detected_keypoint[0][70]) begin
    filter_input_0_0 = buffer_data_3[583:560];
    filter_input_0_1 = buffer_data_2[583:560];
    filter_input_0_2 = blur3x3_dout[583:560];
    current_RowCol_0 = {img_addr, 10'd71};
  end
  else if (detected_keypoint[0][71]) begin
    filter_input_0_0 = buffer_data_3[591:568];
    filter_input_0_1 = buffer_data_2[591:568];
    filter_input_0_2 = blur3x3_dout[591:568];
    current_RowCol_0 = {img_addr, 10'd72};
  end
  else if (detected_keypoint[0][72]) begin
    filter_input_0_0 = buffer_data_3[599:576];
    filter_input_0_1 = buffer_data_2[599:576];
    filter_input_0_2 = blur3x3_dout[599:576];
    current_RowCol_0 = {img_addr, 10'd73};
  end
  else if (detected_keypoint[0][73]) begin
    filter_input_0_0 = buffer_data_3[607:584];
    filter_input_0_1 = buffer_data_2[607:584];
    filter_input_0_2 = blur3x3_dout[607:584];
    current_RowCol_0 = {img_addr, 10'd74};
  end
  else if (detected_keypoint[0][74]) begin
    filter_input_0_0 = buffer_data_3[615:592];
    filter_input_0_1 = buffer_data_2[615:592];
    filter_input_0_2 = blur3x3_dout[615:592];
    current_RowCol_0 = {img_addr, 10'd75};
  end
  else if (detected_keypoint[0][75]) begin
    filter_input_0_0 = buffer_data_3[623:600];
    filter_input_0_1 = buffer_data_2[623:600];
    filter_input_0_2 = blur3x3_dout[623:600];
    current_RowCol_0 = {img_addr, 10'd76};
  end
  else if (detected_keypoint[0][76]) begin
    filter_input_0_0 = buffer_data_3[631:608];
    filter_input_0_1 = buffer_data_2[631:608];
    filter_input_0_2 = blur3x3_dout[631:608];
    current_RowCol_0 = {img_addr, 10'd77};
  end
  else if (detected_keypoint[0][77]) begin
    filter_input_0_0 = buffer_data_3[639:616];
    filter_input_0_1 = buffer_data_2[639:616];
    filter_input_0_2 = blur3x3_dout[639:616];
    current_RowCol_0 = {img_addr, 10'd78};
  end
  else if (detected_keypoint[0][78]) begin
    filter_input_0_0 = buffer_data_3[647:624];
    filter_input_0_1 = buffer_data_2[647:624];
    filter_input_0_2 = blur3x3_dout[647:624];
    current_RowCol_0 = {img_addr, 10'd79};
  end
  else if (detected_keypoint[0][79]) begin
    filter_input_0_0 = buffer_data_3[655:632];
    filter_input_0_1 = buffer_data_2[655:632];
    filter_input_0_2 = blur3x3_dout[655:632];
    current_RowCol_0 = {img_addr, 10'd80};
  end
  else if (detected_keypoint[0][80]) begin
    filter_input_0_0 = buffer_data_3[663:640];
    filter_input_0_1 = buffer_data_2[663:640];
    filter_input_0_2 = blur3x3_dout[663:640];
    current_RowCol_0 = {img_addr, 10'd81};
  end
  else if (detected_keypoint[0][81]) begin
    filter_input_0_0 = buffer_data_3[671:648];
    filter_input_0_1 = buffer_data_2[671:648];
    filter_input_0_2 = blur3x3_dout[671:648];
    current_RowCol_0 = {img_addr, 10'd82};
  end
  else if (detected_keypoint[0][82]) begin
    filter_input_0_0 = buffer_data_3[679:656];
    filter_input_0_1 = buffer_data_2[679:656];
    filter_input_0_2 = blur3x3_dout[679:656];
    current_RowCol_0 = {img_addr, 10'd83};
  end
  else if (detected_keypoint[0][83]) begin
    filter_input_0_0 = buffer_data_3[687:664];
    filter_input_0_1 = buffer_data_2[687:664];
    filter_input_0_2 = blur3x3_dout[687:664];
    current_RowCol_0 = {img_addr, 10'd84};
  end
  else if (detected_keypoint[0][84]) begin
    filter_input_0_0 = buffer_data_3[695:672];
    filter_input_0_1 = buffer_data_2[695:672];
    filter_input_0_2 = blur3x3_dout[695:672];
    current_RowCol_0 = {img_addr, 10'd85};
  end
  else if (detected_keypoint[0][85]) begin
    filter_input_0_0 = buffer_data_3[703:680];
    filter_input_0_1 = buffer_data_2[703:680];
    filter_input_0_2 = blur3x3_dout[703:680];
    current_RowCol_0 = {img_addr, 10'd86};
  end
  else if (detected_keypoint[0][86]) begin
    filter_input_0_0 = buffer_data_3[711:688];
    filter_input_0_1 = buffer_data_2[711:688];
    filter_input_0_2 = blur3x3_dout[711:688];
    current_RowCol_0 = {img_addr, 10'd87};
  end
  else if (detected_keypoint[0][87]) begin
    filter_input_0_0 = buffer_data_3[719:696];
    filter_input_0_1 = buffer_data_2[719:696];
    filter_input_0_2 = blur3x3_dout[719:696];
    current_RowCol_0 = {img_addr, 10'd88};
  end
  else if (detected_keypoint[0][88]) begin
    filter_input_0_0 = buffer_data_3[727:704];
    filter_input_0_1 = buffer_data_2[727:704];
    filter_input_0_2 = blur3x3_dout[727:704];
    current_RowCol_0 = {img_addr, 10'd89};
  end
  else if (detected_keypoint[0][89]) begin
    filter_input_0_0 = buffer_data_3[735:712];
    filter_input_0_1 = buffer_data_2[735:712];
    filter_input_0_2 = blur3x3_dout[735:712];
    current_RowCol_0 = {img_addr, 10'd90};
  end
  else if (detected_keypoint[0][90]) begin
    filter_input_0_0 = buffer_data_3[743:720];
    filter_input_0_1 = buffer_data_2[743:720];
    filter_input_0_2 = blur3x3_dout[743:720];
    current_RowCol_0 = {img_addr, 10'd91};
  end
  else if (detected_keypoint[0][91]) begin
    filter_input_0_0 = buffer_data_3[751:728];
    filter_input_0_1 = buffer_data_2[751:728];
    filter_input_0_2 = blur3x3_dout[751:728];
    current_RowCol_0 = {img_addr, 10'd92};
  end
  else if (detected_keypoint[0][92]) begin
    filter_input_0_0 = buffer_data_3[759:736];
    filter_input_0_1 = buffer_data_2[759:736];
    filter_input_0_2 = blur3x3_dout[759:736];
    current_RowCol_0 = {img_addr, 10'd93};
  end
  else if (detected_keypoint[0][93]) begin
    filter_input_0_0 = buffer_data_3[767:744];
    filter_input_0_1 = buffer_data_2[767:744];
    filter_input_0_2 = blur3x3_dout[767:744];
    current_RowCol_0 = {img_addr, 10'd94};
  end
  else if (detected_keypoint[0][94]) begin
    filter_input_0_0 = buffer_data_3[775:752];
    filter_input_0_1 = buffer_data_2[775:752];
    filter_input_0_2 = blur3x3_dout[775:752];
    current_RowCol_0 = {img_addr, 10'd95};
  end
  else if (detected_keypoint[0][95]) begin
    filter_input_0_0 = buffer_data_3[783:760];
    filter_input_0_1 = buffer_data_2[783:760];
    filter_input_0_2 = blur3x3_dout[783:760];
    current_RowCol_0 = {img_addr, 10'd96};
  end
  else if (detected_keypoint[0][96]) begin
    filter_input_0_0 = buffer_data_3[791:768];
    filter_input_0_1 = buffer_data_2[791:768];
    filter_input_0_2 = blur3x3_dout[791:768];
    current_RowCol_0 = {img_addr, 10'd97};
  end
  else if (detected_keypoint[0][97]) begin
    filter_input_0_0 = buffer_data_3[799:776];
    filter_input_0_1 = buffer_data_2[799:776];
    filter_input_0_2 = blur3x3_dout[799:776];
    current_RowCol_0 = {img_addr, 10'd98};
  end
  else if (detected_keypoint[0][98]) begin
    filter_input_0_0 = buffer_data_3[807:784];
    filter_input_0_1 = buffer_data_2[807:784];
    filter_input_0_2 = blur3x3_dout[807:784];
    current_RowCol_0 = {img_addr, 10'd99};
  end
  else if (detected_keypoint[0][99]) begin
    filter_input_0_0 = buffer_data_3[815:792];
    filter_input_0_1 = buffer_data_2[815:792];
    filter_input_0_2 = blur3x3_dout[815:792];
    current_RowCol_0 = {img_addr, 10'd100};
  end
  else if (detected_keypoint[0][100]) begin
    filter_input_0_0 = buffer_data_3[823:800];
    filter_input_0_1 = buffer_data_2[823:800];
    filter_input_0_2 = blur3x3_dout[823:800];
    current_RowCol_0 = {img_addr, 10'd101};
  end
  else if (detected_keypoint[0][101]) begin
    filter_input_0_0 = buffer_data_3[831:808];
    filter_input_0_1 = buffer_data_2[831:808];
    filter_input_0_2 = blur3x3_dout[831:808];
    current_RowCol_0 = {img_addr, 10'd102};
  end
  else if (detected_keypoint[0][102]) begin
    filter_input_0_0 = buffer_data_3[839:816];
    filter_input_0_1 = buffer_data_2[839:816];
    filter_input_0_2 = blur3x3_dout[839:816];
    current_RowCol_0 = {img_addr, 10'd103};
  end
  else if (detected_keypoint[0][103]) begin
    filter_input_0_0 = buffer_data_3[847:824];
    filter_input_0_1 = buffer_data_2[847:824];
    filter_input_0_2 = blur3x3_dout[847:824];
    current_RowCol_0 = {img_addr, 10'd104};
  end
  else if (detected_keypoint[0][104]) begin
    filter_input_0_0 = buffer_data_3[855:832];
    filter_input_0_1 = buffer_data_2[855:832];
    filter_input_0_2 = blur3x3_dout[855:832];
    current_RowCol_0 = {img_addr, 10'd105};
  end
  else if (detected_keypoint[0][105]) begin
    filter_input_0_0 = buffer_data_3[863:840];
    filter_input_0_1 = buffer_data_2[863:840];
    filter_input_0_2 = blur3x3_dout[863:840];
    current_RowCol_0 = {img_addr, 10'd106};
  end
  else if (detected_keypoint[0][106]) begin
    filter_input_0_0 = buffer_data_3[871:848];
    filter_input_0_1 = buffer_data_2[871:848];
    filter_input_0_2 = blur3x3_dout[871:848];
    current_RowCol_0 = {img_addr, 10'd107};
  end
  else if (detected_keypoint[0][107]) begin
    filter_input_0_0 = buffer_data_3[879:856];
    filter_input_0_1 = buffer_data_2[879:856];
    filter_input_0_2 = blur3x3_dout[879:856];
    current_RowCol_0 = {img_addr, 10'd108};
  end
  else if (detected_keypoint[0][108]) begin
    filter_input_0_0 = buffer_data_3[887:864];
    filter_input_0_1 = buffer_data_2[887:864];
    filter_input_0_2 = blur3x3_dout[887:864];
    current_RowCol_0 = {img_addr, 10'd109};
  end
  else if (detected_keypoint[0][109]) begin
    filter_input_0_0 = buffer_data_3[895:872];
    filter_input_0_1 = buffer_data_2[895:872];
    filter_input_0_2 = blur3x3_dout[895:872];
    current_RowCol_0 = {img_addr, 10'd110};
  end
  else if (detected_keypoint[0][110]) begin
    filter_input_0_0 = buffer_data_3[903:880];
    filter_input_0_1 = buffer_data_2[903:880];
    filter_input_0_2 = blur3x3_dout[903:880];
    current_RowCol_0 = {img_addr, 10'd111};
  end
  else if (detected_keypoint[0][111]) begin
    filter_input_0_0 = buffer_data_3[911:888];
    filter_input_0_1 = buffer_data_2[911:888];
    filter_input_0_2 = blur3x3_dout[911:888];
    current_RowCol_0 = {img_addr, 10'd112};
  end
  else if (detected_keypoint[0][112]) begin
    filter_input_0_0 = buffer_data_3[919:896];
    filter_input_0_1 = buffer_data_2[919:896];
    filter_input_0_2 = blur3x3_dout[919:896];
    current_RowCol_0 = {img_addr, 10'd113};
  end
  else if (detected_keypoint[0][113]) begin
    filter_input_0_0 = buffer_data_3[927:904];
    filter_input_0_1 = buffer_data_2[927:904];
    filter_input_0_2 = blur3x3_dout[927:904];
    current_RowCol_0 = {img_addr, 10'd114};
  end
  else if (detected_keypoint[0][114]) begin
    filter_input_0_0 = buffer_data_3[935:912];
    filter_input_0_1 = buffer_data_2[935:912];
    filter_input_0_2 = blur3x3_dout[935:912];
    current_RowCol_0 = {img_addr, 10'd115};
  end
  else if (detected_keypoint[0][115]) begin
    filter_input_0_0 = buffer_data_3[943:920];
    filter_input_0_1 = buffer_data_2[943:920];
    filter_input_0_2 = blur3x3_dout[943:920];
    current_RowCol_0 = {img_addr, 10'd116};
  end
  else if (detected_keypoint[0][116]) begin
    filter_input_0_0 = buffer_data_3[951:928];
    filter_input_0_1 = buffer_data_2[951:928];
    filter_input_0_2 = blur3x3_dout[951:928];
    current_RowCol_0 = {img_addr, 10'd117};
  end
  else if (detected_keypoint[0][117]) begin
    filter_input_0_0 = buffer_data_3[959:936];
    filter_input_0_1 = buffer_data_2[959:936];
    filter_input_0_2 = blur3x3_dout[959:936];
    current_RowCol_0 = {img_addr, 10'd118};
  end
  else if (detected_keypoint[0][118]) begin
    filter_input_0_0 = buffer_data_3[967:944];
    filter_input_0_1 = buffer_data_2[967:944];
    filter_input_0_2 = blur3x3_dout[967:944];
    current_RowCol_0 = {img_addr, 10'd119};
  end
  else if (detected_keypoint[0][119]) begin
    filter_input_0_0 = buffer_data_3[975:952];
    filter_input_0_1 = buffer_data_2[975:952];
    filter_input_0_2 = blur3x3_dout[975:952];
    current_RowCol_0 = {img_addr, 10'd120};
  end
  else if (detected_keypoint[0][120]) begin
    filter_input_0_0 = buffer_data_3[983:960];
    filter_input_0_1 = buffer_data_2[983:960];
    filter_input_0_2 = blur3x3_dout[983:960];
    current_RowCol_0 = {img_addr, 10'd121};
  end
  else if (detected_keypoint[0][121]) begin
    filter_input_0_0 = buffer_data_3[991:968];
    filter_input_0_1 = buffer_data_2[991:968];
    filter_input_0_2 = blur3x3_dout[991:968];
    current_RowCol_0 = {img_addr, 10'd122};
  end
  else if (detected_keypoint[0][122]) begin
    filter_input_0_0 = buffer_data_3[999:976];
    filter_input_0_1 = buffer_data_2[999:976];
    filter_input_0_2 = blur3x3_dout[999:976];
    current_RowCol_0 = {img_addr, 10'd123};
  end
  else if (detected_keypoint[0][123]) begin
    filter_input_0_0 = buffer_data_3[1007:984];
    filter_input_0_1 = buffer_data_2[1007:984];
    filter_input_0_2 = blur3x3_dout[1007:984];
    current_RowCol_0 = {img_addr, 10'd124};
  end
  else if (detected_keypoint[0][124]) begin
    filter_input_0_0 = buffer_data_3[1015:992];
    filter_input_0_1 = buffer_data_2[1015:992];
    filter_input_0_2 = blur3x3_dout[1015:992];
    current_RowCol_0 = {img_addr, 10'd125};
  end
  else if (detected_keypoint[0][125]) begin
    filter_input_0_0 = buffer_data_3[1023:1000];
    filter_input_0_1 = buffer_data_2[1023:1000];
    filter_input_0_2 = blur3x3_dout[1023:1000];
    current_RowCol_0 = {img_addr, 10'd126};
  end
  else if (detected_keypoint[0][126]) begin
    filter_input_0_0 = buffer_data_3[1031:1008];
    filter_input_0_1 = buffer_data_2[1031:1008];
    filter_input_0_2 = blur3x3_dout[1031:1008];
    current_RowCol_0 = {img_addr, 10'd127};
  end
  else if (detected_keypoint[0][127]) begin
    filter_input_0_0 = buffer_data_3[1039:1016];
    filter_input_0_1 = buffer_data_2[1039:1016];
    filter_input_0_2 = blur3x3_dout[1039:1016];
    current_RowCol_0 = {img_addr, 10'd128};
  end
  else if (detected_keypoint[0][128]) begin
    filter_input_0_0 = buffer_data_3[1047:1024];
    filter_input_0_1 = buffer_data_2[1047:1024];
    filter_input_0_2 = blur3x3_dout[1047:1024];
    current_RowCol_0 = {img_addr, 10'd129};
  end
  else if (detected_keypoint[0][129]) begin
    filter_input_0_0 = buffer_data_3[1055:1032];
    filter_input_0_1 = buffer_data_2[1055:1032];
    filter_input_0_2 = blur3x3_dout[1055:1032];
    current_RowCol_0 = {img_addr, 10'd130};
  end
  else if (detected_keypoint[0][130]) begin
    filter_input_0_0 = buffer_data_3[1063:1040];
    filter_input_0_1 = buffer_data_2[1063:1040];
    filter_input_0_2 = blur3x3_dout[1063:1040];
    current_RowCol_0 = {img_addr, 10'd131};
  end
  else if (detected_keypoint[0][131]) begin
    filter_input_0_0 = buffer_data_3[1071:1048];
    filter_input_0_1 = buffer_data_2[1071:1048];
    filter_input_0_2 = blur3x3_dout[1071:1048];
    current_RowCol_0 = {img_addr, 10'd132};
  end
  else if (detected_keypoint[0][132]) begin
    filter_input_0_0 = buffer_data_3[1079:1056];
    filter_input_0_1 = buffer_data_2[1079:1056];
    filter_input_0_2 = blur3x3_dout[1079:1056];
    current_RowCol_0 = {img_addr, 10'd133};
  end
  else if (detected_keypoint[0][133]) begin
    filter_input_0_0 = buffer_data_3[1087:1064];
    filter_input_0_1 = buffer_data_2[1087:1064];
    filter_input_0_2 = blur3x3_dout[1087:1064];
    current_RowCol_0 = {img_addr, 10'd134};
  end
  else if (detected_keypoint[0][134]) begin
    filter_input_0_0 = buffer_data_3[1095:1072];
    filter_input_0_1 = buffer_data_2[1095:1072];
    filter_input_0_2 = blur3x3_dout[1095:1072];
    current_RowCol_0 = {img_addr, 10'd135};
  end
  else if (detected_keypoint[0][135]) begin
    filter_input_0_0 = buffer_data_3[1103:1080];
    filter_input_0_1 = buffer_data_2[1103:1080];
    filter_input_0_2 = blur3x3_dout[1103:1080];
    current_RowCol_0 = {img_addr, 10'd136};
  end
  else if (detected_keypoint[0][136]) begin
    filter_input_0_0 = buffer_data_3[1111:1088];
    filter_input_0_1 = buffer_data_2[1111:1088];
    filter_input_0_2 = blur3x3_dout[1111:1088];
    current_RowCol_0 = {img_addr, 10'd137};
  end
  else if (detected_keypoint[0][137]) begin
    filter_input_0_0 = buffer_data_3[1119:1096];
    filter_input_0_1 = buffer_data_2[1119:1096];
    filter_input_0_2 = blur3x3_dout[1119:1096];
    current_RowCol_0 = {img_addr, 10'd138};
  end
  else if (detected_keypoint[0][138]) begin
    filter_input_0_0 = buffer_data_3[1127:1104];
    filter_input_0_1 = buffer_data_2[1127:1104];
    filter_input_0_2 = blur3x3_dout[1127:1104];
    current_RowCol_0 = {img_addr, 10'd139};
  end
  else if (detected_keypoint[0][139]) begin
    filter_input_0_0 = buffer_data_3[1135:1112];
    filter_input_0_1 = buffer_data_2[1135:1112];
    filter_input_0_2 = blur3x3_dout[1135:1112];
    current_RowCol_0 = {img_addr, 10'd140};
  end
  else if (detected_keypoint[0][140]) begin
    filter_input_0_0 = buffer_data_3[1143:1120];
    filter_input_0_1 = buffer_data_2[1143:1120];
    filter_input_0_2 = blur3x3_dout[1143:1120];
    current_RowCol_0 = {img_addr, 10'd141};
  end
  else if (detected_keypoint[0][141]) begin
    filter_input_0_0 = buffer_data_3[1151:1128];
    filter_input_0_1 = buffer_data_2[1151:1128];
    filter_input_0_2 = blur3x3_dout[1151:1128];
    current_RowCol_0 = {img_addr, 10'd142};
  end
  else if (detected_keypoint[0][142]) begin
    filter_input_0_0 = buffer_data_3[1159:1136];
    filter_input_0_1 = buffer_data_2[1159:1136];
    filter_input_0_2 = blur3x3_dout[1159:1136];
    current_RowCol_0 = {img_addr, 10'd143};
  end
  else if (detected_keypoint[0][143]) begin
    filter_input_0_0 = buffer_data_3[1167:1144];
    filter_input_0_1 = buffer_data_2[1167:1144];
    filter_input_0_2 = blur3x3_dout[1167:1144];
    current_RowCol_0 = {img_addr, 10'd144};
  end
  else if (detected_keypoint[0][144]) begin
    filter_input_0_0 = buffer_data_3[1175:1152];
    filter_input_0_1 = buffer_data_2[1175:1152];
    filter_input_0_2 = blur3x3_dout[1175:1152];
    current_RowCol_0 = {img_addr, 10'd145};
  end
  else if (detected_keypoint[0][145]) begin
    filter_input_0_0 = buffer_data_3[1183:1160];
    filter_input_0_1 = buffer_data_2[1183:1160];
    filter_input_0_2 = blur3x3_dout[1183:1160];
    current_RowCol_0 = {img_addr, 10'd146};
  end
  else if (detected_keypoint[0][146]) begin
    filter_input_0_0 = buffer_data_3[1191:1168];
    filter_input_0_1 = buffer_data_2[1191:1168];
    filter_input_0_2 = blur3x3_dout[1191:1168];
    current_RowCol_0 = {img_addr, 10'd147};
  end
  else if (detected_keypoint[0][147]) begin
    filter_input_0_0 = buffer_data_3[1199:1176];
    filter_input_0_1 = buffer_data_2[1199:1176];
    filter_input_0_2 = blur3x3_dout[1199:1176];
    current_RowCol_0 = {img_addr, 10'd148};
  end
  else if (detected_keypoint[0][148]) begin
    filter_input_0_0 = buffer_data_3[1207:1184];
    filter_input_0_1 = buffer_data_2[1207:1184];
    filter_input_0_2 = blur3x3_dout[1207:1184];
    current_RowCol_0 = {img_addr, 10'd149};
  end
  else if (detected_keypoint[0][149]) begin
    filter_input_0_0 = buffer_data_3[1215:1192];
    filter_input_0_1 = buffer_data_2[1215:1192];
    filter_input_0_2 = blur3x3_dout[1215:1192];
    current_RowCol_0 = {img_addr, 10'd150};
  end
  else if (detected_keypoint[0][150]) begin
    filter_input_0_0 = buffer_data_3[1223:1200];
    filter_input_0_1 = buffer_data_2[1223:1200];
    filter_input_0_2 = blur3x3_dout[1223:1200];
    current_RowCol_0 = {img_addr, 10'd151};
  end
  else if (detected_keypoint[0][151]) begin
    filter_input_0_0 = buffer_data_3[1231:1208];
    filter_input_0_1 = buffer_data_2[1231:1208];
    filter_input_0_2 = blur3x3_dout[1231:1208];
    current_RowCol_0 = {img_addr, 10'd152};
  end
  else if (detected_keypoint[0][152]) begin
    filter_input_0_0 = buffer_data_3[1239:1216];
    filter_input_0_1 = buffer_data_2[1239:1216];
    filter_input_0_2 = blur3x3_dout[1239:1216];
    current_RowCol_0 = {img_addr, 10'd153};
  end
  else if (detected_keypoint[0][153]) begin
    filter_input_0_0 = buffer_data_3[1247:1224];
    filter_input_0_1 = buffer_data_2[1247:1224];
    filter_input_0_2 = blur3x3_dout[1247:1224];
    current_RowCol_0 = {img_addr, 10'd154};
  end
  else if (detected_keypoint[0][154]) begin
    filter_input_0_0 = buffer_data_3[1255:1232];
    filter_input_0_1 = buffer_data_2[1255:1232];
    filter_input_0_2 = blur3x3_dout[1255:1232];
    current_RowCol_0 = {img_addr, 10'd155};
  end
  else if (detected_keypoint[0][155]) begin
    filter_input_0_0 = buffer_data_3[1263:1240];
    filter_input_0_1 = buffer_data_2[1263:1240];
    filter_input_0_2 = blur3x3_dout[1263:1240];
    current_RowCol_0 = {img_addr, 10'd156};
  end
  else if (detected_keypoint[0][156]) begin
    filter_input_0_0 = buffer_data_3[1271:1248];
    filter_input_0_1 = buffer_data_2[1271:1248];
    filter_input_0_2 = blur3x3_dout[1271:1248];
    current_RowCol_0 = {img_addr, 10'd157};
  end
  else if (detected_keypoint[0][157]) begin
    filter_input_0_0 = buffer_data_3[1279:1256];
    filter_input_0_1 = buffer_data_2[1279:1256];
    filter_input_0_2 = blur3x3_dout[1279:1256];
    current_RowCol_0 = {img_addr, 10'd158};
  end
  else if (detected_keypoint[0][158]) begin
    filter_input_0_0 = buffer_data_3[1287:1264];
    filter_input_0_1 = buffer_data_2[1287:1264];
    filter_input_0_2 = blur3x3_dout[1287:1264];
    current_RowCol_0 = {img_addr, 10'd159};
  end
  else if (detected_keypoint[0][159]) begin
    filter_input_0_0 = buffer_data_3[1295:1272];
    filter_input_0_1 = buffer_data_2[1295:1272];
    filter_input_0_2 = blur3x3_dout[1295:1272];
    current_RowCol_0 = {img_addr, 10'd160};
  end
  else if (detected_keypoint[0][160]) begin
    filter_input_0_0 = buffer_data_3[1303:1280];
    filter_input_0_1 = buffer_data_2[1303:1280];
    filter_input_0_2 = blur3x3_dout[1303:1280];
    current_RowCol_0 = {img_addr, 10'd161};
  end
  else if (detected_keypoint[0][161]) begin
    filter_input_0_0 = buffer_data_3[1311:1288];
    filter_input_0_1 = buffer_data_2[1311:1288];
    filter_input_0_2 = blur3x3_dout[1311:1288];
    current_RowCol_0 = {img_addr, 10'd162};
  end
  else if (detected_keypoint[0][162]) begin
    filter_input_0_0 = buffer_data_3[1319:1296];
    filter_input_0_1 = buffer_data_2[1319:1296];
    filter_input_0_2 = blur3x3_dout[1319:1296];
    current_RowCol_0 = {img_addr, 10'd163};
  end
  else if (detected_keypoint[0][163]) begin
    filter_input_0_0 = buffer_data_3[1327:1304];
    filter_input_0_1 = buffer_data_2[1327:1304];
    filter_input_0_2 = blur3x3_dout[1327:1304];
    current_RowCol_0 = {img_addr, 10'd164};
  end
  else if (detected_keypoint[0][164]) begin
    filter_input_0_0 = buffer_data_3[1335:1312];
    filter_input_0_1 = buffer_data_2[1335:1312];
    filter_input_0_2 = blur3x3_dout[1335:1312];
    current_RowCol_0 = {img_addr, 10'd165};
  end
  else if (detected_keypoint[0][165]) begin
    filter_input_0_0 = buffer_data_3[1343:1320];
    filter_input_0_1 = buffer_data_2[1343:1320];
    filter_input_0_2 = blur3x3_dout[1343:1320];
    current_RowCol_0 = {img_addr, 10'd166};
  end
  else if (detected_keypoint[0][166]) begin
    filter_input_0_0 = buffer_data_3[1351:1328];
    filter_input_0_1 = buffer_data_2[1351:1328];
    filter_input_0_2 = blur3x3_dout[1351:1328];
    current_RowCol_0 = {img_addr, 10'd167};
  end
  else if (detected_keypoint[0][167]) begin
    filter_input_0_0 = buffer_data_3[1359:1336];
    filter_input_0_1 = buffer_data_2[1359:1336];
    filter_input_0_2 = blur3x3_dout[1359:1336];
    current_RowCol_0 = {img_addr, 10'd168};
  end
  else if (detected_keypoint[0][168]) begin
    filter_input_0_0 = buffer_data_3[1367:1344];
    filter_input_0_1 = buffer_data_2[1367:1344];
    filter_input_0_2 = blur3x3_dout[1367:1344];
    current_RowCol_0 = {img_addr, 10'd169};
  end
  else if (detected_keypoint[0][169]) begin
    filter_input_0_0 = buffer_data_3[1375:1352];
    filter_input_0_1 = buffer_data_2[1375:1352];
    filter_input_0_2 = blur3x3_dout[1375:1352];
    current_RowCol_0 = {img_addr, 10'd170};
  end
  else if (detected_keypoint[0][170]) begin
    filter_input_0_0 = buffer_data_3[1383:1360];
    filter_input_0_1 = buffer_data_2[1383:1360];
    filter_input_0_2 = blur3x3_dout[1383:1360];
    current_RowCol_0 = {img_addr, 10'd171};
  end
  else if (detected_keypoint[0][171]) begin
    filter_input_0_0 = buffer_data_3[1391:1368];
    filter_input_0_1 = buffer_data_2[1391:1368];
    filter_input_0_2 = blur3x3_dout[1391:1368];
    current_RowCol_0 = {img_addr, 10'd172};
  end
  else if (detected_keypoint[0][172]) begin
    filter_input_0_0 = buffer_data_3[1399:1376];
    filter_input_0_1 = buffer_data_2[1399:1376];
    filter_input_0_2 = blur3x3_dout[1399:1376];
    current_RowCol_0 = {img_addr, 10'd173};
  end
  else if (detected_keypoint[0][173]) begin
    filter_input_0_0 = buffer_data_3[1407:1384];
    filter_input_0_1 = buffer_data_2[1407:1384];
    filter_input_0_2 = blur3x3_dout[1407:1384];
    current_RowCol_0 = {img_addr, 10'd174};
  end
  else if (detected_keypoint[0][174]) begin
    filter_input_0_0 = buffer_data_3[1415:1392];
    filter_input_0_1 = buffer_data_2[1415:1392];
    filter_input_0_2 = blur3x3_dout[1415:1392];
    current_RowCol_0 = {img_addr, 10'd175};
  end
  else if (detected_keypoint[0][175]) begin
    filter_input_0_0 = buffer_data_3[1423:1400];
    filter_input_0_1 = buffer_data_2[1423:1400];
    filter_input_0_2 = blur3x3_dout[1423:1400];
    current_RowCol_0 = {img_addr, 10'd176};
  end
  else if (detected_keypoint[0][176]) begin
    filter_input_0_0 = buffer_data_3[1431:1408];
    filter_input_0_1 = buffer_data_2[1431:1408];
    filter_input_0_2 = blur3x3_dout[1431:1408];
    current_RowCol_0 = {img_addr, 10'd177};
  end
  else if (detected_keypoint[0][177]) begin
    filter_input_0_0 = buffer_data_3[1439:1416];
    filter_input_0_1 = buffer_data_2[1439:1416];
    filter_input_0_2 = blur3x3_dout[1439:1416];
    current_RowCol_0 = {img_addr, 10'd178};
  end
  else if (detected_keypoint[0][178]) begin
    filter_input_0_0 = buffer_data_3[1447:1424];
    filter_input_0_1 = buffer_data_2[1447:1424];
    filter_input_0_2 = blur3x3_dout[1447:1424];
    current_RowCol_0 = {img_addr, 10'd179};
  end
  else if (detected_keypoint[0][179]) begin
    filter_input_0_0 = buffer_data_3[1455:1432];
    filter_input_0_1 = buffer_data_2[1455:1432];
    filter_input_0_2 = blur3x3_dout[1455:1432];
    current_RowCol_0 = {img_addr, 10'd180};
  end
  else if (detected_keypoint[0][180]) begin
    filter_input_0_0 = buffer_data_3[1463:1440];
    filter_input_0_1 = buffer_data_2[1463:1440];
    filter_input_0_2 = blur3x3_dout[1463:1440];
    current_RowCol_0 = {img_addr, 10'd181};
  end
  else if (detected_keypoint[0][181]) begin
    filter_input_0_0 = buffer_data_3[1471:1448];
    filter_input_0_1 = buffer_data_2[1471:1448];
    filter_input_0_2 = blur3x3_dout[1471:1448];
    current_RowCol_0 = {img_addr, 10'd182};
  end
  else if (detected_keypoint[0][182]) begin
    filter_input_0_0 = buffer_data_3[1479:1456];
    filter_input_0_1 = buffer_data_2[1479:1456];
    filter_input_0_2 = blur3x3_dout[1479:1456];
    current_RowCol_0 = {img_addr, 10'd183};
  end
  else if (detected_keypoint[0][183]) begin
    filter_input_0_0 = buffer_data_3[1487:1464];
    filter_input_0_1 = buffer_data_2[1487:1464];
    filter_input_0_2 = blur3x3_dout[1487:1464];
    current_RowCol_0 = {img_addr, 10'd184};
  end
  else if (detected_keypoint[0][184]) begin
    filter_input_0_0 = buffer_data_3[1495:1472];
    filter_input_0_1 = buffer_data_2[1495:1472];
    filter_input_0_2 = blur3x3_dout[1495:1472];
    current_RowCol_0 = {img_addr, 10'd185};
  end
  else if (detected_keypoint[0][185]) begin
    filter_input_0_0 = buffer_data_3[1503:1480];
    filter_input_0_1 = buffer_data_2[1503:1480];
    filter_input_0_2 = blur3x3_dout[1503:1480];
    current_RowCol_0 = {img_addr, 10'd186};
  end
  else if (detected_keypoint[0][186]) begin
    filter_input_0_0 = buffer_data_3[1511:1488];
    filter_input_0_1 = buffer_data_2[1511:1488];
    filter_input_0_2 = blur3x3_dout[1511:1488];
    current_RowCol_0 = {img_addr, 10'd187};
  end
  else if (detected_keypoint[0][187]) begin
    filter_input_0_0 = buffer_data_3[1519:1496];
    filter_input_0_1 = buffer_data_2[1519:1496];
    filter_input_0_2 = blur3x3_dout[1519:1496];
    current_RowCol_0 = {img_addr, 10'd188};
  end
  else if (detected_keypoint[0][188]) begin
    filter_input_0_0 = buffer_data_3[1527:1504];
    filter_input_0_1 = buffer_data_2[1527:1504];
    filter_input_0_2 = blur3x3_dout[1527:1504];
    current_RowCol_0 = {img_addr, 10'd189};
  end
  else if (detected_keypoint[0][189]) begin
    filter_input_0_0 = buffer_data_3[1535:1512];
    filter_input_0_1 = buffer_data_2[1535:1512];
    filter_input_0_2 = blur3x3_dout[1535:1512];
    current_RowCol_0 = {img_addr, 10'd190};
  end
  else if (detected_keypoint[0][190]) begin
    filter_input_0_0 = buffer_data_3[1543:1520];
    filter_input_0_1 = buffer_data_2[1543:1520];
    filter_input_0_2 = blur3x3_dout[1543:1520];
    current_RowCol_0 = {img_addr, 10'd191};
  end
  else if (detected_keypoint[0][191]) begin
    filter_input_0_0 = buffer_data_3[1551:1528];
    filter_input_0_1 = buffer_data_2[1551:1528];
    filter_input_0_2 = blur3x3_dout[1551:1528];
    current_RowCol_0 = {img_addr, 10'd192};
  end
  else if (detected_keypoint[0][192]) begin
    filter_input_0_0 = buffer_data_3[1559:1536];
    filter_input_0_1 = buffer_data_2[1559:1536];
    filter_input_0_2 = blur3x3_dout[1559:1536];
    current_RowCol_0 = {img_addr, 10'd193};
  end
  else if (detected_keypoint[0][193]) begin
    filter_input_0_0 = buffer_data_3[1567:1544];
    filter_input_0_1 = buffer_data_2[1567:1544];
    filter_input_0_2 = blur3x3_dout[1567:1544];
    current_RowCol_0 = {img_addr, 10'd194};
  end
  else if (detected_keypoint[0][194]) begin
    filter_input_0_0 = buffer_data_3[1575:1552];
    filter_input_0_1 = buffer_data_2[1575:1552];
    filter_input_0_2 = blur3x3_dout[1575:1552];
    current_RowCol_0 = {img_addr, 10'd195};
  end
  else if (detected_keypoint[0][195]) begin
    filter_input_0_0 = buffer_data_3[1583:1560];
    filter_input_0_1 = buffer_data_2[1583:1560];
    filter_input_0_2 = blur3x3_dout[1583:1560];
    current_RowCol_0 = {img_addr, 10'd196};
  end
  else if (detected_keypoint[0][196]) begin
    filter_input_0_0 = buffer_data_3[1591:1568];
    filter_input_0_1 = buffer_data_2[1591:1568];
    filter_input_0_2 = blur3x3_dout[1591:1568];
    current_RowCol_0 = {img_addr, 10'd197};
  end
  else if (detected_keypoint[0][197]) begin
    filter_input_0_0 = buffer_data_3[1599:1576];
    filter_input_0_1 = buffer_data_2[1599:1576];
    filter_input_0_2 = blur3x3_dout[1599:1576];
    current_RowCol_0 = {img_addr, 10'd198};
  end
  else if (detected_keypoint[0][198]) begin
    filter_input_0_0 = buffer_data_3[1607:1584];
    filter_input_0_1 = buffer_data_2[1607:1584];
    filter_input_0_2 = blur3x3_dout[1607:1584];
    current_RowCol_0 = {img_addr, 10'd199};
  end
  else if (detected_keypoint[0][199]) begin
    filter_input_0_0 = buffer_data_3[1615:1592];
    filter_input_0_1 = buffer_data_2[1615:1592];
    filter_input_0_2 = blur3x3_dout[1615:1592];
    current_RowCol_0 = {img_addr, 10'd200};
  end
  else if (detected_keypoint[0][200]) begin
    filter_input_0_0 = buffer_data_3[1623:1600];
    filter_input_0_1 = buffer_data_2[1623:1600];
    filter_input_0_2 = blur3x3_dout[1623:1600];
    current_RowCol_0 = {img_addr, 10'd201};
  end
  else if (detected_keypoint[0][201]) begin
    filter_input_0_0 = buffer_data_3[1631:1608];
    filter_input_0_1 = buffer_data_2[1631:1608];
    filter_input_0_2 = blur3x3_dout[1631:1608];
    current_RowCol_0 = {img_addr, 10'd202};
  end
  else if (detected_keypoint[0][202]) begin
    filter_input_0_0 = buffer_data_3[1639:1616];
    filter_input_0_1 = buffer_data_2[1639:1616];
    filter_input_0_2 = blur3x3_dout[1639:1616];
    current_RowCol_0 = {img_addr, 10'd203};
  end
  else if (detected_keypoint[0][203]) begin
    filter_input_0_0 = buffer_data_3[1647:1624];
    filter_input_0_1 = buffer_data_2[1647:1624];
    filter_input_0_2 = blur3x3_dout[1647:1624];
    current_RowCol_0 = {img_addr, 10'd204};
  end
  else if (detected_keypoint[0][204]) begin
    filter_input_0_0 = buffer_data_3[1655:1632];
    filter_input_0_1 = buffer_data_2[1655:1632];
    filter_input_0_2 = blur3x3_dout[1655:1632];
    current_RowCol_0 = {img_addr, 10'd205};
  end
  else if (detected_keypoint[0][205]) begin
    filter_input_0_0 = buffer_data_3[1663:1640];
    filter_input_0_1 = buffer_data_2[1663:1640];
    filter_input_0_2 = blur3x3_dout[1663:1640];
    current_RowCol_0 = {img_addr, 10'd206};
  end
  else if (detected_keypoint[0][206]) begin
    filter_input_0_0 = buffer_data_3[1671:1648];
    filter_input_0_1 = buffer_data_2[1671:1648];
    filter_input_0_2 = blur3x3_dout[1671:1648];
    current_RowCol_0 = {img_addr, 10'd207};
  end
  else if (detected_keypoint[0][207]) begin
    filter_input_0_0 = buffer_data_3[1679:1656];
    filter_input_0_1 = buffer_data_2[1679:1656];
    filter_input_0_2 = blur3x3_dout[1679:1656];
    current_RowCol_0 = {img_addr, 10'd208};
  end
  else if (detected_keypoint[0][208]) begin
    filter_input_0_0 = buffer_data_3[1687:1664];
    filter_input_0_1 = buffer_data_2[1687:1664];
    filter_input_0_2 = blur3x3_dout[1687:1664];
    current_RowCol_0 = {img_addr, 10'd209};
  end
  else if (detected_keypoint[0][209]) begin
    filter_input_0_0 = buffer_data_3[1695:1672];
    filter_input_0_1 = buffer_data_2[1695:1672];
    filter_input_0_2 = blur3x3_dout[1695:1672];
    current_RowCol_0 = {img_addr, 10'd210};
  end
  else if (detected_keypoint[0][210]) begin
    filter_input_0_0 = buffer_data_3[1703:1680];
    filter_input_0_1 = buffer_data_2[1703:1680];
    filter_input_0_2 = blur3x3_dout[1703:1680];
    current_RowCol_0 = {img_addr, 10'd211};
  end
  else if (detected_keypoint[0][211]) begin
    filter_input_0_0 = buffer_data_3[1711:1688];
    filter_input_0_1 = buffer_data_2[1711:1688];
    filter_input_0_2 = blur3x3_dout[1711:1688];
    current_RowCol_0 = {img_addr, 10'd212};
  end
  else if (detected_keypoint[0][212]) begin
    filter_input_0_0 = buffer_data_3[1719:1696];
    filter_input_0_1 = buffer_data_2[1719:1696];
    filter_input_0_2 = blur3x3_dout[1719:1696];
    current_RowCol_0 = {img_addr, 10'd213};
  end
  else if (detected_keypoint[0][213]) begin
    filter_input_0_0 = buffer_data_3[1727:1704];
    filter_input_0_1 = buffer_data_2[1727:1704];
    filter_input_0_2 = blur3x3_dout[1727:1704];
    current_RowCol_0 = {img_addr, 10'd214};
  end
  else if (detected_keypoint[0][214]) begin
    filter_input_0_0 = buffer_data_3[1735:1712];
    filter_input_0_1 = buffer_data_2[1735:1712];
    filter_input_0_2 = blur3x3_dout[1735:1712];
    current_RowCol_0 = {img_addr, 10'd215};
  end
  else if (detected_keypoint[0][215]) begin
    filter_input_0_0 = buffer_data_3[1743:1720];
    filter_input_0_1 = buffer_data_2[1743:1720];
    filter_input_0_2 = blur3x3_dout[1743:1720];
    current_RowCol_0 = {img_addr, 10'd216};
  end
  else if (detected_keypoint[0][216]) begin
    filter_input_0_0 = buffer_data_3[1751:1728];
    filter_input_0_1 = buffer_data_2[1751:1728];
    filter_input_0_2 = blur3x3_dout[1751:1728];
    current_RowCol_0 = {img_addr, 10'd217};
  end
  else if (detected_keypoint[0][217]) begin
    filter_input_0_0 = buffer_data_3[1759:1736];
    filter_input_0_1 = buffer_data_2[1759:1736];
    filter_input_0_2 = blur3x3_dout[1759:1736];
    current_RowCol_0 = {img_addr, 10'd218};
  end
  else if (detected_keypoint[0][218]) begin
    filter_input_0_0 = buffer_data_3[1767:1744];
    filter_input_0_1 = buffer_data_2[1767:1744];
    filter_input_0_2 = blur3x3_dout[1767:1744];
    current_RowCol_0 = {img_addr, 10'd219};
  end
  else if (detected_keypoint[0][219]) begin
    filter_input_0_0 = buffer_data_3[1775:1752];
    filter_input_0_1 = buffer_data_2[1775:1752];
    filter_input_0_2 = blur3x3_dout[1775:1752];
    current_RowCol_0 = {img_addr, 10'd220};
  end
  else if (detected_keypoint[0][220]) begin
    filter_input_0_0 = buffer_data_3[1783:1760];
    filter_input_0_1 = buffer_data_2[1783:1760];
    filter_input_0_2 = blur3x3_dout[1783:1760];
    current_RowCol_0 = {img_addr, 10'd221};
  end
  else if (detected_keypoint[0][221]) begin
    filter_input_0_0 = buffer_data_3[1791:1768];
    filter_input_0_1 = buffer_data_2[1791:1768];
    filter_input_0_2 = blur3x3_dout[1791:1768];
    current_RowCol_0 = {img_addr, 10'd222};
  end
  else if (detected_keypoint[0][222]) begin
    filter_input_0_0 = buffer_data_3[1799:1776];
    filter_input_0_1 = buffer_data_2[1799:1776];
    filter_input_0_2 = blur3x3_dout[1799:1776];
    current_RowCol_0 = {img_addr, 10'd223};
  end
  else if (detected_keypoint[0][223]) begin
    filter_input_0_0 = buffer_data_3[1807:1784];
    filter_input_0_1 = buffer_data_2[1807:1784];
    filter_input_0_2 = blur3x3_dout[1807:1784];
    current_RowCol_0 = {img_addr, 10'd224};
  end
  else if (detected_keypoint[0][224]) begin
    filter_input_0_0 = buffer_data_3[1815:1792];
    filter_input_0_1 = buffer_data_2[1815:1792];
    filter_input_0_2 = blur3x3_dout[1815:1792];
    current_RowCol_0 = {img_addr, 10'd225};
  end
  else if (detected_keypoint[0][225]) begin
    filter_input_0_0 = buffer_data_3[1823:1800];
    filter_input_0_1 = buffer_data_2[1823:1800];
    filter_input_0_2 = blur3x3_dout[1823:1800];
    current_RowCol_0 = {img_addr, 10'd226};
  end
  else if (detected_keypoint[0][226]) begin
    filter_input_0_0 = buffer_data_3[1831:1808];
    filter_input_0_1 = buffer_data_2[1831:1808];
    filter_input_0_2 = blur3x3_dout[1831:1808];
    current_RowCol_0 = {img_addr, 10'd227};
  end
  else if (detected_keypoint[0][227]) begin
    filter_input_0_0 = buffer_data_3[1839:1816];
    filter_input_0_1 = buffer_data_2[1839:1816];
    filter_input_0_2 = blur3x3_dout[1839:1816];
    current_RowCol_0 = {img_addr, 10'd228};
  end
  else if (detected_keypoint[0][228]) begin
    filter_input_0_0 = buffer_data_3[1847:1824];
    filter_input_0_1 = buffer_data_2[1847:1824];
    filter_input_0_2 = blur3x3_dout[1847:1824];
    current_RowCol_0 = {img_addr, 10'd229};
  end
  else if (detected_keypoint[0][229]) begin
    filter_input_0_0 = buffer_data_3[1855:1832];
    filter_input_0_1 = buffer_data_2[1855:1832];
    filter_input_0_2 = blur3x3_dout[1855:1832];
    current_RowCol_0 = {img_addr, 10'd230};
  end
  else if (detected_keypoint[0][230]) begin
    filter_input_0_0 = buffer_data_3[1863:1840];
    filter_input_0_1 = buffer_data_2[1863:1840];
    filter_input_0_2 = blur3x3_dout[1863:1840];
    current_RowCol_0 = {img_addr, 10'd231};
  end
  else if (detected_keypoint[0][231]) begin
    filter_input_0_0 = buffer_data_3[1871:1848];
    filter_input_0_1 = buffer_data_2[1871:1848];
    filter_input_0_2 = blur3x3_dout[1871:1848];
    current_RowCol_0 = {img_addr, 10'd232};
  end
  else if (detected_keypoint[0][232]) begin
    filter_input_0_0 = buffer_data_3[1879:1856];
    filter_input_0_1 = buffer_data_2[1879:1856];
    filter_input_0_2 = blur3x3_dout[1879:1856];
    current_RowCol_0 = {img_addr, 10'd233};
  end
  else if (detected_keypoint[0][233]) begin
    filter_input_0_0 = buffer_data_3[1887:1864];
    filter_input_0_1 = buffer_data_2[1887:1864];
    filter_input_0_2 = blur3x3_dout[1887:1864];
    current_RowCol_0 = {img_addr, 10'd234};
  end
  else if (detected_keypoint[0][234]) begin
    filter_input_0_0 = buffer_data_3[1895:1872];
    filter_input_0_1 = buffer_data_2[1895:1872];
    filter_input_0_2 = blur3x3_dout[1895:1872];
    current_RowCol_0 = {img_addr, 10'd235};
  end
  else if (detected_keypoint[0][235]) begin
    filter_input_0_0 = buffer_data_3[1903:1880];
    filter_input_0_1 = buffer_data_2[1903:1880];
    filter_input_0_2 = blur3x3_dout[1903:1880];
    current_RowCol_0 = {img_addr, 10'd236};
  end
  else if (detected_keypoint[0][236]) begin
    filter_input_0_0 = buffer_data_3[1911:1888];
    filter_input_0_1 = buffer_data_2[1911:1888];
    filter_input_0_2 = blur3x3_dout[1911:1888];
    current_RowCol_0 = {img_addr, 10'd237};
  end
  else if (detected_keypoint[0][237]) begin
    filter_input_0_0 = buffer_data_3[1919:1896];
    filter_input_0_1 = buffer_data_2[1919:1896];
    filter_input_0_2 = blur3x3_dout[1919:1896];
    current_RowCol_0 = {img_addr, 10'd238};
  end
  else if (detected_keypoint[0][238]) begin
    filter_input_0_0 = buffer_data_3[1927:1904];
    filter_input_0_1 = buffer_data_2[1927:1904];
    filter_input_0_2 = blur3x3_dout[1927:1904];
    current_RowCol_0 = {img_addr, 10'd239};
  end
  else if (detected_keypoint[0][239]) begin
    filter_input_0_0 = buffer_data_3[1935:1912];
    filter_input_0_1 = buffer_data_2[1935:1912];
    filter_input_0_2 = blur3x3_dout[1935:1912];
    current_RowCol_0 = {img_addr, 10'd240};
  end
  else if (detected_keypoint[0][240]) begin
    filter_input_0_0 = buffer_data_3[1943:1920];
    filter_input_0_1 = buffer_data_2[1943:1920];
    filter_input_0_2 = blur3x3_dout[1943:1920];
    current_RowCol_0 = {img_addr, 10'd241};
  end
  else if (detected_keypoint[0][241]) begin
    filter_input_0_0 = buffer_data_3[1951:1928];
    filter_input_0_1 = buffer_data_2[1951:1928];
    filter_input_0_2 = blur3x3_dout[1951:1928];
    current_RowCol_0 = {img_addr, 10'd242};
  end
  else if (detected_keypoint[0][242]) begin
    filter_input_0_0 = buffer_data_3[1959:1936];
    filter_input_0_1 = buffer_data_2[1959:1936];
    filter_input_0_2 = blur3x3_dout[1959:1936];
    current_RowCol_0 = {img_addr, 10'd243};
  end
  else if (detected_keypoint[0][243]) begin
    filter_input_0_0 = buffer_data_3[1967:1944];
    filter_input_0_1 = buffer_data_2[1967:1944];
    filter_input_0_2 = blur3x3_dout[1967:1944];
    current_RowCol_0 = {img_addr, 10'd244};
  end
  else if (detected_keypoint[0][244]) begin
    filter_input_0_0 = buffer_data_3[1975:1952];
    filter_input_0_1 = buffer_data_2[1975:1952];
    filter_input_0_2 = blur3x3_dout[1975:1952];
    current_RowCol_0 = {img_addr, 10'd245};
  end
  else if (detected_keypoint[0][245]) begin
    filter_input_0_0 = buffer_data_3[1983:1960];
    filter_input_0_1 = buffer_data_2[1983:1960];
    filter_input_0_2 = blur3x3_dout[1983:1960];
    current_RowCol_0 = {img_addr, 10'd246};
  end
  else if (detected_keypoint[0][246]) begin
    filter_input_0_0 = buffer_data_3[1991:1968];
    filter_input_0_1 = buffer_data_2[1991:1968];
    filter_input_0_2 = blur3x3_dout[1991:1968];
    current_RowCol_0 = {img_addr, 10'd247};
  end
  else if (detected_keypoint[0][247]) begin
    filter_input_0_0 = buffer_data_3[1999:1976];
    filter_input_0_1 = buffer_data_2[1999:1976];
    filter_input_0_2 = blur3x3_dout[1999:1976];
    current_RowCol_0 = {img_addr, 10'd248};
  end
  else if (detected_keypoint[0][248]) begin
    filter_input_0_0 = buffer_data_3[2007:1984];
    filter_input_0_1 = buffer_data_2[2007:1984];
    filter_input_0_2 = blur3x3_dout[2007:1984];
    current_RowCol_0 = {img_addr, 10'd249};
  end
  else if (detected_keypoint[0][249]) begin
    filter_input_0_0 = buffer_data_3[2015:1992];
    filter_input_0_1 = buffer_data_2[2015:1992];
    filter_input_0_2 = blur3x3_dout[2015:1992];
    current_RowCol_0 = {img_addr, 10'd250};
  end
  else if (detected_keypoint[0][250]) begin
    filter_input_0_0 = buffer_data_3[2023:2000];
    filter_input_0_1 = buffer_data_2[2023:2000];
    filter_input_0_2 = blur3x3_dout[2023:2000];
    current_RowCol_0 = {img_addr, 10'd251};
  end
  else if (detected_keypoint[0][251]) begin
    filter_input_0_0 = buffer_data_3[2031:2008];
    filter_input_0_1 = buffer_data_2[2031:2008];
    filter_input_0_2 = blur3x3_dout[2031:2008];
    current_RowCol_0 = {img_addr, 10'd252};
  end
  else if (detected_keypoint[0][252]) begin
    filter_input_0_0 = buffer_data_3[2039:2016];
    filter_input_0_1 = buffer_data_2[2039:2016];
    filter_input_0_2 = blur3x3_dout[2039:2016];
    current_RowCol_0 = {img_addr, 10'd253};
  end
  else if (detected_keypoint[0][253]) begin
    filter_input_0_0 = buffer_data_3[2047:2024];
    filter_input_0_1 = buffer_data_2[2047:2024];
    filter_input_0_2 = blur3x3_dout[2047:2024];
    current_RowCol_0 = {img_addr, 10'd254};
  end
  else if (detected_keypoint[0][254]) begin
    filter_input_0_0 = buffer_data_3[2055:2032];
    filter_input_0_1 = buffer_data_2[2055:2032];
    filter_input_0_2 = blur3x3_dout[2055:2032];
    current_RowCol_0 = {img_addr, 10'd255};
  end
  else if (detected_keypoint[0][255]) begin
    filter_input_0_0 = buffer_data_3[2063:2040];
    filter_input_0_1 = buffer_data_2[2063:2040];
    filter_input_0_2 = blur3x3_dout[2063:2040];
    current_RowCol_0 = {img_addr, 10'd256};
  end
  else if (detected_keypoint[0][256]) begin
    filter_input_0_0 = buffer_data_3[2071:2048];
    filter_input_0_1 = buffer_data_2[2071:2048];
    filter_input_0_2 = blur3x3_dout[2071:2048];
    current_RowCol_0 = {img_addr, 10'd257};
  end
  else if (detected_keypoint[0][257]) begin
    filter_input_0_0 = buffer_data_3[2079:2056];
    filter_input_0_1 = buffer_data_2[2079:2056];
    filter_input_0_2 = blur3x3_dout[2079:2056];
    current_RowCol_0 = {img_addr, 10'd258};
  end
  else if (detected_keypoint[0][258]) begin
    filter_input_0_0 = buffer_data_3[2087:2064];
    filter_input_0_1 = buffer_data_2[2087:2064];
    filter_input_0_2 = blur3x3_dout[2087:2064];
    current_RowCol_0 = {img_addr, 10'd259};
  end
  else if (detected_keypoint[0][259]) begin
    filter_input_0_0 = buffer_data_3[2095:2072];
    filter_input_0_1 = buffer_data_2[2095:2072];
    filter_input_0_2 = blur3x3_dout[2095:2072];
    current_RowCol_0 = {img_addr, 10'd260};
  end
  else if (detected_keypoint[0][260]) begin
    filter_input_0_0 = buffer_data_3[2103:2080];
    filter_input_0_1 = buffer_data_2[2103:2080];
    filter_input_0_2 = blur3x3_dout[2103:2080];
    current_RowCol_0 = {img_addr, 10'd261};
  end
  else if (detected_keypoint[0][261]) begin
    filter_input_0_0 = buffer_data_3[2111:2088];
    filter_input_0_1 = buffer_data_2[2111:2088];
    filter_input_0_2 = blur3x3_dout[2111:2088];
    current_RowCol_0 = {img_addr, 10'd262};
  end
  else if (detected_keypoint[0][262]) begin
    filter_input_0_0 = buffer_data_3[2119:2096];
    filter_input_0_1 = buffer_data_2[2119:2096];
    filter_input_0_2 = blur3x3_dout[2119:2096];
    current_RowCol_0 = {img_addr, 10'd263};
  end
  else if (detected_keypoint[0][263]) begin
    filter_input_0_0 = buffer_data_3[2127:2104];
    filter_input_0_1 = buffer_data_2[2127:2104];
    filter_input_0_2 = blur3x3_dout[2127:2104];
    current_RowCol_0 = {img_addr, 10'd264};
  end
  else if (detected_keypoint[0][264]) begin
    filter_input_0_0 = buffer_data_3[2135:2112];
    filter_input_0_1 = buffer_data_2[2135:2112];
    filter_input_0_2 = blur3x3_dout[2135:2112];
    current_RowCol_0 = {img_addr, 10'd265};
  end
  else if (detected_keypoint[0][265]) begin
    filter_input_0_0 = buffer_data_3[2143:2120];
    filter_input_0_1 = buffer_data_2[2143:2120];
    filter_input_0_2 = blur3x3_dout[2143:2120];
    current_RowCol_0 = {img_addr, 10'd266};
  end
  else if (detected_keypoint[0][266]) begin
    filter_input_0_0 = buffer_data_3[2151:2128];
    filter_input_0_1 = buffer_data_2[2151:2128];
    filter_input_0_2 = blur3x3_dout[2151:2128];
    current_RowCol_0 = {img_addr, 10'd267};
  end
  else if (detected_keypoint[0][267]) begin
    filter_input_0_0 = buffer_data_3[2159:2136];
    filter_input_0_1 = buffer_data_2[2159:2136];
    filter_input_0_2 = blur3x3_dout[2159:2136];
    current_RowCol_0 = {img_addr, 10'd268};
  end
  else if (detected_keypoint[0][268]) begin
    filter_input_0_0 = buffer_data_3[2167:2144];
    filter_input_0_1 = buffer_data_2[2167:2144];
    filter_input_0_2 = blur3x3_dout[2167:2144];
    current_RowCol_0 = {img_addr, 10'd269};
  end
  else if (detected_keypoint[0][269]) begin
    filter_input_0_0 = buffer_data_3[2175:2152];
    filter_input_0_1 = buffer_data_2[2175:2152];
    filter_input_0_2 = blur3x3_dout[2175:2152];
    current_RowCol_0 = {img_addr, 10'd270};
  end
  else if (detected_keypoint[0][270]) begin
    filter_input_0_0 = buffer_data_3[2183:2160];
    filter_input_0_1 = buffer_data_2[2183:2160];
    filter_input_0_2 = blur3x3_dout[2183:2160];
    current_RowCol_0 = {img_addr, 10'd271};
  end
  else if (detected_keypoint[0][271]) begin
    filter_input_0_0 = buffer_data_3[2191:2168];
    filter_input_0_1 = buffer_data_2[2191:2168];
    filter_input_0_2 = blur3x3_dout[2191:2168];
    current_RowCol_0 = {img_addr, 10'd272};
  end
  else if (detected_keypoint[0][272]) begin
    filter_input_0_0 = buffer_data_3[2199:2176];
    filter_input_0_1 = buffer_data_2[2199:2176];
    filter_input_0_2 = blur3x3_dout[2199:2176];
    current_RowCol_0 = {img_addr, 10'd273};
  end
  else if (detected_keypoint[0][273]) begin
    filter_input_0_0 = buffer_data_3[2207:2184];
    filter_input_0_1 = buffer_data_2[2207:2184];
    filter_input_0_2 = blur3x3_dout[2207:2184];
    current_RowCol_0 = {img_addr, 10'd274};
  end
  else if (detected_keypoint[0][274]) begin
    filter_input_0_0 = buffer_data_3[2215:2192];
    filter_input_0_1 = buffer_data_2[2215:2192];
    filter_input_0_2 = blur3x3_dout[2215:2192];
    current_RowCol_0 = {img_addr, 10'd275};
  end
  else if (detected_keypoint[0][275]) begin
    filter_input_0_0 = buffer_data_3[2223:2200];
    filter_input_0_1 = buffer_data_2[2223:2200];
    filter_input_0_2 = blur3x3_dout[2223:2200];
    current_RowCol_0 = {img_addr, 10'd276};
  end
  else if (detected_keypoint[0][276]) begin
    filter_input_0_0 = buffer_data_3[2231:2208];
    filter_input_0_1 = buffer_data_2[2231:2208];
    filter_input_0_2 = blur3x3_dout[2231:2208];
    current_RowCol_0 = {img_addr, 10'd277};
  end
  else if (detected_keypoint[0][277]) begin
    filter_input_0_0 = buffer_data_3[2239:2216];
    filter_input_0_1 = buffer_data_2[2239:2216];
    filter_input_0_2 = blur3x3_dout[2239:2216];
    current_RowCol_0 = {img_addr, 10'd278};
  end
  else if (detected_keypoint[0][278]) begin
    filter_input_0_0 = buffer_data_3[2247:2224];
    filter_input_0_1 = buffer_data_2[2247:2224];
    filter_input_0_2 = blur3x3_dout[2247:2224];
    current_RowCol_0 = {img_addr, 10'd279};
  end
  else if (detected_keypoint[0][279]) begin
    filter_input_0_0 = buffer_data_3[2255:2232];
    filter_input_0_1 = buffer_data_2[2255:2232];
    filter_input_0_2 = blur3x3_dout[2255:2232];
    current_RowCol_0 = {img_addr, 10'd280};
  end
  else if (detected_keypoint[0][280]) begin
    filter_input_0_0 = buffer_data_3[2263:2240];
    filter_input_0_1 = buffer_data_2[2263:2240];
    filter_input_0_2 = blur3x3_dout[2263:2240];
    current_RowCol_0 = {img_addr, 10'd281};
  end
  else if (detected_keypoint[0][281]) begin
    filter_input_0_0 = buffer_data_3[2271:2248];
    filter_input_0_1 = buffer_data_2[2271:2248];
    filter_input_0_2 = blur3x3_dout[2271:2248];
    current_RowCol_0 = {img_addr, 10'd282};
  end
  else if (detected_keypoint[0][282]) begin
    filter_input_0_0 = buffer_data_3[2279:2256];
    filter_input_0_1 = buffer_data_2[2279:2256];
    filter_input_0_2 = blur3x3_dout[2279:2256];
    current_RowCol_0 = {img_addr, 10'd283};
  end
  else if (detected_keypoint[0][283]) begin
    filter_input_0_0 = buffer_data_3[2287:2264];
    filter_input_0_1 = buffer_data_2[2287:2264];
    filter_input_0_2 = blur3x3_dout[2287:2264];
    current_RowCol_0 = {img_addr, 10'd284};
  end
  else if (detected_keypoint[0][284]) begin
    filter_input_0_0 = buffer_data_3[2295:2272];
    filter_input_0_1 = buffer_data_2[2295:2272];
    filter_input_0_2 = blur3x3_dout[2295:2272];
    current_RowCol_0 = {img_addr, 10'd285};
  end
  else if (detected_keypoint[0][285]) begin
    filter_input_0_0 = buffer_data_3[2303:2280];
    filter_input_0_1 = buffer_data_2[2303:2280];
    filter_input_0_2 = blur3x3_dout[2303:2280];
    current_RowCol_0 = {img_addr, 10'd286};
  end
  else if (detected_keypoint[0][286]) begin
    filter_input_0_0 = buffer_data_3[2311:2288];
    filter_input_0_1 = buffer_data_2[2311:2288];
    filter_input_0_2 = blur3x3_dout[2311:2288];
    current_RowCol_0 = {img_addr, 10'd287};
  end
  else if (detected_keypoint[0][287]) begin
    filter_input_0_0 = buffer_data_3[2319:2296];
    filter_input_0_1 = buffer_data_2[2319:2296];
    filter_input_0_2 = blur3x3_dout[2319:2296];
    current_RowCol_0 = {img_addr, 10'd288};
  end
  else if (detected_keypoint[0][288]) begin
    filter_input_0_0 = buffer_data_3[2327:2304];
    filter_input_0_1 = buffer_data_2[2327:2304];
    filter_input_0_2 = blur3x3_dout[2327:2304];
    current_RowCol_0 = {img_addr, 10'd289};
  end
  else if (detected_keypoint[0][289]) begin
    filter_input_0_0 = buffer_data_3[2335:2312];
    filter_input_0_1 = buffer_data_2[2335:2312];
    filter_input_0_2 = blur3x3_dout[2335:2312];
    current_RowCol_0 = {img_addr, 10'd290};
  end
  else if (detected_keypoint[0][290]) begin
    filter_input_0_0 = buffer_data_3[2343:2320];
    filter_input_0_1 = buffer_data_2[2343:2320];
    filter_input_0_2 = blur3x3_dout[2343:2320];
    current_RowCol_0 = {img_addr, 10'd291};
  end
  else if (detected_keypoint[0][291]) begin
    filter_input_0_0 = buffer_data_3[2351:2328];
    filter_input_0_1 = buffer_data_2[2351:2328];
    filter_input_0_2 = blur3x3_dout[2351:2328];
    current_RowCol_0 = {img_addr, 10'd292};
  end
  else if (detected_keypoint[0][292]) begin
    filter_input_0_0 = buffer_data_3[2359:2336];
    filter_input_0_1 = buffer_data_2[2359:2336];
    filter_input_0_2 = blur3x3_dout[2359:2336];
    current_RowCol_0 = {img_addr, 10'd293};
  end
  else if (detected_keypoint[0][293]) begin
    filter_input_0_0 = buffer_data_3[2367:2344];
    filter_input_0_1 = buffer_data_2[2367:2344];
    filter_input_0_2 = blur3x3_dout[2367:2344];
    current_RowCol_0 = {img_addr, 10'd294};
  end
  else if (detected_keypoint[0][294]) begin
    filter_input_0_0 = buffer_data_3[2375:2352];
    filter_input_0_1 = buffer_data_2[2375:2352];
    filter_input_0_2 = blur3x3_dout[2375:2352];
    current_RowCol_0 = {img_addr, 10'd295};
  end
  else if (detected_keypoint[0][295]) begin
    filter_input_0_0 = buffer_data_3[2383:2360];
    filter_input_0_1 = buffer_data_2[2383:2360];
    filter_input_0_2 = blur3x3_dout[2383:2360];
    current_RowCol_0 = {img_addr, 10'd296};
  end
  else if (detected_keypoint[0][296]) begin
    filter_input_0_0 = buffer_data_3[2391:2368];
    filter_input_0_1 = buffer_data_2[2391:2368];
    filter_input_0_2 = blur3x3_dout[2391:2368];
    current_RowCol_0 = {img_addr, 10'd297};
  end
  else if (detected_keypoint[0][297]) begin
    filter_input_0_0 = buffer_data_3[2399:2376];
    filter_input_0_1 = buffer_data_2[2399:2376];
    filter_input_0_2 = blur3x3_dout[2399:2376];
    current_RowCol_0 = {img_addr, 10'd298};
  end
  else if (detected_keypoint[0][298]) begin
    filter_input_0_0 = buffer_data_3[2407:2384];
    filter_input_0_1 = buffer_data_2[2407:2384];
    filter_input_0_2 = blur3x3_dout[2407:2384];
    current_RowCol_0 = {img_addr, 10'd299};
  end
  else if (detected_keypoint[0][299]) begin
    filter_input_0_0 = buffer_data_3[2415:2392];
    filter_input_0_1 = buffer_data_2[2415:2392];
    filter_input_0_2 = blur3x3_dout[2415:2392];
    current_RowCol_0 = {img_addr, 10'd300};
  end
  else if (detected_keypoint[0][300]) begin
    filter_input_0_0 = buffer_data_3[2423:2400];
    filter_input_0_1 = buffer_data_2[2423:2400];
    filter_input_0_2 = blur3x3_dout[2423:2400];
    current_RowCol_0 = {img_addr, 10'd301};
  end
  else if (detected_keypoint[0][301]) begin
    filter_input_0_0 = buffer_data_3[2431:2408];
    filter_input_0_1 = buffer_data_2[2431:2408];
    filter_input_0_2 = blur3x3_dout[2431:2408];
    current_RowCol_0 = {img_addr, 10'd302};
  end
  else if (detected_keypoint[0][302]) begin
    filter_input_0_0 = buffer_data_3[2439:2416];
    filter_input_0_1 = buffer_data_2[2439:2416];
    filter_input_0_2 = blur3x3_dout[2439:2416];
    current_RowCol_0 = {img_addr, 10'd303};
  end
  else if (detected_keypoint[0][303]) begin
    filter_input_0_0 = buffer_data_3[2447:2424];
    filter_input_0_1 = buffer_data_2[2447:2424];
    filter_input_0_2 = blur3x3_dout[2447:2424];
    current_RowCol_0 = {img_addr, 10'd304};
  end
  else if (detected_keypoint[0][304]) begin
    filter_input_0_0 = buffer_data_3[2455:2432];
    filter_input_0_1 = buffer_data_2[2455:2432];
    filter_input_0_2 = blur3x3_dout[2455:2432];
    current_RowCol_0 = {img_addr, 10'd305};
  end
  else if (detected_keypoint[0][305]) begin
    filter_input_0_0 = buffer_data_3[2463:2440];
    filter_input_0_1 = buffer_data_2[2463:2440];
    filter_input_0_2 = blur3x3_dout[2463:2440];
    current_RowCol_0 = {img_addr, 10'd306};
  end
  else if (detected_keypoint[0][306]) begin
    filter_input_0_0 = buffer_data_3[2471:2448];
    filter_input_0_1 = buffer_data_2[2471:2448];
    filter_input_0_2 = blur3x3_dout[2471:2448];
    current_RowCol_0 = {img_addr, 10'd307};
  end
  else if (detected_keypoint[0][307]) begin
    filter_input_0_0 = buffer_data_3[2479:2456];
    filter_input_0_1 = buffer_data_2[2479:2456];
    filter_input_0_2 = blur3x3_dout[2479:2456];
    current_RowCol_0 = {img_addr, 10'd308};
  end
  else if (detected_keypoint[0][308]) begin
    filter_input_0_0 = buffer_data_3[2487:2464];
    filter_input_0_1 = buffer_data_2[2487:2464];
    filter_input_0_2 = blur3x3_dout[2487:2464];
    current_RowCol_0 = {img_addr, 10'd309};
  end
  else if (detected_keypoint[0][309]) begin
    filter_input_0_0 = buffer_data_3[2495:2472];
    filter_input_0_1 = buffer_data_2[2495:2472];
    filter_input_0_2 = blur3x3_dout[2495:2472];
    current_RowCol_0 = {img_addr, 10'd310};
  end
  else if (detected_keypoint[0][310]) begin
    filter_input_0_0 = buffer_data_3[2503:2480];
    filter_input_0_1 = buffer_data_2[2503:2480];
    filter_input_0_2 = blur3x3_dout[2503:2480];
    current_RowCol_0 = {img_addr, 10'd311};
  end
  else if (detected_keypoint[0][311]) begin
    filter_input_0_0 = buffer_data_3[2511:2488];
    filter_input_0_1 = buffer_data_2[2511:2488];
    filter_input_0_2 = blur3x3_dout[2511:2488];
    current_RowCol_0 = {img_addr, 10'd312};
  end
  else if (detected_keypoint[0][312]) begin
    filter_input_0_0 = buffer_data_3[2519:2496];
    filter_input_0_1 = buffer_data_2[2519:2496];
    filter_input_0_2 = blur3x3_dout[2519:2496];
    current_RowCol_0 = {img_addr, 10'd313};
  end
  else if (detected_keypoint[0][313]) begin
    filter_input_0_0 = buffer_data_3[2527:2504];
    filter_input_0_1 = buffer_data_2[2527:2504];
    filter_input_0_2 = blur3x3_dout[2527:2504];
    current_RowCol_0 = {img_addr, 10'd314};
  end
  else if (detected_keypoint[0][314]) begin
    filter_input_0_0 = buffer_data_3[2535:2512];
    filter_input_0_1 = buffer_data_2[2535:2512];
    filter_input_0_2 = blur3x3_dout[2535:2512];
    current_RowCol_0 = {img_addr, 10'd315};
  end
  else if (detected_keypoint[0][315]) begin
    filter_input_0_0 = buffer_data_3[2543:2520];
    filter_input_0_1 = buffer_data_2[2543:2520];
    filter_input_0_2 = blur3x3_dout[2543:2520];
    current_RowCol_0 = {img_addr, 10'd316};
  end
  else if (detected_keypoint[0][316]) begin
    filter_input_0_0 = buffer_data_3[2551:2528];
    filter_input_0_1 = buffer_data_2[2551:2528];
    filter_input_0_2 = blur3x3_dout[2551:2528];
    current_RowCol_0 = {img_addr, 10'd317};
  end
  else if (detected_keypoint[0][317]) begin
    filter_input_0_0 = buffer_data_3[2559:2536];
    filter_input_0_1 = buffer_data_2[2559:2536];
    filter_input_0_2 = blur3x3_dout[2559:2536];
    current_RowCol_0 = {img_addr, 10'd318};
  end
  else if (detected_keypoint[0][318]) begin
    filter_input_0_0 = buffer_data_3[2567:2544];
    filter_input_0_1 = buffer_data_2[2567:2544];
    filter_input_0_2 = blur3x3_dout[2567:2544];
    current_RowCol_0 = {img_addr, 10'd319};
  end
  else if (detected_keypoint[0][319]) begin
    filter_input_0_0 = buffer_data_3[2575:2552];
    filter_input_0_1 = buffer_data_2[2575:2552];
    filter_input_0_2 = blur3x3_dout[2575:2552];
    current_RowCol_0 = {img_addr, 10'd320};
  end
  else if (detected_keypoint[0][320]) begin
    filter_input_0_0 = buffer_data_3[2583:2560];
    filter_input_0_1 = buffer_data_2[2583:2560];
    filter_input_0_2 = blur3x3_dout[2583:2560];
    current_RowCol_0 = {img_addr, 10'd321};
  end
  else if (detected_keypoint[0][321]) begin
    filter_input_0_0 = buffer_data_3[2591:2568];
    filter_input_0_1 = buffer_data_2[2591:2568];
    filter_input_0_2 = blur3x3_dout[2591:2568];
    current_RowCol_0 = {img_addr, 10'd322};
  end
  else if (detected_keypoint[0][322]) begin
    filter_input_0_0 = buffer_data_3[2599:2576];
    filter_input_0_1 = buffer_data_2[2599:2576];
    filter_input_0_2 = blur3x3_dout[2599:2576];
    current_RowCol_0 = {img_addr, 10'd323};
  end
  else if (detected_keypoint[0][323]) begin
    filter_input_0_0 = buffer_data_3[2607:2584];
    filter_input_0_1 = buffer_data_2[2607:2584];
    filter_input_0_2 = blur3x3_dout[2607:2584];
    current_RowCol_0 = {img_addr, 10'd324};
  end
  else if (detected_keypoint[0][324]) begin
    filter_input_0_0 = buffer_data_3[2615:2592];
    filter_input_0_1 = buffer_data_2[2615:2592];
    filter_input_0_2 = blur3x3_dout[2615:2592];
    current_RowCol_0 = {img_addr, 10'd325};
  end
  else if (detected_keypoint[0][325]) begin
    filter_input_0_0 = buffer_data_3[2623:2600];
    filter_input_0_1 = buffer_data_2[2623:2600];
    filter_input_0_2 = blur3x3_dout[2623:2600];
    current_RowCol_0 = {img_addr, 10'd326};
  end
  else if (detected_keypoint[0][326]) begin
    filter_input_0_0 = buffer_data_3[2631:2608];
    filter_input_0_1 = buffer_data_2[2631:2608];
    filter_input_0_2 = blur3x3_dout[2631:2608];
    current_RowCol_0 = {img_addr, 10'd327};
  end
  else if (detected_keypoint[0][327]) begin
    filter_input_0_0 = buffer_data_3[2639:2616];
    filter_input_0_1 = buffer_data_2[2639:2616];
    filter_input_0_2 = blur3x3_dout[2639:2616];
    current_RowCol_0 = {img_addr, 10'd328};
  end
  else if (detected_keypoint[0][328]) begin
    filter_input_0_0 = buffer_data_3[2647:2624];
    filter_input_0_1 = buffer_data_2[2647:2624];
    filter_input_0_2 = blur3x3_dout[2647:2624];
    current_RowCol_0 = {img_addr, 10'd329};
  end
  else if (detected_keypoint[0][329]) begin
    filter_input_0_0 = buffer_data_3[2655:2632];
    filter_input_0_1 = buffer_data_2[2655:2632];
    filter_input_0_2 = blur3x3_dout[2655:2632];
    current_RowCol_0 = {img_addr, 10'd330};
  end
  else if (detected_keypoint[0][330]) begin
    filter_input_0_0 = buffer_data_3[2663:2640];
    filter_input_0_1 = buffer_data_2[2663:2640];
    filter_input_0_2 = blur3x3_dout[2663:2640];
    current_RowCol_0 = {img_addr, 10'd331};
  end
  else if (detected_keypoint[0][331]) begin
    filter_input_0_0 = buffer_data_3[2671:2648];
    filter_input_0_1 = buffer_data_2[2671:2648];
    filter_input_0_2 = blur3x3_dout[2671:2648];
    current_RowCol_0 = {img_addr, 10'd332};
  end
  else if (detected_keypoint[0][332]) begin
    filter_input_0_0 = buffer_data_3[2679:2656];
    filter_input_0_1 = buffer_data_2[2679:2656];
    filter_input_0_2 = blur3x3_dout[2679:2656];
    current_RowCol_0 = {img_addr, 10'd333};
  end
  else if (detected_keypoint[0][333]) begin
    filter_input_0_0 = buffer_data_3[2687:2664];
    filter_input_0_1 = buffer_data_2[2687:2664];
    filter_input_0_2 = blur3x3_dout[2687:2664];
    current_RowCol_0 = {img_addr, 10'd334};
  end
  else if (detected_keypoint[0][334]) begin
    filter_input_0_0 = buffer_data_3[2695:2672];
    filter_input_0_1 = buffer_data_2[2695:2672];
    filter_input_0_2 = blur3x3_dout[2695:2672];
    current_RowCol_0 = {img_addr, 10'd335};
  end
  else if (detected_keypoint[0][335]) begin
    filter_input_0_0 = buffer_data_3[2703:2680];
    filter_input_0_1 = buffer_data_2[2703:2680];
    filter_input_0_2 = blur3x3_dout[2703:2680];
    current_RowCol_0 = {img_addr, 10'd336};
  end
  else if (detected_keypoint[0][336]) begin
    filter_input_0_0 = buffer_data_3[2711:2688];
    filter_input_0_1 = buffer_data_2[2711:2688];
    filter_input_0_2 = blur3x3_dout[2711:2688];
    current_RowCol_0 = {img_addr, 10'd337};
  end
  else if (detected_keypoint[0][337]) begin
    filter_input_0_0 = buffer_data_3[2719:2696];
    filter_input_0_1 = buffer_data_2[2719:2696];
    filter_input_0_2 = blur3x3_dout[2719:2696];
    current_RowCol_0 = {img_addr, 10'd338};
  end
  else if (detected_keypoint[0][338]) begin
    filter_input_0_0 = buffer_data_3[2727:2704];
    filter_input_0_1 = buffer_data_2[2727:2704];
    filter_input_0_2 = blur3x3_dout[2727:2704];
    current_RowCol_0 = {img_addr, 10'd339};
  end
  else if (detected_keypoint[0][339]) begin
    filter_input_0_0 = buffer_data_3[2735:2712];
    filter_input_0_1 = buffer_data_2[2735:2712];
    filter_input_0_2 = blur3x3_dout[2735:2712];
    current_RowCol_0 = {img_addr, 10'd340};
  end
  else if (detected_keypoint[0][340]) begin
    filter_input_0_0 = buffer_data_3[2743:2720];
    filter_input_0_1 = buffer_data_2[2743:2720];
    filter_input_0_2 = blur3x3_dout[2743:2720];
    current_RowCol_0 = {img_addr, 10'd341};
  end
  else if (detected_keypoint[0][341]) begin
    filter_input_0_0 = buffer_data_3[2751:2728];
    filter_input_0_1 = buffer_data_2[2751:2728];
    filter_input_0_2 = blur3x3_dout[2751:2728];
    current_RowCol_0 = {img_addr, 10'd342};
  end
  else if (detected_keypoint[0][342]) begin
    filter_input_0_0 = buffer_data_3[2759:2736];
    filter_input_0_1 = buffer_data_2[2759:2736];
    filter_input_0_2 = blur3x3_dout[2759:2736];
    current_RowCol_0 = {img_addr, 10'd343};
  end
  else if (detected_keypoint[0][343]) begin
    filter_input_0_0 = buffer_data_3[2767:2744];
    filter_input_0_1 = buffer_data_2[2767:2744];
    filter_input_0_2 = blur3x3_dout[2767:2744];
    current_RowCol_0 = {img_addr, 10'd344};
  end
  else if (detected_keypoint[0][344]) begin
    filter_input_0_0 = buffer_data_3[2775:2752];
    filter_input_0_1 = buffer_data_2[2775:2752];
    filter_input_0_2 = blur3x3_dout[2775:2752];
    current_RowCol_0 = {img_addr, 10'd345};
  end
  else if (detected_keypoint[0][345]) begin
    filter_input_0_0 = buffer_data_3[2783:2760];
    filter_input_0_1 = buffer_data_2[2783:2760];
    filter_input_0_2 = blur3x3_dout[2783:2760];
    current_RowCol_0 = {img_addr, 10'd346};
  end
  else if (detected_keypoint[0][346]) begin
    filter_input_0_0 = buffer_data_3[2791:2768];
    filter_input_0_1 = buffer_data_2[2791:2768];
    filter_input_0_2 = blur3x3_dout[2791:2768];
    current_RowCol_0 = {img_addr, 10'd347};
  end
  else if (detected_keypoint[0][347]) begin
    filter_input_0_0 = buffer_data_3[2799:2776];
    filter_input_0_1 = buffer_data_2[2799:2776];
    filter_input_0_2 = blur3x3_dout[2799:2776];
    current_RowCol_0 = {img_addr, 10'd348};
  end
  else if (detected_keypoint[0][348]) begin
    filter_input_0_0 = buffer_data_3[2807:2784];
    filter_input_0_1 = buffer_data_2[2807:2784];
    filter_input_0_2 = blur3x3_dout[2807:2784];
    current_RowCol_0 = {img_addr, 10'd349};
  end
  else if (detected_keypoint[0][349]) begin
    filter_input_0_0 = buffer_data_3[2815:2792];
    filter_input_0_1 = buffer_data_2[2815:2792];
    filter_input_0_2 = blur3x3_dout[2815:2792];
    current_RowCol_0 = {img_addr, 10'd350};
  end
  else if (detected_keypoint[0][350]) begin
    filter_input_0_0 = buffer_data_3[2823:2800];
    filter_input_0_1 = buffer_data_2[2823:2800];
    filter_input_0_2 = blur3x3_dout[2823:2800];
    current_RowCol_0 = {img_addr, 10'd351};
  end
  else if (detected_keypoint[0][351]) begin
    filter_input_0_0 = buffer_data_3[2831:2808];
    filter_input_0_1 = buffer_data_2[2831:2808];
    filter_input_0_2 = blur3x3_dout[2831:2808];
    current_RowCol_0 = {img_addr, 10'd352};
  end
  else if (detected_keypoint[0][352]) begin
    filter_input_0_0 = buffer_data_3[2839:2816];
    filter_input_0_1 = buffer_data_2[2839:2816];
    filter_input_0_2 = blur3x3_dout[2839:2816];
    current_RowCol_0 = {img_addr, 10'd353};
  end
  else if (detected_keypoint[0][353]) begin
    filter_input_0_0 = buffer_data_3[2847:2824];
    filter_input_0_1 = buffer_data_2[2847:2824];
    filter_input_0_2 = blur3x3_dout[2847:2824];
    current_RowCol_0 = {img_addr, 10'd354};
  end
  else if (detected_keypoint[0][354]) begin
    filter_input_0_0 = buffer_data_3[2855:2832];
    filter_input_0_1 = buffer_data_2[2855:2832];
    filter_input_0_2 = blur3x3_dout[2855:2832];
    current_RowCol_0 = {img_addr, 10'd355};
  end
  else if (detected_keypoint[0][355]) begin
    filter_input_0_0 = buffer_data_3[2863:2840];
    filter_input_0_1 = buffer_data_2[2863:2840];
    filter_input_0_2 = blur3x3_dout[2863:2840];
    current_RowCol_0 = {img_addr, 10'd356};
  end
  else if (detected_keypoint[0][356]) begin
    filter_input_0_0 = buffer_data_3[2871:2848];
    filter_input_0_1 = buffer_data_2[2871:2848];
    filter_input_0_2 = blur3x3_dout[2871:2848];
    current_RowCol_0 = {img_addr, 10'd357};
  end
  else if (detected_keypoint[0][357]) begin
    filter_input_0_0 = buffer_data_3[2879:2856];
    filter_input_0_1 = buffer_data_2[2879:2856];
    filter_input_0_2 = blur3x3_dout[2879:2856];
    current_RowCol_0 = {img_addr, 10'd358};
  end
  else if (detected_keypoint[0][358]) begin
    filter_input_0_0 = buffer_data_3[2887:2864];
    filter_input_0_1 = buffer_data_2[2887:2864];
    filter_input_0_2 = blur3x3_dout[2887:2864];
    current_RowCol_0 = {img_addr, 10'd359};
  end
  else if (detected_keypoint[0][359]) begin
    filter_input_0_0 = buffer_data_3[2895:2872];
    filter_input_0_1 = buffer_data_2[2895:2872];
    filter_input_0_2 = blur3x3_dout[2895:2872];
    current_RowCol_0 = {img_addr, 10'd360};
  end
  else if (detected_keypoint[0][360]) begin
    filter_input_0_0 = buffer_data_3[2903:2880];
    filter_input_0_1 = buffer_data_2[2903:2880];
    filter_input_0_2 = blur3x3_dout[2903:2880];
    current_RowCol_0 = {img_addr, 10'd361};
  end
  else if (detected_keypoint[0][361]) begin
    filter_input_0_0 = buffer_data_3[2911:2888];
    filter_input_0_1 = buffer_data_2[2911:2888];
    filter_input_0_2 = blur3x3_dout[2911:2888];
    current_RowCol_0 = {img_addr, 10'd362};
  end
  else if (detected_keypoint[0][362]) begin
    filter_input_0_0 = buffer_data_3[2919:2896];
    filter_input_0_1 = buffer_data_2[2919:2896];
    filter_input_0_2 = blur3x3_dout[2919:2896];
    current_RowCol_0 = {img_addr, 10'd363};
  end
  else if (detected_keypoint[0][363]) begin
    filter_input_0_0 = buffer_data_3[2927:2904];
    filter_input_0_1 = buffer_data_2[2927:2904];
    filter_input_0_2 = blur3x3_dout[2927:2904];
    current_RowCol_0 = {img_addr, 10'd364};
  end
  else if (detected_keypoint[0][364]) begin
    filter_input_0_0 = buffer_data_3[2935:2912];
    filter_input_0_1 = buffer_data_2[2935:2912];
    filter_input_0_2 = blur3x3_dout[2935:2912];
    current_RowCol_0 = {img_addr, 10'd365};
  end
  else if (detected_keypoint[0][365]) begin
    filter_input_0_0 = buffer_data_3[2943:2920];
    filter_input_0_1 = buffer_data_2[2943:2920];
    filter_input_0_2 = blur3x3_dout[2943:2920];
    current_RowCol_0 = {img_addr, 10'd366};
  end
  else if (detected_keypoint[0][366]) begin
    filter_input_0_0 = buffer_data_3[2951:2928];
    filter_input_0_1 = buffer_data_2[2951:2928];
    filter_input_0_2 = blur3x3_dout[2951:2928];
    current_RowCol_0 = {img_addr, 10'd367};
  end
  else if (detected_keypoint[0][367]) begin
    filter_input_0_0 = buffer_data_3[2959:2936];
    filter_input_0_1 = buffer_data_2[2959:2936];
    filter_input_0_2 = blur3x3_dout[2959:2936];
    current_RowCol_0 = {img_addr, 10'd368};
  end
  else if (detected_keypoint[0][368]) begin
    filter_input_0_0 = buffer_data_3[2967:2944];
    filter_input_0_1 = buffer_data_2[2967:2944];
    filter_input_0_2 = blur3x3_dout[2967:2944];
    current_RowCol_0 = {img_addr, 10'd369};
  end
  else if (detected_keypoint[0][369]) begin
    filter_input_0_0 = buffer_data_3[2975:2952];
    filter_input_0_1 = buffer_data_2[2975:2952];
    filter_input_0_2 = blur3x3_dout[2975:2952];
    current_RowCol_0 = {img_addr, 10'd370};
  end
  else if (detected_keypoint[0][370]) begin
    filter_input_0_0 = buffer_data_3[2983:2960];
    filter_input_0_1 = buffer_data_2[2983:2960];
    filter_input_0_2 = blur3x3_dout[2983:2960];
    current_RowCol_0 = {img_addr, 10'd371};
  end
  else if (detected_keypoint[0][371]) begin
    filter_input_0_0 = buffer_data_3[2991:2968];
    filter_input_0_1 = buffer_data_2[2991:2968];
    filter_input_0_2 = blur3x3_dout[2991:2968];
    current_RowCol_0 = {img_addr, 10'd372};
  end
  else if (detected_keypoint[0][372]) begin
    filter_input_0_0 = buffer_data_3[2999:2976];
    filter_input_0_1 = buffer_data_2[2999:2976];
    filter_input_0_2 = blur3x3_dout[2999:2976];
    current_RowCol_0 = {img_addr, 10'd373};
  end
  else if (detected_keypoint[0][373]) begin
    filter_input_0_0 = buffer_data_3[3007:2984];
    filter_input_0_1 = buffer_data_2[3007:2984];
    filter_input_0_2 = blur3x3_dout[3007:2984];
    current_RowCol_0 = {img_addr, 10'd374};
  end
  else if (detected_keypoint[0][374]) begin
    filter_input_0_0 = buffer_data_3[3015:2992];
    filter_input_0_1 = buffer_data_2[3015:2992];
    filter_input_0_2 = blur3x3_dout[3015:2992];
    current_RowCol_0 = {img_addr, 10'd375};
  end
  else if (detected_keypoint[0][375]) begin
    filter_input_0_0 = buffer_data_3[3023:3000];
    filter_input_0_1 = buffer_data_2[3023:3000];
    filter_input_0_2 = blur3x3_dout[3023:3000];
    current_RowCol_0 = {img_addr, 10'd376};
  end
  else if (detected_keypoint[0][376]) begin
    filter_input_0_0 = buffer_data_3[3031:3008];
    filter_input_0_1 = buffer_data_2[3031:3008];
    filter_input_0_2 = blur3x3_dout[3031:3008];
    current_RowCol_0 = {img_addr, 10'd377};
  end
  else if (detected_keypoint[0][377]) begin
    filter_input_0_0 = buffer_data_3[3039:3016];
    filter_input_0_1 = buffer_data_2[3039:3016];
    filter_input_0_2 = blur3x3_dout[3039:3016];
    current_RowCol_0 = {img_addr, 10'd378};
  end
  else if (detected_keypoint[0][378]) begin
    filter_input_0_0 = buffer_data_3[3047:3024];
    filter_input_0_1 = buffer_data_2[3047:3024];
    filter_input_0_2 = blur3x3_dout[3047:3024];
    current_RowCol_0 = {img_addr, 10'd379};
  end
  else if (detected_keypoint[0][379]) begin
    filter_input_0_0 = buffer_data_3[3055:3032];
    filter_input_0_1 = buffer_data_2[3055:3032];
    filter_input_0_2 = blur3x3_dout[3055:3032];
    current_RowCol_0 = {img_addr, 10'd380};
  end
  else if (detected_keypoint[0][380]) begin
    filter_input_0_0 = buffer_data_3[3063:3040];
    filter_input_0_1 = buffer_data_2[3063:3040];
    filter_input_0_2 = blur3x3_dout[3063:3040];
    current_RowCol_0 = {img_addr, 10'd381};
  end
  else if (detected_keypoint[0][381]) begin
    filter_input_0_0 = buffer_data_3[3071:3048];
    filter_input_0_1 = buffer_data_2[3071:3048];
    filter_input_0_2 = blur3x3_dout[3071:3048];
    current_RowCol_0 = {img_addr, 10'd382};
  end
  else if (detected_keypoint[0][382]) begin
    filter_input_0_0 = buffer_data_3[3079:3056];
    filter_input_0_1 = buffer_data_2[3079:3056];
    filter_input_0_2 = blur3x3_dout[3079:3056];
    current_RowCol_0 = {img_addr, 10'd383};
  end
  else if (detected_keypoint[0][383]) begin
    filter_input_0_0 = buffer_data_3[3087:3064];
    filter_input_0_1 = buffer_data_2[3087:3064];
    filter_input_0_2 = blur3x3_dout[3087:3064];
    current_RowCol_0 = {img_addr, 10'd384};
  end
  else if (detected_keypoint[0][384]) begin
    filter_input_0_0 = buffer_data_3[3095:3072];
    filter_input_0_1 = buffer_data_2[3095:3072];
    filter_input_0_2 = blur3x3_dout[3095:3072];
    current_RowCol_0 = {img_addr, 10'd385};
  end
  else if (detected_keypoint[0][385]) begin
    filter_input_0_0 = buffer_data_3[3103:3080];
    filter_input_0_1 = buffer_data_2[3103:3080];
    filter_input_0_2 = blur3x3_dout[3103:3080];
    current_RowCol_0 = {img_addr, 10'd386};
  end
  else if (detected_keypoint[0][386]) begin
    filter_input_0_0 = buffer_data_3[3111:3088];
    filter_input_0_1 = buffer_data_2[3111:3088];
    filter_input_0_2 = blur3x3_dout[3111:3088];
    current_RowCol_0 = {img_addr, 10'd387};
  end
  else if (detected_keypoint[0][387]) begin
    filter_input_0_0 = buffer_data_3[3119:3096];
    filter_input_0_1 = buffer_data_2[3119:3096];
    filter_input_0_2 = blur3x3_dout[3119:3096];
    current_RowCol_0 = {img_addr, 10'd388};
  end
  else if (detected_keypoint[0][388]) begin
    filter_input_0_0 = buffer_data_3[3127:3104];
    filter_input_0_1 = buffer_data_2[3127:3104];
    filter_input_0_2 = blur3x3_dout[3127:3104];
    current_RowCol_0 = {img_addr, 10'd389};
  end
  else if (detected_keypoint[0][389]) begin
    filter_input_0_0 = buffer_data_3[3135:3112];
    filter_input_0_1 = buffer_data_2[3135:3112];
    filter_input_0_2 = blur3x3_dout[3135:3112];
    current_RowCol_0 = {img_addr, 10'd390};
  end
  else if (detected_keypoint[0][390]) begin
    filter_input_0_0 = buffer_data_3[3143:3120];
    filter_input_0_1 = buffer_data_2[3143:3120];
    filter_input_0_2 = blur3x3_dout[3143:3120];
    current_RowCol_0 = {img_addr, 10'd391};
  end
  else if (detected_keypoint[0][391]) begin
    filter_input_0_0 = buffer_data_3[3151:3128];
    filter_input_0_1 = buffer_data_2[3151:3128];
    filter_input_0_2 = blur3x3_dout[3151:3128];
    current_RowCol_0 = {img_addr, 10'd392};
  end
  else if (detected_keypoint[0][392]) begin
    filter_input_0_0 = buffer_data_3[3159:3136];
    filter_input_0_1 = buffer_data_2[3159:3136];
    filter_input_0_2 = blur3x3_dout[3159:3136];
    current_RowCol_0 = {img_addr, 10'd393};
  end
  else if (detected_keypoint[0][393]) begin
    filter_input_0_0 = buffer_data_3[3167:3144];
    filter_input_0_1 = buffer_data_2[3167:3144];
    filter_input_0_2 = blur3x3_dout[3167:3144];
    current_RowCol_0 = {img_addr, 10'd394};
  end
  else if (detected_keypoint[0][394]) begin
    filter_input_0_0 = buffer_data_3[3175:3152];
    filter_input_0_1 = buffer_data_2[3175:3152];
    filter_input_0_2 = blur3x3_dout[3175:3152];
    current_RowCol_0 = {img_addr, 10'd395};
  end
  else if (detected_keypoint[0][395]) begin
    filter_input_0_0 = buffer_data_3[3183:3160];
    filter_input_0_1 = buffer_data_2[3183:3160];
    filter_input_0_2 = blur3x3_dout[3183:3160];
    current_RowCol_0 = {img_addr, 10'd396};
  end
  else if (detected_keypoint[0][396]) begin
    filter_input_0_0 = buffer_data_3[3191:3168];
    filter_input_0_1 = buffer_data_2[3191:3168];
    filter_input_0_2 = blur3x3_dout[3191:3168];
    current_RowCol_0 = {img_addr, 10'd397};
  end
  else if (detected_keypoint[0][397]) begin
    filter_input_0_0 = buffer_data_3[3199:3176];
    filter_input_0_1 = buffer_data_2[3199:3176];
    filter_input_0_2 = blur3x3_dout[3199:3176];
    current_RowCol_0 = {img_addr, 10'd398};
  end
  else if (detected_keypoint[0][398]) begin
    filter_input_0_0 = buffer_data_3[3207:3184];
    filter_input_0_1 = buffer_data_2[3207:3184];
    filter_input_0_2 = blur3x3_dout[3207:3184];
    current_RowCol_0 = {img_addr, 10'd399};
  end
  else if (detected_keypoint[0][399]) begin
    filter_input_0_0 = buffer_data_3[3215:3192];
    filter_input_0_1 = buffer_data_2[3215:3192];
    filter_input_0_2 = blur3x3_dout[3215:3192];
    current_RowCol_0 = {img_addr, 10'd400};
  end
  else if (detected_keypoint[0][400]) begin
    filter_input_0_0 = buffer_data_3[3223:3200];
    filter_input_0_1 = buffer_data_2[3223:3200];
    filter_input_0_2 = blur3x3_dout[3223:3200];
    current_RowCol_0 = {img_addr, 10'd401};
  end
  else if (detected_keypoint[0][401]) begin
    filter_input_0_0 = buffer_data_3[3231:3208];
    filter_input_0_1 = buffer_data_2[3231:3208];
    filter_input_0_2 = blur3x3_dout[3231:3208];
    current_RowCol_0 = {img_addr, 10'd402};
  end
  else if (detected_keypoint[0][402]) begin
    filter_input_0_0 = buffer_data_3[3239:3216];
    filter_input_0_1 = buffer_data_2[3239:3216];
    filter_input_0_2 = blur3x3_dout[3239:3216];
    current_RowCol_0 = {img_addr, 10'd403};
  end
  else if (detected_keypoint[0][403]) begin
    filter_input_0_0 = buffer_data_3[3247:3224];
    filter_input_0_1 = buffer_data_2[3247:3224];
    filter_input_0_2 = blur3x3_dout[3247:3224];
    current_RowCol_0 = {img_addr, 10'd404};
  end
  else if (detected_keypoint[0][404]) begin
    filter_input_0_0 = buffer_data_3[3255:3232];
    filter_input_0_1 = buffer_data_2[3255:3232];
    filter_input_0_2 = blur3x3_dout[3255:3232];
    current_RowCol_0 = {img_addr, 10'd405};
  end
  else if (detected_keypoint[0][405]) begin
    filter_input_0_0 = buffer_data_3[3263:3240];
    filter_input_0_1 = buffer_data_2[3263:3240];
    filter_input_0_2 = blur3x3_dout[3263:3240];
    current_RowCol_0 = {img_addr, 10'd406};
  end
  else if (detected_keypoint[0][406]) begin
    filter_input_0_0 = buffer_data_3[3271:3248];
    filter_input_0_1 = buffer_data_2[3271:3248];
    filter_input_0_2 = blur3x3_dout[3271:3248];
    current_RowCol_0 = {img_addr, 10'd407};
  end
  else if (detected_keypoint[0][407]) begin
    filter_input_0_0 = buffer_data_3[3279:3256];
    filter_input_0_1 = buffer_data_2[3279:3256];
    filter_input_0_2 = blur3x3_dout[3279:3256];
    current_RowCol_0 = {img_addr, 10'd408};
  end
  else if (detected_keypoint[0][408]) begin
    filter_input_0_0 = buffer_data_3[3287:3264];
    filter_input_0_1 = buffer_data_2[3287:3264];
    filter_input_0_2 = blur3x3_dout[3287:3264];
    current_RowCol_0 = {img_addr, 10'd409};
  end
  else if (detected_keypoint[0][409]) begin
    filter_input_0_0 = buffer_data_3[3295:3272];
    filter_input_0_1 = buffer_data_2[3295:3272];
    filter_input_0_2 = blur3x3_dout[3295:3272];
    current_RowCol_0 = {img_addr, 10'd410};
  end
  else if (detected_keypoint[0][410]) begin
    filter_input_0_0 = buffer_data_3[3303:3280];
    filter_input_0_1 = buffer_data_2[3303:3280];
    filter_input_0_2 = blur3x3_dout[3303:3280];
    current_RowCol_0 = {img_addr, 10'd411};
  end
  else if (detected_keypoint[0][411]) begin
    filter_input_0_0 = buffer_data_3[3311:3288];
    filter_input_0_1 = buffer_data_2[3311:3288];
    filter_input_0_2 = blur3x3_dout[3311:3288];
    current_RowCol_0 = {img_addr, 10'd412};
  end
  else if (detected_keypoint[0][412]) begin
    filter_input_0_0 = buffer_data_3[3319:3296];
    filter_input_0_1 = buffer_data_2[3319:3296];
    filter_input_0_2 = blur3x3_dout[3319:3296];
    current_RowCol_0 = {img_addr, 10'd413};
  end
  else if (detected_keypoint[0][413]) begin
    filter_input_0_0 = buffer_data_3[3327:3304];
    filter_input_0_1 = buffer_data_2[3327:3304];
    filter_input_0_2 = blur3x3_dout[3327:3304];
    current_RowCol_0 = {img_addr, 10'd414};
  end
  else if (detected_keypoint[0][414]) begin
    filter_input_0_0 = buffer_data_3[3335:3312];
    filter_input_0_1 = buffer_data_2[3335:3312];
    filter_input_0_2 = blur3x3_dout[3335:3312];
    current_RowCol_0 = {img_addr, 10'd415};
  end
  else if (detected_keypoint[0][415]) begin
    filter_input_0_0 = buffer_data_3[3343:3320];
    filter_input_0_1 = buffer_data_2[3343:3320];
    filter_input_0_2 = blur3x3_dout[3343:3320];
    current_RowCol_0 = {img_addr, 10'd416};
  end
  else if (detected_keypoint[0][416]) begin
    filter_input_0_0 = buffer_data_3[3351:3328];
    filter_input_0_1 = buffer_data_2[3351:3328];
    filter_input_0_2 = blur3x3_dout[3351:3328];
    current_RowCol_0 = {img_addr, 10'd417};
  end
  else if (detected_keypoint[0][417]) begin
    filter_input_0_0 = buffer_data_3[3359:3336];
    filter_input_0_1 = buffer_data_2[3359:3336];
    filter_input_0_2 = blur3x3_dout[3359:3336];
    current_RowCol_0 = {img_addr, 10'd418};
  end
  else if (detected_keypoint[0][418]) begin
    filter_input_0_0 = buffer_data_3[3367:3344];
    filter_input_0_1 = buffer_data_2[3367:3344];
    filter_input_0_2 = blur3x3_dout[3367:3344];
    current_RowCol_0 = {img_addr, 10'd419};
  end
  else if (detected_keypoint[0][419]) begin
    filter_input_0_0 = buffer_data_3[3375:3352];
    filter_input_0_1 = buffer_data_2[3375:3352];
    filter_input_0_2 = blur3x3_dout[3375:3352];
    current_RowCol_0 = {img_addr, 10'd420};
  end
  else if (detected_keypoint[0][420]) begin
    filter_input_0_0 = buffer_data_3[3383:3360];
    filter_input_0_1 = buffer_data_2[3383:3360];
    filter_input_0_2 = blur3x3_dout[3383:3360];
    current_RowCol_0 = {img_addr, 10'd421};
  end
  else if (detected_keypoint[0][421]) begin
    filter_input_0_0 = buffer_data_3[3391:3368];
    filter_input_0_1 = buffer_data_2[3391:3368];
    filter_input_0_2 = blur3x3_dout[3391:3368];
    current_RowCol_0 = {img_addr, 10'd422};
  end
  else if (detected_keypoint[0][422]) begin
    filter_input_0_0 = buffer_data_3[3399:3376];
    filter_input_0_1 = buffer_data_2[3399:3376];
    filter_input_0_2 = blur3x3_dout[3399:3376];
    current_RowCol_0 = {img_addr, 10'd423};
  end
  else if (detected_keypoint[0][423]) begin
    filter_input_0_0 = buffer_data_3[3407:3384];
    filter_input_0_1 = buffer_data_2[3407:3384];
    filter_input_0_2 = blur3x3_dout[3407:3384];
    current_RowCol_0 = {img_addr, 10'd424};
  end
  else if (detected_keypoint[0][424]) begin
    filter_input_0_0 = buffer_data_3[3415:3392];
    filter_input_0_1 = buffer_data_2[3415:3392];
    filter_input_0_2 = blur3x3_dout[3415:3392];
    current_RowCol_0 = {img_addr, 10'd425};
  end
  else if (detected_keypoint[0][425]) begin
    filter_input_0_0 = buffer_data_3[3423:3400];
    filter_input_0_1 = buffer_data_2[3423:3400];
    filter_input_0_2 = blur3x3_dout[3423:3400];
    current_RowCol_0 = {img_addr, 10'd426};
  end
  else if (detected_keypoint[0][426]) begin
    filter_input_0_0 = buffer_data_3[3431:3408];
    filter_input_0_1 = buffer_data_2[3431:3408];
    filter_input_0_2 = blur3x3_dout[3431:3408];
    current_RowCol_0 = {img_addr, 10'd427};
  end
  else if (detected_keypoint[0][427]) begin
    filter_input_0_0 = buffer_data_3[3439:3416];
    filter_input_0_1 = buffer_data_2[3439:3416];
    filter_input_0_2 = blur3x3_dout[3439:3416];
    current_RowCol_0 = {img_addr, 10'd428};
  end
  else if (detected_keypoint[0][428]) begin
    filter_input_0_0 = buffer_data_3[3447:3424];
    filter_input_0_1 = buffer_data_2[3447:3424];
    filter_input_0_2 = blur3x3_dout[3447:3424];
    current_RowCol_0 = {img_addr, 10'd429};
  end
  else if (detected_keypoint[0][429]) begin
    filter_input_0_0 = buffer_data_3[3455:3432];
    filter_input_0_1 = buffer_data_2[3455:3432];
    filter_input_0_2 = blur3x3_dout[3455:3432];
    current_RowCol_0 = {img_addr, 10'd430};
  end
  else if (detected_keypoint[0][430]) begin
    filter_input_0_0 = buffer_data_3[3463:3440];
    filter_input_0_1 = buffer_data_2[3463:3440];
    filter_input_0_2 = blur3x3_dout[3463:3440];
    current_RowCol_0 = {img_addr, 10'd431};
  end
  else if (detected_keypoint[0][431]) begin
    filter_input_0_0 = buffer_data_3[3471:3448];
    filter_input_0_1 = buffer_data_2[3471:3448];
    filter_input_0_2 = blur3x3_dout[3471:3448];
    current_RowCol_0 = {img_addr, 10'd432};
  end
  else if (detected_keypoint[0][432]) begin
    filter_input_0_0 = buffer_data_3[3479:3456];
    filter_input_0_1 = buffer_data_2[3479:3456];
    filter_input_0_2 = blur3x3_dout[3479:3456];
    current_RowCol_0 = {img_addr, 10'd433};
  end
  else if (detected_keypoint[0][433]) begin
    filter_input_0_0 = buffer_data_3[3487:3464];
    filter_input_0_1 = buffer_data_2[3487:3464];
    filter_input_0_2 = blur3x3_dout[3487:3464];
    current_RowCol_0 = {img_addr, 10'd434};
  end
  else if (detected_keypoint[0][434]) begin
    filter_input_0_0 = buffer_data_3[3495:3472];
    filter_input_0_1 = buffer_data_2[3495:3472];
    filter_input_0_2 = blur3x3_dout[3495:3472];
    current_RowCol_0 = {img_addr, 10'd435};
  end
  else if (detected_keypoint[0][435]) begin
    filter_input_0_0 = buffer_data_3[3503:3480];
    filter_input_0_1 = buffer_data_2[3503:3480];
    filter_input_0_2 = blur3x3_dout[3503:3480];
    current_RowCol_0 = {img_addr, 10'd436};
  end
  else if (detected_keypoint[0][436]) begin
    filter_input_0_0 = buffer_data_3[3511:3488];
    filter_input_0_1 = buffer_data_2[3511:3488];
    filter_input_0_2 = blur3x3_dout[3511:3488];
    current_RowCol_0 = {img_addr, 10'd437};
  end
  else if (detected_keypoint[0][437]) begin
    filter_input_0_0 = buffer_data_3[3519:3496];
    filter_input_0_1 = buffer_data_2[3519:3496];
    filter_input_0_2 = blur3x3_dout[3519:3496];
    current_RowCol_0 = {img_addr, 10'd438};
  end
  else if (detected_keypoint[0][438]) begin
    filter_input_0_0 = buffer_data_3[3527:3504];
    filter_input_0_1 = buffer_data_2[3527:3504];
    filter_input_0_2 = blur3x3_dout[3527:3504];
    current_RowCol_0 = {img_addr, 10'd439};
  end
  else if (detected_keypoint[0][439]) begin
    filter_input_0_0 = buffer_data_3[3535:3512];
    filter_input_0_1 = buffer_data_2[3535:3512];
    filter_input_0_2 = blur3x3_dout[3535:3512];
    current_RowCol_0 = {img_addr, 10'd440};
  end
  else if (detected_keypoint[0][440]) begin
    filter_input_0_0 = buffer_data_3[3543:3520];
    filter_input_0_1 = buffer_data_2[3543:3520];
    filter_input_0_2 = blur3x3_dout[3543:3520];
    current_RowCol_0 = {img_addr, 10'd441};
  end
  else if (detected_keypoint[0][441]) begin
    filter_input_0_0 = buffer_data_3[3551:3528];
    filter_input_0_1 = buffer_data_2[3551:3528];
    filter_input_0_2 = blur3x3_dout[3551:3528];
    current_RowCol_0 = {img_addr, 10'd442};
  end
  else if (detected_keypoint[0][442]) begin
    filter_input_0_0 = buffer_data_3[3559:3536];
    filter_input_0_1 = buffer_data_2[3559:3536];
    filter_input_0_2 = blur3x3_dout[3559:3536];
    current_RowCol_0 = {img_addr, 10'd443};
  end
  else if (detected_keypoint[0][443]) begin
    filter_input_0_0 = buffer_data_3[3567:3544];
    filter_input_0_1 = buffer_data_2[3567:3544];
    filter_input_0_2 = blur3x3_dout[3567:3544];
    current_RowCol_0 = {img_addr, 10'd444};
  end
  else if (detected_keypoint[0][444]) begin
    filter_input_0_0 = buffer_data_3[3575:3552];
    filter_input_0_1 = buffer_data_2[3575:3552];
    filter_input_0_2 = blur3x3_dout[3575:3552];
    current_RowCol_0 = {img_addr, 10'd445};
  end
  else if (detected_keypoint[0][445]) begin
    filter_input_0_0 = buffer_data_3[3583:3560];
    filter_input_0_1 = buffer_data_2[3583:3560];
    filter_input_0_2 = blur3x3_dout[3583:3560];
    current_RowCol_0 = {img_addr, 10'd446};
  end
  else if (detected_keypoint[0][446]) begin
    filter_input_0_0 = buffer_data_3[3591:3568];
    filter_input_0_1 = buffer_data_2[3591:3568];
    filter_input_0_2 = blur3x3_dout[3591:3568];
    current_RowCol_0 = {img_addr, 10'd447};
  end
  else if (detected_keypoint[0][447]) begin
    filter_input_0_0 = buffer_data_3[3599:3576];
    filter_input_0_1 = buffer_data_2[3599:3576];
    filter_input_0_2 = blur3x3_dout[3599:3576];
    current_RowCol_0 = {img_addr, 10'd448};
  end
  else if (detected_keypoint[0][448]) begin
    filter_input_0_0 = buffer_data_3[3607:3584];
    filter_input_0_1 = buffer_data_2[3607:3584];
    filter_input_0_2 = blur3x3_dout[3607:3584];
    current_RowCol_0 = {img_addr, 10'd449};
  end
  else if (detected_keypoint[0][449]) begin
    filter_input_0_0 = buffer_data_3[3615:3592];
    filter_input_0_1 = buffer_data_2[3615:3592];
    filter_input_0_2 = blur3x3_dout[3615:3592];
    current_RowCol_0 = {img_addr, 10'd450};
  end
  else if (detected_keypoint[0][450]) begin
    filter_input_0_0 = buffer_data_3[3623:3600];
    filter_input_0_1 = buffer_data_2[3623:3600];
    filter_input_0_2 = blur3x3_dout[3623:3600];
    current_RowCol_0 = {img_addr, 10'd451};
  end
  else if (detected_keypoint[0][451]) begin
    filter_input_0_0 = buffer_data_3[3631:3608];
    filter_input_0_1 = buffer_data_2[3631:3608];
    filter_input_0_2 = blur3x3_dout[3631:3608];
    current_RowCol_0 = {img_addr, 10'd452};
  end
  else if (detected_keypoint[0][452]) begin
    filter_input_0_0 = buffer_data_3[3639:3616];
    filter_input_0_1 = buffer_data_2[3639:3616];
    filter_input_0_2 = blur3x3_dout[3639:3616];
    current_RowCol_0 = {img_addr, 10'd453};
  end
  else if (detected_keypoint[0][453]) begin
    filter_input_0_0 = buffer_data_3[3647:3624];
    filter_input_0_1 = buffer_data_2[3647:3624];
    filter_input_0_2 = blur3x3_dout[3647:3624];
    current_RowCol_0 = {img_addr, 10'd454};
  end
  else if (detected_keypoint[0][454]) begin
    filter_input_0_0 = buffer_data_3[3655:3632];
    filter_input_0_1 = buffer_data_2[3655:3632];
    filter_input_0_2 = blur3x3_dout[3655:3632];
    current_RowCol_0 = {img_addr, 10'd455};
  end
  else if (detected_keypoint[0][455]) begin
    filter_input_0_0 = buffer_data_3[3663:3640];
    filter_input_0_1 = buffer_data_2[3663:3640];
    filter_input_0_2 = blur3x3_dout[3663:3640];
    current_RowCol_0 = {img_addr, 10'd456};
  end
  else if (detected_keypoint[0][456]) begin
    filter_input_0_0 = buffer_data_3[3671:3648];
    filter_input_0_1 = buffer_data_2[3671:3648];
    filter_input_0_2 = blur3x3_dout[3671:3648];
    current_RowCol_0 = {img_addr, 10'd457};
  end
  else if (detected_keypoint[0][457]) begin
    filter_input_0_0 = buffer_data_3[3679:3656];
    filter_input_0_1 = buffer_data_2[3679:3656];
    filter_input_0_2 = blur3x3_dout[3679:3656];
    current_RowCol_0 = {img_addr, 10'd458};
  end
  else if (detected_keypoint[0][458]) begin
    filter_input_0_0 = buffer_data_3[3687:3664];
    filter_input_0_1 = buffer_data_2[3687:3664];
    filter_input_0_2 = blur3x3_dout[3687:3664];
    current_RowCol_0 = {img_addr, 10'd459};
  end
  else if (detected_keypoint[0][459]) begin
    filter_input_0_0 = buffer_data_3[3695:3672];
    filter_input_0_1 = buffer_data_2[3695:3672];
    filter_input_0_2 = blur3x3_dout[3695:3672];
    current_RowCol_0 = {img_addr, 10'd460};
  end
  else if (detected_keypoint[0][460]) begin
    filter_input_0_0 = buffer_data_3[3703:3680];
    filter_input_0_1 = buffer_data_2[3703:3680];
    filter_input_0_2 = blur3x3_dout[3703:3680];
    current_RowCol_0 = {img_addr, 10'd461};
  end
  else if (detected_keypoint[0][461]) begin
    filter_input_0_0 = buffer_data_3[3711:3688];
    filter_input_0_1 = buffer_data_2[3711:3688];
    filter_input_0_2 = blur3x3_dout[3711:3688];
    current_RowCol_0 = {img_addr, 10'd462};
  end
  else if (detected_keypoint[0][462]) begin
    filter_input_0_0 = buffer_data_3[3719:3696];
    filter_input_0_1 = buffer_data_2[3719:3696];
    filter_input_0_2 = blur3x3_dout[3719:3696];
    current_RowCol_0 = {img_addr, 10'd463};
  end
  else if (detected_keypoint[0][463]) begin
    filter_input_0_0 = buffer_data_3[3727:3704];
    filter_input_0_1 = buffer_data_2[3727:3704];
    filter_input_0_2 = blur3x3_dout[3727:3704];
    current_RowCol_0 = {img_addr, 10'd464};
  end
  else if (detected_keypoint[0][464]) begin
    filter_input_0_0 = buffer_data_3[3735:3712];
    filter_input_0_1 = buffer_data_2[3735:3712];
    filter_input_0_2 = blur3x3_dout[3735:3712];
    current_RowCol_0 = {img_addr, 10'd465};
  end
  else if (detected_keypoint[0][465]) begin
    filter_input_0_0 = buffer_data_3[3743:3720];
    filter_input_0_1 = buffer_data_2[3743:3720];
    filter_input_0_2 = blur3x3_dout[3743:3720];
    current_RowCol_0 = {img_addr, 10'd466};
  end
  else if (detected_keypoint[0][466]) begin
    filter_input_0_0 = buffer_data_3[3751:3728];
    filter_input_0_1 = buffer_data_2[3751:3728];
    filter_input_0_2 = blur3x3_dout[3751:3728];
    current_RowCol_0 = {img_addr, 10'd467};
  end
  else if (detected_keypoint[0][467]) begin
    filter_input_0_0 = buffer_data_3[3759:3736];
    filter_input_0_1 = buffer_data_2[3759:3736];
    filter_input_0_2 = blur3x3_dout[3759:3736];
    current_RowCol_0 = {img_addr, 10'd468};
  end
  else if (detected_keypoint[0][468]) begin
    filter_input_0_0 = buffer_data_3[3767:3744];
    filter_input_0_1 = buffer_data_2[3767:3744];
    filter_input_0_2 = blur3x3_dout[3767:3744];
    current_RowCol_0 = {img_addr, 10'd469};
  end
  else if (detected_keypoint[0][469]) begin
    filter_input_0_0 = buffer_data_3[3775:3752];
    filter_input_0_1 = buffer_data_2[3775:3752];
    filter_input_0_2 = blur3x3_dout[3775:3752];
    current_RowCol_0 = {img_addr, 10'd470};
  end
  else if (detected_keypoint[0][470]) begin
    filter_input_0_0 = buffer_data_3[3783:3760];
    filter_input_0_1 = buffer_data_2[3783:3760];
    filter_input_0_2 = blur3x3_dout[3783:3760];
    current_RowCol_0 = {img_addr, 10'd471};
  end
  else if (detected_keypoint[0][471]) begin
    filter_input_0_0 = buffer_data_3[3791:3768];
    filter_input_0_1 = buffer_data_2[3791:3768];
    filter_input_0_2 = blur3x3_dout[3791:3768];
    current_RowCol_0 = {img_addr, 10'd472};
  end
  else if (detected_keypoint[0][472]) begin
    filter_input_0_0 = buffer_data_3[3799:3776];
    filter_input_0_1 = buffer_data_2[3799:3776];
    filter_input_0_2 = blur3x3_dout[3799:3776];
    current_RowCol_0 = {img_addr, 10'd473};
  end
  else if (detected_keypoint[0][473]) begin
    filter_input_0_0 = buffer_data_3[3807:3784];
    filter_input_0_1 = buffer_data_2[3807:3784];
    filter_input_0_2 = blur3x3_dout[3807:3784];
    current_RowCol_0 = {img_addr, 10'd474};
  end
  else if (detected_keypoint[0][474]) begin
    filter_input_0_0 = buffer_data_3[3815:3792];
    filter_input_0_1 = buffer_data_2[3815:3792];
    filter_input_0_2 = blur3x3_dout[3815:3792];
    current_RowCol_0 = {img_addr, 10'd475};
  end
  else if (detected_keypoint[0][475]) begin
    filter_input_0_0 = buffer_data_3[3823:3800];
    filter_input_0_1 = buffer_data_2[3823:3800];
    filter_input_0_2 = blur3x3_dout[3823:3800];
    current_RowCol_0 = {img_addr, 10'd476};
  end
  else if (detected_keypoint[0][476]) begin
    filter_input_0_0 = buffer_data_3[3831:3808];
    filter_input_0_1 = buffer_data_2[3831:3808];
    filter_input_0_2 = blur3x3_dout[3831:3808];
    current_RowCol_0 = {img_addr, 10'd477};
  end
  else if (detected_keypoint[0][477]) begin
    filter_input_0_0 = buffer_data_3[3839:3816];
    filter_input_0_1 = buffer_data_2[3839:3816];
    filter_input_0_2 = blur3x3_dout[3839:3816];
    current_RowCol_0 = {img_addr, 10'd478};
  end
  else if (detected_keypoint[0][478]) begin
    filter_input_0_0 = buffer_data_3[3847:3824];
    filter_input_0_1 = buffer_data_2[3847:3824];
    filter_input_0_2 = blur3x3_dout[3847:3824];
    current_RowCol_0 = {img_addr, 10'd479};
  end
  else if (detected_keypoint[0][479]) begin
    filter_input_0_0 = buffer_data_3[3855:3832];
    filter_input_0_1 = buffer_data_2[3855:3832];
    filter_input_0_2 = blur3x3_dout[3855:3832];
    current_RowCol_0 = {img_addr, 10'd480};
  end
  else if (detected_keypoint[0][480]) begin
    filter_input_0_0 = buffer_data_3[3863:3840];
    filter_input_0_1 = buffer_data_2[3863:3840];
    filter_input_0_2 = blur3x3_dout[3863:3840];
    current_RowCol_0 = {img_addr, 10'd481};
  end
  else if (detected_keypoint[0][481]) begin
    filter_input_0_0 = buffer_data_3[3871:3848];
    filter_input_0_1 = buffer_data_2[3871:3848];
    filter_input_0_2 = blur3x3_dout[3871:3848];
    current_RowCol_0 = {img_addr, 10'd482};
  end
  else if (detected_keypoint[0][482]) begin
    filter_input_0_0 = buffer_data_3[3879:3856];
    filter_input_0_1 = buffer_data_2[3879:3856];
    filter_input_0_2 = blur3x3_dout[3879:3856];
    current_RowCol_0 = {img_addr, 10'd483};
  end
  else if (detected_keypoint[0][483]) begin
    filter_input_0_0 = buffer_data_3[3887:3864];
    filter_input_0_1 = buffer_data_2[3887:3864];
    filter_input_0_2 = blur3x3_dout[3887:3864];
    current_RowCol_0 = {img_addr, 10'd484};
  end
  else if (detected_keypoint[0][484]) begin
    filter_input_0_0 = buffer_data_3[3895:3872];
    filter_input_0_1 = buffer_data_2[3895:3872];
    filter_input_0_2 = blur3x3_dout[3895:3872];
    current_RowCol_0 = {img_addr, 10'd485};
  end
  else if (detected_keypoint[0][485]) begin
    filter_input_0_0 = buffer_data_3[3903:3880];
    filter_input_0_1 = buffer_data_2[3903:3880];
    filter_input_0_2 = blur3x3_dout[3903:3880];
    current_RowCol_0 = {img_addr, 10'd486};
  end
  else if (detected_keypoint[0][486]) begin
    filter_input_0_0 = buffer_data_3[3911:3888];
    filter_input_0_1 = buffer_data_2[3911:3888];
    filter_input_0_2 = blur3x3_dout[3911:3888];
    current_RowCol_0 = {img_addr, 10'd487};
  end
  else if (detected_keypoint[0][487]) begin
    filter_input_0_0 = buffer_data_3[3919:3896];
    filter_input_0_1 = buffer_data_2[3919:3896];
    filter_input_0_2 = blur3x3_dout[3919:3896];
    current_RowCol_0 = {img_addr, 10'd488};
  end
  else if (detected_keypoint[0][488]) begin
    filter_input_0_0 = buffer_data_3[3927:3904];
    filter_input_0_1 = buffer_data_2[3927:3904];
    filter_input_0_2 = blur3x3_dout[3927:3904];
    current_RowCol_0 = {img_addr, 10'd489};
  end
  else if (detected_keypoint[0][489]) begin
    filter_input_0_0 = buffer_data_3[3935:3912];
    filter_input_0_1 = buffer_data_2[3935:3912];
    filter_input_0_2 = blur3x3_dout[3935:3912];
    current_RowCol_0 = {img_addr, 10'd490};
  end
  else if (detected_keypoint[0][490]) begin
    filter_input_0_0 = buffer_data_3[3943:3920];
    filter_input_0_1 = buffer_data_2[3943:3920];
    filter_input_0_2 = blur3x3_dout[3943:3920];
    current_RowCol_0 = {img_addr, 10'd491};
  end
  else if (detected_keypoint[0][491]) begin
    filter_input_0_0 = buffer_data_3[3951:3928];
    filter_input_0_1 = buffer_data_2[3951:3928];
    filter_input_0_2 = blur3x3_dout[3951:3928];
    current_RowCol_0 = {img_addr, 10'd492};
  end
  else if (detected_keypoint[0][492]) begin
    filter_input_0_0 = buffer_data_3[3959:3936];
    filter_input_0_1 = buffer_data_2[3959:3936];
    filter_input_0_2 = blur3x3_dout[3959:3936];
    current_RowCol_0 = {img_addr, 10'd493};
  end
  else if (detected_keypoint[0][493]) begin
    filter_input_0_0 = buffer_data_3[3967:3944];
    filter_input_0_1 = buffer_data_2[3967:3944];
    filter_input_0_2 = blur3x3_dout[3967:3944];
    current_RowCol_0 = {img_addr, 10'd494};
  end
  else if (detected_keypoint[0][494]) begin
    filter_input_0_0 = buffer_data_3[3975:3952];
    filter_input_0_1 = buffer_data_2[3975:3952];
    filter_input_0_2 = blur3x3_dout[3975:3952];
    current_RowCol_0 = {img_addr, 10'd495};
  end
  else if (detected_keypoint[0][495]) begin
    filter_input_0_0 = buffer_data_3[3983:3960];
    filter_input_0_1 = buffer_data_2[3983:3960];
    filter_input_0_2 = blur3x3_dout[3983:3960];
    current_RowCol_0 = {img_addr, 10'd496};
  end
  else if (detected_keypoint[0][496]) begin
    filter_input_0_0 = buffer_data_3[3991:3968];
    filter_input_0_1 = buffer_data_2[3991:3968];
    filter_input_0_2 = blur3x3_dout[3991:3968];
    current_RowCol_0 = {img_addr, 10'd497};
  end
  else if (detected_keypoint[0][497]) begin
    filter_input_0_0 = buffer_data_3[3999:3976];
    filter_input_0_1 = buffer_data_2[3999:3976];
    filter_input_0_2 = blur3x3_dout[3999:3976];
    current_RowCol_0 = {img_addr, 10'd498};
  end
  else if (detected_keypoint[0][498]) begin
    filter_input_0_0 = buffer_data_3[4007:3984];
    filter_input_0_1 = buffer_data_2[4007:3984];
    filter_input_0_2 = blur3x3_dout[4007:3984];
    current_RowCol_0 = {img_addr, 10'd499};
  end
  else if (detected_keypoint[0][499]) begin
    filter_input_0_0 = buffer_data_3[4015:3992];
    filter_input_0_1 = buffer_data_2[4015:3992];
    filter_input_0_2 = blur3x3_dout[4015:3992];
    current_RowCol_0 = {img_addr, 10'd500};
  end
  else if (detected_keypoint[0][500]) begin
    filter_input_0_0 = buffer_data_3[4023:4000];
    filter_input_0_1 = buffer_data_2[4023:4000];
    filter_input_0_2 = blur3x3_dout[4023:4000];
    current_RowCol_0 = {img_addr, 10'd501};
  end
  else if (detected_keypoint[0][501]) begin
    filter_input_0_0 = buffer_data_3[4031:4008];
    filter_input_0_1 = buffer_data_2[4031:4008];
    filter_input_0_2 = blur3x3_dout[4031:4008];
    current_RowCol_0 = {img_addr, 10'd502};
  end
  else if (detected_keypoint[0][502]) begin
    filter_input_0_0 = buffer_data_3[4039:4016];
    filter_input_0_1 = buffer_data_2[4039:4016];
    filter_input_0_2 = blur3x3_dout[4039:4016];
    current_RowCol_0 = {img_addr, 10'd503};
  end
  else if (detected_keypoint[0][503]) begin
    filter_input_0_0 = buffer_data_3[4047:4024];
    filter_input_0_1 = buffer_data_2[4047:4024];
    filter_input_0_2 = blur3x3_dout[4047:4024];
    current_RowCol_0 = {img_addr, 10'd504};
  end
  else if (detected_keypoint[0][504]) begin
    filter_input_0_0 = buffer_data_3[4055:4032];
    filter_input_0_1 = buffer_data_2[4055:4032];
    filter_input_0_2 = blur3x3_dout[4055:4032];
    current_RowCol_0 = {img_addr, 10'd505};
  end
  else if (detected_keypoint[0][505]) begin
    filter_input_0_0 = buffer_data_3[4063:4040];
    filter_input_0_1 = buffer_data_2[4063:4040];
    filter_input_0_2 = blur3x3_dout[4063:4040];
    current_RowCol_0 = {img_addr, 10'd506};
  end
  else if (detected_keypoint[0][506]) begin
    filter_input_0_0 = buffer_data_3[4071:4048];
    filter_input_0_1 = buffer_data_2[4071:4048];
    filter_input_0_2 = blur3x3_dout[4071:4048];
    current_RowCol_0 = {img_addr, 10'd507};
  end
  else if (detected_keypoint[0][507]) begin
    filter_input_0_0 = buffer_data_3[4079:4056];
    filter_input_0_1 = buffer_data_2[4079:4056];
    filter_input_0_2 = blur3x3_dout[4079:4056];
    current_RowCol_0 = {img_addr, 10'd508};
  end
  else if (detected_keypoint[0][508]) begin
    filter_input_0_0 = buffer_data_3[4087:4064];
    filter_input_0_1 = buffer_data_2[4087:4064];
    filter_input_0_2 = blur3x3_dout[4087:4064];
    current_RowCol_0 = {img_addr, 10'd509};
  end
  else if (detected_keypoint[0][509]) begin
    filter_input_0_0 = buffer_data_3[4095:4072];
    filter_input_0_1 = buffer_data_2[4095:4072];
    filter_input_0_2 = blur3x3_dout[4095:4072];
    current_RowCol_0 = {img_addr, 10'd510};
  end
  else if (detected_keypoint[0][510]) begin
    filter_input_0_0 = buffer_data_3[4103:4080];
    filter_input_0_1 = buffer_data_2[4103:4080];
    filter_input_0_2 = blur3x3_dout[4103:4080];
    current_RowCol_0 = {img_addr, 10'd511};
  end
  else if (detected_keypoint[0][511]) begin
    filter_input_0_0 = buffer_data_3[4111:4088];
    filter_input_0_1 = buffer_data_2[4111:4088];
    filter_input_0_2 = blur3x3_dout[4111:4088];
    current_RowCol_0 = {img_addr, 10'd512};
  end
  else if (detected_keypoint[0][512]) begin
    filter_input_0_0 = buffer_data_3[4119:4096];
    filter_input_0_1 = buffer_data_2[4119:4096];
    filter_input_0_2 = blur3x3_dout[4119:4096];
    current_RowCol_0 = {img_addr, 10'd513};
  end
  else if (detected_keypoint[0][513]) begin
    filter_input_0_0 = buffer_data_3[4127:4104];
    filter_input_0_1 = buffer_data_2[4127:4104];
    filter_input_0_2 = blur3x3_dout[4127:4104];
    current_RowCol_0 = {img_addr, 10'd514};
  end
  else if (detected_keypoint[0][514]) begin
    filter_input_0_0 = buffer_data_3[4135:4112];
    filter_input_0_1 = buffer_data_2[4135:4112];
    filter_input_0_2 = blur3x3_dout[4135:4112];
    current_RowCol_0 = {img_addr, 10'd515};
  end
  else if (detected_keypoint[0][515]) begin
    filter_input_0_0 = buffer_data_3[4143:4120];
    filter_input_0_1 = buffer_data_2[4143:4120];
    filter_input_0_2 = blur3x3_dout[4143:4120];
    current_RowCol_0 = {img_addr, 10'd516};
  end
  else if (detected_keypoint[0][516]) begin
    filter_input_0_0 = buffer_data_3[4151:4128];
    filter_input_0_1 = buffer_data_2[4151:4128];
    filter_input_0_2 = blur3x3_dout[4151:4128];
    current_RowCol_0 = {img_addr, 10'd517};
  end
  else if (detected_keypoint[0][517]) begin
    filter_input_0_0 = buffer_data_3[4159:4136];
    filter_input_0_1 = buffer_data_2[4159:4136];
    filter_input_0_2 = blur3x3_dout[4159:4136];
    current_RowCol_0 = {img_addr, 10'd518};
  end
  else if (detected_keypoint[0][518]) begin
    filter_input_0_0 = buffer_data_3[4167:4144];
    filter_input_0_1 = buffer_data_2[4167:4144];
    filter_input_0_2 = blur3x3_dout[4167:4144];
    current_RowCol_0 = {img_addr, 10'd519};
  end
  else if (detected_keypoint[0][519]) begin
    filter_input_0_0 = buffer_data_3[4175:4152];
    filter_input_0_1 = buffer_data_2[4175:4152];
    filter_input_0_2 = blur3x3_dout[4175:4152];
    current_RowCol_0 = {img_addr, 10'd520};
  end
  else if (detected_keypoint[0][520]) begin
    filter_input_0_0 = buffer_data_3[4183:4160];
    filter_input_0_1 = buffer_data_2[4183:4160];
    filter_input_0_2 = blur3x3_dout[4183:4160];
    current_RowCol_0 = {img_addr, 10'd521};
  end
  else if (detected_keypoint[0][521]) begin
    filter_input_0_0 = buffer_data_3[4191:4168];
    filter_input_0_1 = buffer_data_2[4191:4168];
    filter_input_0_2 = blur3x3_dout[4191:4168];
    current_RowCol_0 = {img_addr, 10'd522};
  end
  else if (detected_keypoint[0][522]) begin
    filter_input_0_0 = buffer_data_3[4199:4176];
    filter_input_0_1 = buffer_data_2[4199:4176];
    filter_input_0_2 = blur3x3_dout[4199:4176];
    current_RowCol_0 = {img_addr, 10'd523};
  end
  else if (detected_keypoint[0][523]) begin
    filter_input_0_0 = buffer_data_3[4207:4184];
    filter_input_0_1 = buffer_data_2[4207:4184];
    filter_input_0_2 = blur3x3_dout[4207:4184];
    current_RowCol_0 = {img_addr, 10'd524};
  end
  else if (detected_keypoint[0][524]) begin
    filter_input_0_0 = buffer_data_3[4215:4192];
    filter_input_0_1 = buffer_data_2[4215:4192];
    filter_input_0_2 = blur3x3_dout[4215:4192];
    current_RowCol_0 = {img_addr, 10'd525};
  end
  else if (detected_keypoint[0][525]) begin
    filter_input_0_0 = buffer_data_3[4223:4200];
    filter_input_0_1 = buffer_data_2[4223:4200];
    filter_input_0_2 = blur3x3_dout[4223:4200];
    current_RowCol_0 = {img_addr, 10'd526};
  end
  else if (detected_keypoint[0][526]) begin
    filter_input_0_0 = buffer_data_3[4231:4208];
    filter_input_0_1 = buffer_data_2[4231:4208];
    filter_input_0_2 = blur3x3_dout[4231:4208];
    current_RowCol_0 = {img_addr, 10'd527};
  end
  else if (detected_keypoint[0][527]) begin
    filter_input_0_0 = buffer_data_3[4239:4216];
    filter_input_0_1 = buffer_data_2[4239:4216];
    filter_input_0_2 = blur3x3_dout[4239:4216];
    current_RowCol_0 = {img_addr, 10'd528};
  end
  else if (detected_keypoint[0][528]) begin
    filter_input_0_0 = buffer_data_3[4247:4224];
    filter_input_0_1 = buffer_data_2[4247:4224];
    filter_input_0_2 = blur3x3_dout[4247:4224];
    current_RowCol_0 = {img_addr, 10'd529};
  end
  else if (detected_keypoint[0][529]) begin
    filter_input_0_0 = buffer_data_3[4255:4232];
    filter_input_0_1 = buffer_data_2[4255:4232];
    filter_input_0_2 = blur3x3_dout[4255:4232];
    current_RowCol_0 = {img_addr, 10'd530};
  end
  else if (detected_keypoint[0][530]) begin
    filter_input_0_0 = buffer_data_3[4263:4240];
    filter_input_0_1 = buffer_data_2[4263:4240];
    filter_input_0_2 = blur3x3_dout[4263:4240];
    current_RowCol_0 = {img_addr, 10'd531};
  end
  else if (detected_keypoint[0][531]) begin
    filter_input_0_0 = buffer_data_3[4271:4248];
    filter_input_0_1 = buffer_data_2[4271:4248];
    filter_input_0_2 = blur3x3_dout[4271:4248];
    current_RowCol_0 = {img_addr, 10'd532};
  end
  else if (detected_keypoint[0][532]) begin
    filter_input_0_0 = buffer_data_3[4279:4256];
    filter_input_0_1 = buffer_data_2[4279:4256];
    filter_input_0_2 = blur3x3_dout[4279:4256];
    current_RowCol_0 = {img_addr, 10'd533};
  end
  else if (detected_keypoint[0][533]) begin
    filter_input_0_0 = buffer_data_3[4287:4264];
    filter_input_0_1 = buffer_data_2[4287:4264];
    filter_input_0_2 = blur3x3_dout[4287:4264];
    current_RowCol_0 = {img_addr, 10'd534};
  end
  else if (detected_keypoint[0][534]) begin
    filter_input_0_0 = buffer_data_3[4295:4272];
    filter_input_0_1 = buffer_data_2[4295:4272];
    filter_input_0_2 = blur3x3_dout[4295:4272];
    current_RowCol_0 = {img_addr, 10'd535};
  end
  else if (detected_keypoint[0][535]) begin
    filter_input_0_0 = buffer_data_3[4303:4280];
    filter_input_0_1 = buffer_data_2[4303:4280];
    filter_input_0_2 = blur3x3_dout[4303:4280];
    current_RowCol_0 = {img_addr, 10'd536};
  end
  else if (detected_keypoint[0][536]) begin
    filter_input_0_0 = buffer_data_3[4311:4288];
    filter_input_0_1 = buffer_data_2[4311:4288];
    filter_input_0_2 = blur3x3_dout[4311:4288];
    current_RowCol_0 = {img_addr, 10'd537};
  end
  else if (detected_keypoint[0][537]) begin
    filter_input_0_0 = buffer_data_3[4319:4296];
    filter_input_0_1 = buffer_data_2[4319:4296];
    filter_input_0_2 = blur3x3_dout[4319:4296];
    current_RowCol_0 = {img_addr, 10'd538};
  end
  else if (detected_keypoint[0][538]) begin
    filter_input_0_0 = buffer_data_3[4327:4304];
    filter_input_0_1 = buffer_data_2[4327:4304];
    filter_input_0_2 = blur3x3_dout[4327:4304];
    current_RowCol_0 = {img_addr, 10'd539};
  end
  else if (detected_keypoint[0][539]) begin
    filter_input_0_0 = buffer_data_3[4335:4312];
    filter_input_0_1 = buffer_data_2[4335:4312];
    filter_input_0_2 = blur3x3_dout[4335:4312];
    current_RowCol_0 = {img_addr, 10'd540};
  end
  else if (detected_keypoint[0][540]) begin
    filter_input_0_0 = buffer_data_3[4343:4320];
    filter_input_0_1 = buffer_data_2[4343:4320];
    filter_input_0_2 = blur3x3_dout[4343:4320];
    current_RowCol_0 = {img_addr, 10'd541};
  end
  else if (detected_keypoint[0][541]) begin
    filter_input_0_0 = buffer_data_3[4351:4328];
    filter_input_0_1 = buffer_data_2[4351:4328];
    filter_input_0_2 = blur3x3_dout[4351:4328];
    current_RowCol_0 = {img_addr, 10'd542};
  end
  else if (detected_keypoint[0][542]) begin
    filter_input_0_0 = buffer_data_3[4359:4336];
    filter_input_0_1 = buffer_data_2[4359:4336];
    filter_input_0_2 = blur3x3_dout[4359:4336];
    current_RowCol_0 = {img_addr, 10'd543};
  end
  else if (detected_keypoint[0][543]) begin
    filter_input_0_0 = buffer_data_3[4367:4344];
    filter_input_0_1 = buffer_data_2[4367:4344];
    filter_input_0_2 = blur3x3_dout[4367:4344];
    current_RowCol_0 = {img_addr, 10'd544};
  end
  else if (detected_keypoint[0][544]) begin
    filter_input_0_0 = buffer_data_3[4375:4352];
    filter_input_0_1 = buffer_data_2[4375:4352];
    filter_input_0_2 = blur3x3_dout[4375:4352];
    current_RowCol_0 = {img_addr, 10'd545};
  end
  else if (detected_keypoint[0][545]) begin
    filter_input_0_0 = buffer_data_3[4383:4360];
    filter_input_0_1 = buffer_data_2[4383:4360];
    filter_input_0_2 = blur3x3_dout[4383:4360];
    current_RowCol_0 = {img_addr, 10'd546};
  end
  else if (detected_keypoint[0][546]) begin
    filter_input_0_0 = buffer_data_3[4391:4368];
    filter_input_0_1 = buffer_data_2[4391:4368];
    filter_input_0_2 = blur3x3_dout[4391:4368];
    current_RowCol_0 = {img_addr, 10'd547};
  end
  else if (detected_keypoint[0][547]) begin
    filter_input_0_0 = buffer_data_3[4399:4376];
    filter_input_0_1 = buffer_data_2[4399:4376];
    filter_input_0_2 = blur3x3_dout[4399:4376];
    current_RowCol_0 = {img_addr, 10'd548};
  end
  else if (detected_keypoint[0][548]) begin
    filter_input_0_0 = buffer_data_3[4407:4384];
    filter_input_0_1 = buffer_data_2[4407:4384];
    filter_input_0_2 = blur3x3_dout[4407:4384];
    current_RowCol_0 = {img_addr, 10'd549};
  end
  else if (detected_keypoint[0][549]) begin
    filter_input_0_0 = buffer_data_3[4415:4392];
    filter_input_0_1 = buffer_data_2[4415:4392];
    filter_input_0_2 = blur3x3_dout[4415:4392];
    current_RowCol_0 = {img_addr, 10'd550};
  end
  else if (detected_keypoint[0][550]) begin
    filter_input_0_0 = buffer_data_3[4423:4400];
    filter_input_0_1 = buffer_data_2[4423:4400];
    filter_input_0_2 = blur3x3_dout[4423:4400];
    current_RowCol_0 = {img_addr, 10'd551};
  end
  else if (detected_keypoint[0][551]) begin
    filter_input_0_0 = buffer_data_3[4431:4408];
    filter_input_0_1 = buffer_data_2[4431:4408];
    filter_input_0_2 = blur3x3_dout[4431:4408];
    current_RowCol_0 = {img_addr, 10'd552};
  end
  else if (detected_keypoint[0][552]) begin
    filter_input_0_0 = buffer_data_3[4439:4416];
    filter_input_0_1 = buffer_data_2[4439:4416];
    filter_input_0_2 = blur3x3_dout[4439:4416];
    current_RowCol_0 = {img_addr, 10'd553};
  end
  else if (detected_keypoint[0][553]) begin
    filter_input_0_0 = buffer_data_3[4447:4424];
    filter_input_0_1 = buffer_data_2[4447:4424];
    filter_input_0_2 = blur3x3_dout[4447:4424];
    current_RowCol_0 = {img_addr, 10'd554};
  end
  else if (detected_keypoint[0][554]) begin
    filter_input_0_0 = buffer_data_3[4455:4432];
    filter_input_0_1 = buffer_data_2[4455:4432];
    filter_input_0_2 = blur3x3_dout[4455:4432];
    current_RowCol_0 = {img_addr, 10'd555};
  end
  else if (detected_keypoint[0][555]) begin
    filter_input_0_0 = buffer_data_3[4463:4440];
    filter_input_0_1 = buffer_data_2[4463:4440];
    filter_input_0_2 = blur3x3_dout[4463:4440];
    current_RowCol_0 = {img_addr, 10'd556};
  end
  else if (detected_keypoint[0][556]) begin
    filter_input_0_0 = buffer_data_3[4471:4448];
    filter_input_0_1 = buffer_data_2[4471:4448];
    filter_input_0_2 = blur3x3_dout[4471:4448];
    current_RowCol_0 = {img_addr, 10'd557};
  end
  else if (detected_keypoint[0][557]) begin
    filter_input_0_0 = buffer_data_3[4479:4456];
    filter_input_0_1 = buffer_data_2[4479:4456];
    filter_input_0_2 = blur3x3_dout[4479:4456];
    current_RowCol_0 = {img_addr, 10'd558};
  end
  else if (detected_keypoint[0][558]) begin
    filter_input_0_0 = buffer_data_3[4487:4464];
    filter_input_0_1 = buffer_data_2[4487:4464];
    filter_input_0_2 = blur3x3_dout[4487:4464];
    current_RowCol_0 = {img_addr, 10'd559};
  end
  else if (detected_keypoint[0][559]) begin
    filter_input_0_0 = buffer_data_3[4495:4472];
    filter_input_0_1 = buffer_data_2[4495:4472];
    filter_input_0_2 = blur3x3_dout[4495:4472];
    current_RowCol_0 = {img_addr, 10'd560};
  end
  else if (detected_keypoint[0][560]) begin
    filter_input_0_0 = buffer_data_3[4503:4480];
    filter_input_0_1 = buffer_data_2[4503:4480];
    filter_input_0_2 = blur3x3_dout[4503:4480];
    current_RowCol_0 = {img_addr, 10'd561};
  end
  else if (detected_keypoint[0][561]) begin
    filter_input_0_0 = buffer_data_3[4511:4488];
    filter_input_0_1 = buffer_data_2[4511:4488];
    filter_input_0_2 = blur3x3_dout[4511:4488];
    current_RowCol_0 = {img_addr, 10'd562};
  end
  else if (detected_keypoint[0][562]) begin
    filter_input_0_0 = buffer_data_3[4519:4496];
    filter_input_0_1 = buffer_data_2[4519:4496];
    filter_input_0_2 = blur3x3_dout[4519:4496];
    current_RowCol_0 = {img_addr, 10'd563};
  end
  else if (detected_keypoint[0][563]) begin
    filter_input_0_0 = buffer_data_3[4527:4504];
    filter_input_0_1 = buffer_data_2[4527:4504];
    filter_input_0_2 = blur3x3_dout[4527:4504];
    current_RowCol_0 = {img_addr, 10'd564};
  end
  else if (detected_keypoint[0][564]) begin
    filter_input_0_0 = buffer_data_3[4535:4512];
    filter_input_0_1 = buffer_data_2[4535:4512];
    filter_input_0_2 = blur3x3_dout[4535:4512];
    current_RowCol_0 = {img_addr, 10'd565};
  end
  else if (detected_keypoint[0][565]) begin
    filter_input_0_0 = buffer_data_3[4543:4520];
    filter_input_0_1 = buffer_data_2[4543:4520];
    filter_input_0_2 = blur3x3_dout[4543:4520];
    current_RowCol_0 = {img_addr, 10'd566};
  end
  else if (detected_keypoint[0][566]) begin
    filter_input_0_0 = buffer_data_3[4551:4528];
    filter_input_0_1 = buffer_data_2[4551:4528];
    filter_input_0_2 = blur3x3_dout[4551:4528];
    current_RowCol_0 = {img_addr, 10'd567};
  end
  else if (detected_keypoint[0][567]) begin
    filter_input_0_0 = buffer_data_3[4559:4536];
    filter_input_0_1 = buffer_data_2[4559:4536];
    filter_input_0_2 = blur3x3_dout[4559:4536];
    current_RowCol_0 = {img_addr, 10'd568};
  end
  else if (detected_keypoint[0][568]) begin
    filter_input_0_0 = buffer_data_3[4567:4544];
    filter_input_0_1 = buffer_data_2[4567:4544];
    filter_input_0_2 = blur3x3_dout[4567:4544];
    current_RowCol_0 = {img_addr, 10'd569};
  end
  else if (detected_keypoint[0][569]) begin
    filter_input_0_0 = buffer_data_3[4575:4552];
    filter_input_0_1 = buffer_data_2[4575:4552];
    filter_input_0_2 = blur3x3_dout[4575:4552];
    current_RowCol_0 = {img_addr, 10'd570};
  end
  else if (detected_keypoint[0][570]) begin
    filter_input_0_0 = buffer_data_3[4583:4560];
    filter_input_0_1 = buffer_data_2[4583:4560];
    filter_input_0_2 = blur3x3_dout[4583:4560];
    current_RowCol_0 = {img_addr, 10'd571};
  end
  else if (detected_keypoint[0][571]) begin
    filter_input_0_0 = buffer_data_3[4591:4568];
    filter_input_0_1 = buffer_data_2[4591:4568];
    filter_input_0_2 = blur3x3_dout[4591:4568];
    current_RowCol_0 = {img_addr, 10'd572};
  end
  else if (detected_keypoint[0][572]) begin
    filter_input_0_0 = buffer_data_3[4599:4576];
    filter_input_0_1 = buffer_data_2[4599:4576];
    filter_input_0_2 = blur3x3_dout[4599:4576];
    current_RowCol_0 = {img_addr, 10'd573};
  end
  else if (detected_keypoint[0][573]) begin
    filter_input_0_0 = buffer_data_3[4607:4584];
    filter_input_0_1 = buffer_data_2[4607:4584];
    filter_input_0_2 = blur3x3_dout[4607:4584];
    current_RowCol_0 = {img_addr, 10'd574};
  end
  else if (detected_keypoint[0][574]) begin
    filter_input_0_0 = buffer_data_3[4615:4592];
    filter_input_0_1 = buffer_data_2[4615:4592];
    filter_input_0_2 = blur3x3_dout[4615:4592];
    current_RowCol_0 = {img_addr, 10'd575};
  end
  else if (detected_keypoint[0][575]) begin
    filter_input_0_0 = buffer_data_3[4623:4600];
    filter_input_0_1 = buffer_data_2[4623:4600];
    filter_input_0_2 = blur3x3_dout[4623:4600];
    current_RowCol_0 = {img_addr, 10'd576};
  end
  else if (detected_keypoint[0][576]) begin
    filter_input_0_0 = buffer_data_3[4631:4608];
    filter_input_0_1 = buffer_data_2[4631:4608];
    filter_input_0_2 = blur3x3_dout[4631:4608];
    current_RowCol_0 = {img_addr, 10'd577};
  end
  else if (detected_keypoint[0][577]) begin
    filter_input_0_0 = buffer_data_3[4639:4616];
    filter_input_0_1 = buffer_data_2[4639:4616];
    filter_input_0_2 = blur3x3_dout[4639:4616];
    current_RowCol_0 = {img_addr, 10'd578};
  end
  else if (detected_keypoint[0][578]) begin
    filter_input_0_0 = buffer_data_3[4647:4624];
    filter_input_0_1 = buffer_data_2[4647:4624];
    filter_input_0_2 = blur3x3_dout[4647:4624];
    current_RowCol_0 = {img_addr, 10'd579};
  end
  else if (detected_keypoint[0][579]) begin
    filter_input_0_0 = buffer_data_3[4655:4632];
    filter_input_0_1 = buffer_data_2[4655:4632];
    filter_input_0_2 = blur3x3_dout[4655:4632];
    current_RowCol_0 = {img_addr, 10'd580};
  end
  else if (detected_keypoint[0][580]) begin
    filter_input_0_0 = buffer_data_3[4663:4640];
    filter_input_0_1 = buffer_data_2[4663:4640];
    filter_input_0_2 = blur3x3_dout[4663:4640];
    current_RowCol_0 = {img_addr, 10'd581};
  end
  else if (detected_keypoint[0][581]) begin
    filter_input_0_0 = buffer_data_3[4671:4648];
    filter_input_0_1 = buffer_data_2[4671:4648];
    filter_input_0_2 = blur3x3_dout[4671:4648];
    current_RowCol_0 = {img_addr, 10'd582};
  end
  else if (detected_keypoint[0][582]) begin
    filter_input_0_0 = buffer_data_3[4679:4656];
    filter_input_0_1 = buffer_data_2[4679:4656];
    filter_input_0_2 = blur3x3_dout[4679:4656];
    current_RowCol_0 = {img_addr, 10'd583};
  end
  else if (detected_keypoint[0][583]) begin
    filter_input_0_0 = buffer_data_3[4687:4664];
    filter_input_0_1 = buffer_data_2[4687:4664];
    filter_input_0_2 = blur3x3_dout[4687:4664];
    current_RowCol_0 = {img_addr, 10'd584};
  end
  else if (detected_keypoint[0][584]) begin
    filter_input_0_0 = buffer_data_3[4695:4672];
    filter_input_0_1 = buffer_data_2[4695:4672];
    filter_input_0_2 = blur3x3_dout[4695:4672];
    current_RowCol_0 = {img_addr, 10'd585};
  end
  else if (detected_keypoint[0][585]) begin
    filter_input_0_0 = buffer_data_3[4703:4680];
    filter_input_0_1 = buffer_data_2[4703:4680];
    filter_input_0_2 = blur3x3_dout[4703:4680];
    current_RowCol_0 = {img_addr, 10'd586};
  end
  else if (detected_keypoint[0][586]) begin
    filter_input_0_0 = buffer_data_3[4711:4688];
    filter_input_0_1 = buffer_data_2[4711:4688];
    filter_input_0_2 = blur3x3_dout[4711:4688];
    current_RowCol_0 = {img_addr, 10'd587};
  end
  else if (detected_keypoint[0][587]) begin
    filter_input_0_0 = buffer_data_3[4719:4696];
    filter_input_0_1 = buffer_data_2[4719:4696];
    filter_input_0_2 = blur3x3_dout[4719:4696];
    current_RowCol_0 = {img_addr, 10'd588};
  end
  else if (detected_keypoint[0][588]) begin
    filter_input_0_0 = buffer_data_3[4727:4704];
    filter_input_0_1 = buffer_data_2[4727:4704];
    filter_input_0_2 = blur3x3_dout[4727:4704];
    current_RowCol_0 = {img_addr, 10'd589};
  end
  else if (detected_keypoint[0][589]) begin
    filter_input_0_0 = buffer_data_3[4735:4712];
    filter_input_0_1 = buffer_data_2[4735:4712];
    filter_input_0_2 = blur3x3_dout[4735:4712];
    current_RowCol_0 = {img_addr, 10'd590};
  end
  else if (detected_keypoint[0][590]) begin
    filter_input_0_0 = buffer_data_3[4743:4720];
    filter_input_0_1 = buffer_data_2[4743:4720];
    filter_input_0_2 = blur3x3_dout[4743:4720];
    current_RowCol_0 = {img_addr, 10'd591};
  end
  else if (detected_keypoint[0][591]) begin
    filter_input_0_0 = buffer_data_3[4751:4728];
    filter_input_0_1 = buffer_data_2[4751:4728];
    filter_input_0_2 = blur3x3_dout[4751:4728];
    current_RowCol_0 = {img_addr, 10'd592};
  end
  else if (detected_keypoint[0][592]) begin
    filter_input_0_0 = buffer_data_3[4759:4736];
    filter_input_0_1 = buffer_data_2[4759:4736];
    filter_input_0_2 = blur3x3_dout[4759:4736];
    current_RowCol_0 = {img_addr, 10'd593};
  end
  else if (detected_keypoint[0][593]) begin
    filter_input_0_0 = buffer_data_3[4767:4744];
    filter_input_0_1 = buffer_data_2[4767:4744];
    filter_input_0_2 = blur3x3_dout[4767:4744];
    current_RowCol_0 = {img_addr, 10'd594};
  end
  else if (detected_keypoint[0][594]) begin
    filter_input_0_0 = buffer_data_3[4775:4752];
    filter_input_0_1 = buffer_data_2[4775:4752];
    filter_input_0_2 = blur3x3_dout[4775:4752];
    current_RowCol_0 = {img_addr, 10'd595};
  end
  else if (detected_keypoint[0][595]) begin
    filter_input_0_0 = buffer_data_3[4783:4760];
    filter_input_0_1 = buffer_data_2[4783:4760];
    filter_input_0_2 = blur3x3_dout[4783:4760];
    current_RowCol_0 = {img_addr, 10'd596};
  end
  else if (detected_keypoint[0][596]) begin
    filter_input_0_0 = buffer_data_3[4791:4768];
    filter_input_0_1 = buffer_data_2[4791:4768];
    filter_input_0_2 = blur3x3_dout[4791:4768];
    current_RowCol_0 = {img_addr, 10'd597};
  end
  else if (detected_keypoint[0][597]) begin
    filter_input_0_0 = buffer_data_3[4799:4776];
    filter_input_0_1 = buffer_data_2[4799:4776];
    filter_input_0_2 = blur3x3_dout[4799:4776];
    current_RowCol_0 = {img_addr, 10'd598};
  end
  else if (detected_keypoint[0][598]) begin
    filter_input_0_0 = buffer_data_3[4807:4784];
    filter_input_0_1 = buffer_data_2[4807:4784];
    filter_input_0_2 = blur3x3_dout[4807:4784];
    current_RowCol_0 = {img_addr, 10'd599};
  end
  else if (detected_keypoint[0][599]) begin
    filter_input_0_0 = buffer_data_3[4815:4792];
    filter_input_0_1 = buffer_data_2[4815:4792];
    filter_input_0_2 = blur3x3_dout[4815:4792];
    current_RowCol_0 = {img_addr, 10'd600};
  end
  else if (detected_keypoint[0][600]) begin
    filter_input_0_0 = buffer_data_3[4823:4800];
    filter_input_0_1 = buffer_data_2[4823:4800];
    filter_input_0_2 = blur3x3_dout[4823:4800];
    current_RowCol_0 = {img_addr, 10'd601};
  end
  else if (detected_keypoint[0][601]) begin
    filter_input_0_0 = buffer_data_3[4831:4808];
    filter_input_0_1 = buffer_data_2[4831:4808];
    filter_input_0_2 = blur3x3_dout[4831:4808];
    current_RowCol_0 = {img_addr, 10'd602};
  end
  else if (detected_keypoint[0][602]) begin
    filter_input_0_0 = buffer_data_3[4839:4816];
    filter_input_0_1 = buffer_data_2[4839:4816];
    filter_input_0_2 = blur3x3_dout[4839:4816];
    current_RowCol_0 = {img_addr, 10'd603};
  end
  else if (detected_keypoint[0][603]) begin
    filter_input_0_0 = buffer_data_3[4847:4824];
    filter_input_0_1 = buffer_data_2[4847:4824];
    filter_input_0_2 = blur3x3_dout[4847:4824];
    current_RowCol_0 = {img_addr, 10'd604};
  end
  else if (detected_keypoint[0][604]) begin
    filter_input_0_0 = buffer_data_3[4855:4832];
    filter_input_0_1 = buffer_data_2[4855:4832];
    filter_input_0_2 = blur3x3_dout[4855:4832];
    current_RowCol_0 = {img_addr, 10'd605};
  end
  else if (detected_keypoint[0][605]) begin
    filter_input_0_0 = buffer_data_3[4863:4840];
    filter_input_0_1 = buffer_data_2[4863:4840];
    filter_input_0_2 = blur3x3_dout[4863:4840];
    current_RowCol_0 = {img_addr, 10'd606};
  end
  else if (detected_keypoint[0][606]) begin
    filter_input_0_0 = buffer_data_3[4871:4848];
    filter_input_0_1 = buffer_data_2[4871:4848];
    filter_input_0_2 = blur3x3_dout[4871:4848];
    current_RowCol_0 = {img_addr, 10'd607};
  end
  else if (detected_keypoint[0][607]) begin
    filter_input_0_0 = buffer_data_3[4879:4856];
    filter_input_0_1 = buffer_data_2[4879:4856];
    filter_input_0_2 = blur3x3_dout[4879:4856];
    current_RowCol_0 = {img_addr, 10'd608};
  end
  else if (detected_keypoint[0][608]) begin
    filter_input_0_0 = buffer_data_3[4887:4864];
    filter_input_0_1 = buffer_data_2[4887:4864];
    filter_input_0_2 = blur3x3_dout[4887:4864];
    current_RowCol_0 = {img_addr, 10'd609};
  end
  else if (detected_keypoint[0][609]) begin
    filter_input_0_0 = buffer_data_3[4895:4872];
    filter_input_0_1 = buffer_data_2[4895:4872];
    filter_input_0_2 = blur3x3_dout[4895:4872];
    current_RowCol_0 = {img_addr, 10'd610};
  end
  else if (detected_keypoint[0][610]) begin
    filter_input_0_0 = buffer_data_3[4903:4880];
    filter_input_0_1 = buffer_data_2[4903:4880];
    filter_input_0_2 = blur3x3_dout[4903:4880];
    current_RowCol_0 = {img_addr, 10'd611};
  end
  else if (detected_keypoint[0][611]) begin
    filter_input_0_0 = buffer_data_3[4911:4888];
    filter_input_0_1 = buffer_data_2[4911:4888];
    filter_input_0_2 = blur3x3_dout[4911:4888];
    current_RowCol_0 = {img_addr, 10'd612};
  end
  else if (detected_keypoint[0][612]) begin
    filter_input_0_0 = buffer_data_3[4919:4896];
    filter_input_0_1 = buffer_data_2[4919:4896];
    filter_input_0_2 = blur3x3_dout[4919:4896];
    current_RowCol_0 = {img_addr, 10'd613};
  end
  else if (detected_keypoint[0][613]) begin
    filter_input_0_0 = buffer_data_3[4927:4904];
    filter_input_0_1 = buffer_data_2[4927:4904];
    filter_input_0_2 = blur3x3_dout[4927:4904];
    current_RowCol_0 = {img_addr, 10'd614};
  end
  else if (detected_keypoint[0][614]) begin
    filter_input_0_0 = buffer_data_3[4935:4912];
    filter_input_0_1 = buffer_data_2[4935:4912];
    filter_input_0_2 = blur3x3_dout[4935:4912];
    current_RowCol_0 = {img_addr, 10'd615};
  end
  else if (detected_keypoint[0][615]) begin
    filter_input_0_0 = buffer_data_3[4943:4920];
    filter_input_0_1 = buffer_data_2[4943:4920];
    filter_input_0_2 = blur3x3_dout[4943:4920];
    current_RowCol_0 = {img_addr, 10'd616};
  end
  else if (detected_keypoint[0][616]) begin
    filter_input_0_0 = buffer_data_3[4951:4928];
    filter_input_0_1 = buffer_data_2[4951:4928];
    filter_input_0_2 = blur3x3_dout[4951:4928];
    current_RowCol_0 = {img_addr, 10'd617};
  end
  else if (detected_keypoint[0][617]) begin
    filter_input_0_0 = buffer_data_3[4959:4936];
    filter_input_0_1 = buffer_data_2[4959:4936];
    filter_input_0_2 = blur3x3_dout[4959:4936];
    current_RowCol_0 = {img_addr, 10'd618};
  end
  else if (detected_keypoint[0][618]) begin
    filter_input_0_0 = buffer_data_3[4967:4944];
    filter_input_0_1 = buffer_data_2[4967:4944];
    filter_input_0_2 = blur3x3_dout[4967:4944];
    current_RowCol_0 = {img_addr, 10'd619};
  end
  else if (detected_keypoint[0][619]) begin
    filter_input_0_0 = buffer_data_3[4975:4952];
    filter_input_0_1 = buffer_data_2[4975:4952];
    filter_input_0_2 = blur3x3_dout[4975:4952];
    current_RowCol_0 = {img_addr, 10'd620};
  end
  else if (detected_keypoint[0][620]) begin
    filter_input_0_0 = buffer_data_3[4983:4960];
    filter_input_0_1 = buffer_data_2[4983:4960];
    filter_input_0_2 = blur3x3_dout[4983:4960];
    current_RowCol_0 = {img_addr, 10'd621};
  end
  else if (detected_keypoint[0][621]) begin
    filter_input_0_0 = buffer_data_3[4991:4968];
    filter_input_0_1 = buffer_data_2[4991:4968];
    filter_input_0_2 = blur3x3_dout[4991:4968];
    current_RowCol_0 = {img_addr, 10'd622};
  end
  else if (detected_keypoint[0][622]) begin
    filter_input_0_0 = buffer_data_3[4999:4976];
    filter_input_0_1 = buffer_data_2[4999:4976];
    filter_input_0_2 = blur3x3_dout[4999:4976];
    current_RowCol_0 = {img_addr, 10'd623};
  end
  else if (detected_keypoint[0][623]) begin
    filter_input_0_0 = buffer_data_3[5007:4984];
    filter_input_0_1 = buffer_data_2[5007:4984];
    filter_input_0_2 = blur3x3_dout[5007:4984];
    current_RowCol_0 = {img_addr, 10'd624};
  end
  else if (detected_keypoint[0][624]) begin
    filter_input_0_0 = buffer_data_3[5015:4992];
    filter_input_0_1 = buffer_data_2[5015:4992];
    filter_input_0_2 = blur3x3_dout[5015:4992];
    current_RowCol_0 = {img_addr, 10'd625};
  end
  else if (detected_keypoint[0][625]) begin
    filter_input_0_0 = buffer_data_3[5023:5000];
    filter_input_0_1 = buffer_data_2[5023:5000];
    filter_input_0_2 = blur3x3_dout[5023:5000];
    current_RowCol_0 = {img_addr, 10'd626};
  end
  else if (detected_keypoint[0][626]) begin
    filter_input_0_0 = buffer_data_3[5031:5008];
    filter_input_0_1 = buffer_data_2[5031:5008];
    filter_input_0_2 = blur3x3_dout[5031:5008];
    current_RowCol_0 = {img_addr, 10'd627};
  end
  else if (detected_keypoint[0][627]) begin
    filter_input_0_0 = buffer_data_3[5039:5016];
    filter_input_0_1 = buffer_data_2[5039:5016];
    filter_input_0_2 = blur3x3_dout[5039:5016];
    current_RowCol_0 = {img_addr, 10'd628};
  end
  else if (detected_keypoint[0][628]) begin
    filter_input_0_0 = buffer_data_3[5047:5024];
    filter_input_0_1 = buffer_data_2[5047:5024];
    filter_input_0_2 = blur3x3_dout[5047:5024];
    current_RowCol_0 = {img_addr, 10'd629};
  end
  else if (detected_keypoint[0][629]) begin
    filter_input_0_0 = buffer_data_3[5055:5032];
    filter_input_0_1 = buffer_data_2[5055:5032];
    filter_input_0_2 = blur3x3_dout[5055:5032];
    current_RowCol_0 = {img_addr, 10'd630};
  end
  else if (detected_keypoint[0][630]) begin
    filter_input_0_0 = buffer_data_3[5063:5040];
    filter_input_0_1 = buffer_data_2[5063:5040];
    filter_input_0_2 = blur3x3_dout[5063:5040];
    current_RowCol_0 = {img_addr, 10'd631};
  end
  else if (detected_keypoint[0][631]) begin
    filter_input_0_0 = buffer_data_3[5071:5048];
    filter_input_0_1 = buffer_data_2[5071:5048];
    filter_input_0_2 = blur3x3_dout[5071:5048];
    current_RowCol_0 = {img_addr, 10'd632};
  end
  else if (detected_keypoint[0][632]) begin
    filter_input_0_0 = buffer_data_3[5079:5056];
    filter_input_0_1 = buffer_data_2[5079:5056];
    filter_input_0_2 = blur3x3_dout[5079:5056];
    current_RowCol_0 = {img_addr, 10'd633};
  end
  else if (detected_keypoint[0][633]) begin
    filter_input_0_0 = buffer_data_3[5087:5064];
    filter_input_0_1 = buffer_data_2[5087:5064];
    filter_input_0_2 = blur3x3_dout[5087:5064];
    current_RowCol_0 = {img_addr, 10'd634};
  end
  else if (detected_keypoint[0][634]) begin
    filter_input_0_0 = buffer_data_3[5095:5072];
    filter_input_0_1 = buffer_data_2[5095:5072];
    filter_input_0_2 = blur3x3_dout[5095:5072];
    current_RowCol_0 = {img_addr, 10'd635};
  end
  else if (detected_keypoint[0][635]) begin
    filter_input_0_0 = buffer_data_3[5103:5080];
    filter_input_0_1 = buffer_data_2[5103:5080];
    filter_input_0_2 = blur3x3_dout[5103:5080];
    current_RowCol_0 = {img_addr, 10'd636};
  end
  else if (detected_keypoint[0][636]) begin
    filter_input_0_0 = buffer_data_3[5111:5088];
    filter_input_0_1 = buffer_data_2[5111:5088];
    filter_input_0_2 = blur3x3_dout[5111:5088];
    current_RowCol_0 = {img_addr, 10'd637};
  end
  else if (detected_keypoint[0][637]) begin
    filter_input_0_0 = buffer_data_3[5119:5096];
    filter_input_0_1 = buffer_data_2[5119:5096];
    filter_input_0_2 = blur3x3_dout[5119:5096];
    current_RowCol_0 = {img_addr, 10'd638};
  end
  else begin
    filter_input_0_0 = 'd0;
    filter_input_0_1 = 'd0;
    filter_input_0_2 = 'd0;
    current_RowCol_0 = 'd0;
  end

always @(*) begin
  if (detected_keypoint[1][0]) begin
    filter_input_1_0 = buffer_data_5[23:0];
    filter_input_1_1 = buffer_data_4[23:0];
    filter_input_1_2 = blur5x5_1_dout[23:0];
    current_RowCol_1 = {img_addr, 10'd1};
  end
  else if (detected_keypoint[1][1]) begin
    filter_input_1_0 = buffer_data_5[31:8];
    filter_input_1_1 = buffer_data_4[31:8];
    filter_input_1_2 = blur5x5_1_dout[31:8];
    current_RowCol_1 = {img_addr, 10'd2};
  end
  else if (detected_keypoint[1][2]) begin
    filter_input_1_0 = buffer_data_5[39:16];
    filter_input_1_1 = buffer_data_4[39:16];
    filter_input_1_2 = blur5x5_1_dout[39:16];
    current_RowCol_1 = {img_addr, 10'd3};
  end
  else if (detected_keypoint[1][3]) begin
    filter_input_1_0 = buffer_data_5[47:24];
    filter_input_1_1 = buffer_data_4[47:24];
    filter_input_1_2 = blur5x5_1_dout[47:24];
    current_RowCol_1 = {img_addr, 10'd4};
  end
  else if (detected_keypoint[1][4]) begin
    filter_input_1_0 = buffer_data_5[55:32];
    filter_input_1_1 = buffer_data_4[55:32];
    filter_input_1_2 = blur5x5_1_dout[55:32];
    current_RowCol_1 = {img_addr, 10'd5};
  end
  else if (detected_keypoint[1][5]) begin
    filter_input_1_0 = buffer_data_5[63:40];
    filter_input_1_1 = buffer_data_4[63:40];
    filter_input_1_2 = blur5x5_1_dout[63:40];
    current_RowCol_1 = {img_addr, 10'd6};
  end
  else if (detected_keypoint[1][6]) begin
    filter_input_1_0 = buffer_data_5[71:48];
    filter_input_1_1 = buffer_data_4[71:48];
    filter_input_1_2 = blur5x5_1_dout[71:48];
    current_RowCol_1 = {img_addr, 10'd7};
  end
  else if (detected_keypoint[1][7]) begin
    filter_input_1_0 = buffer_data_5[79:56];
    filter_input_1_1 = buffer_data_4[79:56];
    filter_input_1_2 = blur5x5_1_dout[79:56];
    current_RowCol_1 = {img_addr, 10'd8};
  end
  else if (detected_keypoint[1][8]) begin
    filter_input_1_0 = buffer_data_5[87:64];
    filter_input_1_1 = buffer_data_4[87:64];
    filter_input_1_2 = blur5x5_1_dout[87:64];
    current_RowCol_1 = {img_addr, 10'd9};
  end
  else if (detected_keypoint[1][9]) begin
    filter_input_1_0 = buffer_data_5[95:72];
    filter_input_1_1 = buffer_data_4[95:72];
    filter_input_1_2 = blur5x5_1_dout[95:72];
    current_RowCol_1 = {img_addr, 10'd10};
  end
  else if (detected_keypoint[1][10]) begin
    filter_input_1_0 = buffer_data_5[103:80];
    filter_input_1_1 = buffer_data_4[103:80];
    filter_input_1_2 = blur5x5_1_dout[103:80];
    current_RowCol_1 = {img_addr, 10'd11};
  end
  else if (detected_keypoint[1][11]) begin
    filter_input_1_0 = buffer_data_5[111:88];
    filter_input_1_1 = buffer_data_4[111:88];
    filter_input_1_2 = blur5x5_1_dout[111:88];
    current_RowCol_1 = {img_addr, 10'd12};
  end
  else if (detected_keypoint[1][12]) begin
    filter_input_1_0 = buffer_data_5[119:96];
    filter_input_1_1 = buffer_data_4[119:96];
    filter_input_1_2 = blur5x5_1_dout[119:96];
    current_RowCol_1 = {img_addr, 10'd13};
  end
  else if (detected_keypoint[1][13]) begin
    filter_input_1_0 = buffer_data_5[127:104];
    filter_input_1_1 = buffer_data_4[127:104];
    filter_input_1_2 = blur5x5_1_dout[127:104];
    current_RowCol_1 = {img_addr, 10'd14};
  end
  else if (detected_keypoint[1][14]) begin
    filter_input_1_0 = buffer_data_5[135:112];
    filter_input_1_1 = buffer_data_4[135:112];
    filter_input_1_2 = blur5x5_1_dout[135:112];
    current_RowCol_1 = {img_addr, 10'd15};
  end
  else if (detected_keypoint[1][15]) begin
    filter_input_1_0 = buffer_data_5[143:120];
    filter_input_1_1 = buffer_data_4[143:120];
    filter_input_1_2 = blur5x5_1_dout[143:120];
    current_RowCol_1 = {img_addr, 10'd16};
  end
  else if (detected_keypoint[1][16]) begin
    filter_input_1_0 = buffer_data_5[151:128];
    filter_input_1_1 = buffer_data_4[151:128];
    filter_input_1_2 = blur5x5_1_dout[151:128];
    current_RowCol_1 = {img_addr, 10'd17};
  end
  else if (detected_keypoint[1][17]) begin
    filter_input_1_0 = buffer_data_5[159:136];
    filter_input_1_1 = buffer_data_4[159:136];
    filter_input_1_2 = blur5x5_1_dout[159:136];
    current_RowCol_1 = {img_addr, 10'd18};
  end
  else if (detected_keypoint[1][18]) begin
    filter_input_1_0 = buffer_data_5[167:144];
    filter_input_1_1 = buffer_data_4[167:144];
    filter_input_1_2 = blur5x5_1_dout[167:144];
    current_RowCol_1 = {img_addr, 10'd19};
  end
  else if (detected_keypoint[1][19]) begin
    filter_input_1_0 = buffer_data_5[175:152];
    filter_input_1_1 = buffer_data_4[175:152];
    filter_input_1_2 = blur5x5_1_dout[175:152];
    current_RowCol_1 = {img_addr, 10'd20};
  end
  else if (detected_keypoint[1][20]) begin
    filter_input_1_0 = buffer_data_5[183:160];
    filter_input_1_1 = buffer_data_4[183:160];
    filter_input_1_2 = blur5x5_1_dout[183:160];
    current_RowCol_1 = {img_addr, 10'd21};
  end
  else if (detected_keypoint[1][21]) begin
    filter_input_1_0 = buffer_data_5[191:168];
    filter_input_1_1 = buffer_data_4[191:168];
    filter_input_1_2 = blur5x5_1_dout[191:168];
    current_RowCol_1 = {img_addr, 10'd22};
  end
  else if (detected_keypoint[1][22]) begin
    filter_input_1_0 = buffer_data_5[199:176];
    filter_input_1_1 = buffer_data_4[199:176];
    filter_input_1_2 = blur5x5_1_dout[199:176];
    current_RowCol_1 = {img_addr, 10'd23};
  end
  else if (detected_keypoint[1][23]) begin
    filter_input_1_0 = buffer_data_5[207:184];
    filter_input_1_1 = buffer_data_4[207:184];
    filter_input_1_2 = blur5x5_1_dout[207:184];
    current_RowCol_1 = {img_addr, 10'd24};
  end
  else if (detected_keypoint[1][24]) begin
    filter_input_1_0 = buffer_data_5[215:192];
    filter_input_1_1 = buffer_data_4[215:192];
    filter_input_1_2 = blur5x5_1_dout[215:192];
    current_RowCol_1 = {img_addr, 10'd25};
  end
  else if (detected_keypoint[1][25]) begin
    filter_input_1_0 = buffer_data_5[223:200];
    filter_input_1_1 = buffer_data_4[223:200];
    filter_input_1_2 = blur5x5_1_dout[223:200];
    current_RowCol_1 = {img_addr, 10'd26};
  end
  else if (detected_keypoint[1][26]) begin
    filter_input_1_0 = buffer_data_5[231:208];
    filter_input_1_1 = buffer_data_4[231:208];
    filter_input_1_2 = blur5x5_1_dout[231:208];
    current_RowCol_1 = {img_addr, 10'd27};
  end
  else if (detected_keypoint[1][27]) begin
    filter_input_1_0 = buffer_data_5[239:216];
    filter_input_1_1 = buffer_data_4[239:216];
    filter_input_1_2 = blur5x5_1_dout[239:216];
    current_RowCol_1 = {img_addr, 10'd28};
  end
  else if (detected_keypoint[1][28]) begin
    filter_input_1_0 = buffer_data_5[247:224];
    filter_input_1_1 = buffer_data_4[247:224];
    filter_input_1_2 = blur5x5_1_dout[247:224];
    current_RowCol_1 = {img_addr, 10'd29};
  end
  else if (detected_keypoint[1][29]) begin
    filter_input_1_0 = buffer_data_5[255:232];
    filter_input_1_1 = buffer_data_4[255:232];
    filter_input_1_2 = blur5x5_1_dout[255:232];
    current_RowCol_1 = {img_addr, 10'd30};
  end
  else if (detected_keypoint[1][30]) begin
    filter_input_1_0 = buffer_data_5[263:240];
    filter_input_1_1 = buffer_data_4[263:240];
    filter_input_1_2 = blur5x5_1_dout[263:240];
    current_RowCol_1 = {img_addr, 10'd31};
  end
  else if (detected_keypoint[1][31]) begin
    filter_input_1_0 = buffer_data_5[271:248];
    filter_input_1_1 = buffer_data_4[271:248];
    filter_input_1_2 = blur5x5_1_dout[271:248];
    current_RowCol_1 = {img_addr, 10'd32};
  end
  else if (detected_keypoint[1][32]) begin
    filter_input_1_0 = buffer_data_5[279:256];
    filter_input_1_1 = buffer_data_4[279:256];
    filter_input_1_2 = blur5x5_1_dout[279:256];
    current_RowCol_1 = {img_addr, 10'd33};
  end
  else if (detected_keypoint[1][33]) begin
    filter_input_1_0 = buffer_data_5[287:264];
    filter_input_1_1 = buffer_data_4[287:264];
    filter_input_1_2 = blur5x5_1_dout[287:264];
    current_RowCol_1 = {img_addr, 10'd34};
  end
  else if (detected_keypoint[1][34]) begin
    filter_input_1_0 = buffer_data_5[295:272];
    filter_input_1_1 = buffer_data_4[295:272];
    filter_input_1_2 = blur5x5_1_dout[295:272];
    current_RowCol_1 = {img_addr, 10'd35};
  end
  else if (detected_keypoint[1][35]) begin
    filter_input_1_0 = buffer_data_5[303:280];
    filter_input_1_1 = buffer_data_4[303:280];
    filter_input_1_2 = blur5x5_1_dout[303:280];
    current_RowCol_1 = {img_addr, 10'd36};
  end
  else if (detected_keypoint[1][36]) begin
    filter_input_1_0 = buffer_data_5[311:288];
    filter_input_1_1 = buffer_data_4[311:288];
    filter_input_1_2 = blur5x5_1_dout[311:288];
    current_RowCol_1 = {img_addr, 10'd37};
  end
  else if (detected_keypoint[1][37]) begin
    filter_input_1_0 = buffer_data_5[319:296];
    filter_input_1_1 = buffer_data_4[319:296];
    filter_input_1_2 = blur5x5_1_dout[319:296];
    current_RowCol_1 = {img_addr, 10'd38};
  end
  else if (detected_keypoint[1][38]) begin
    filter_input_1_0 = buffer_data_5[327:304];
    filter_input_1_1 = buffer_data_4[327:304];
    filter_input_1_2 = blur5x5_1_dout[327:304];
    current_RowCol_1 = {img_addr, 10'd39};
  end
  else if (detected_keypoint[1][39]) begin
    filter_input_1_0 = buffer_data_5[335:312];
    filter_input_1_1 = buffer_data_4[335:312];
    filter_input_1_2 = blur5x5_1_dout[335:312];
    current_RowCol_1 = {img_addr, 10'd40};
  end
  else if (detected_keypoint[1][40]) begin
    filter_input_1_0 = buffer_data_5[343:320];
    filter_input_1_1 = buffer_data_4[343:320];
    filter_input_1_2 = blur5x5_1_dout[343:320];
    current_RowCol_1 = {img_addr, 10'd41};
  end
  else if (detected_keypoint[1][41]) begin
    filter_input_1_0 = buffer_data_5[351:328];
    filter_input_1_1 = buffer_data_4[351:328];
    filter_input_1_2 = blur5x5_1_dout[351:328];
    current_RowCol_1 = {img_addr, 10'd42};
  end
  else if (detected_keypoint[1][42]) begin
    filter_input_1_0 = buffer_data_5[359:336];
    filter_input_1_1 = buffer_data_4[359:336];
    filter_input_1_2 = blur5x5_1_dout[359:336];
    current_RowCol_1 = {img_addr, 10'd43};
  end
  else if (detected_keypoint[1][43]) begin
    filter_input_1_0 = buffer_data_5[367:344];
    filter_input_1_1 = buffer_data_4[367:344];
    filter_input_1_2 = blur5x5_1_dout[367:344];
    current_RowCol_1 = {img_addr, 10'd44};
  end
  else if (detected_keypoint[1][44]) begin
    filter_input_1_0 = buffer_data_5[375:352];
    filter_input_1_1 = buffer_data_4[375:352];
    filter_input_1_2 = blur5x5_1_dout[375:352];
    current_RowCol_1 = {img_addr, 10'd45};
  end
  else if (detected_keypoint[1][45]) begin
    filter_input_1_0 = buffer_data_5[383:360];
    filter_input_1_1 = buffer_data_4[383:360];
    filter_input_1_2 = blur5x5_1_dout[383:360];
    current_RowCol_1 = {img_addr, 10'd46};
  end
  else if (detected_keypoint[1][46]) begin
    filter_input_1_0 = buffer_data_5[391:368];
    filter_input_1_1 = buffer_data_4[391:368];
    filter_input_1_2 = blur5x5_1_dout[391:368];
    current_RowCol_1 = {img_addr, 10'd47};
  end
  else if (detected_keypoint[1][47]) begin
    filter_input_1_0 = buffer_data_5[399:376];
    filter_input_1_1 = buffer_data_4[399:376];
    filter_input_1_2 = blur5x5_1_dout[399:376];
    current_RowCol_1 = {img_addr, 10'd48};
  end
  else if (detected_keypoint[1][48]) begin
    filter_input_1_0 = buffer_data_5[407:384];
    filter_input_1_1 = buffer_data_4[407:384];
    filter_input_1_2 = blur5x5_1_dout[407:384];
    current_RowCol_1 = {img_addr, 10'd49};
  end
  else if (detected_keypoint[1][49]) begin
    filter_input_1_0 = buffer_data_5[415:392];
    filter_input_1_1 = buffer_data_4[415:392];
    filter_input_1_2 = blur5x5_1_dout[415:392];
    current_RowCol_1 = {img_addr, 10'd50};
  end
  else if (detected_keypoint[1][50]) begin
    filter_input_1_0 = buffer_data_5[423:400];
    filter_input_1_1 = buffer_data_4[423:400];
    filter_input_1_2 = blur5x5_1_dout[423:400];
    current_RowCol_1 = {img_addr, 10'd51};
  end
  else if (detected_keypoint[1][51]) begin
    filter_input_1_0 = buffer_data_5[431:408];
    filter_input_1_1 = buffer_data_4[431:408];
    filter_input_1_2 = blur5x5_1_dout[431:408];
    current_RowCol_1 = {img_addr, 10'd52};
  end
  else if (detected_keypoint[1][52]) begin
    filter_input_1_0 = buffer_data_5[439:416];
    filter_input_1_1 = buffer_data_4[439:416];
    filter_input_1_2 = blur5x5_1_dout[439:416];
    current_RowCol_1 = {img_addr, 10'd53};
  end
  else if (detected_keypoint[1][53]) begin
    filter_input_1_0 = buffer_data_5[447:424];
    filter_input_1_1 = buffer_data_4[447:424];
    filter_input_1_2 = blur5x5_1_dout[447:424];
    current_RowCol_1 = {img_addr, 10'd54};
  end
  else if (detected_keypoint[1][54]) begin
    filter_input_1_0 = buffer_data_5[455:432];
    filter_input_1_1 = buffer_data_4[455:432];
    filter_input_1_2 = blur5x5_1_dout[455:432];
    current_RowCol_1 = {img_addr, 10'd55};
  end
  else if (detected_keypoint[1][55]) begin
    filter_input_1_0 = buffer_data_5[463:440];
    filter_input_1_1 = buffer_data_4[463:440];
    filter_input_1_2 = blur5x5_1_dout[463:440];
    current_RowCol_1 = {img_addr, 10'd56};
  end
  else if (detected_keypoint[1][56]) begin
    filter_input_1_0 = buffer_data_5[471:448];
    filter_input_1_1 = buffer_data_4[471:448];
    filter_input_1_2 = blur5x5_1_dout[471:448];
    current_RowCol_1 = {img_addr, 10'd57};
  end
  else if (detected_keypoint[1][57]) begin
    filter_input_1_0 = buffer_data_5[479:456];
    filter_input_1_1 = buffer_data_4[479:456];
    filter_input_1_2 = blur5x5_1_dout[479:456];
    current_RowCol_1 = {img_addr, 10'd58};
  end
  else if (detected_keypoint[1][58]) begin
    filter_input_1_0 = buffer_data_5[487:464];
    filter_input_1_1 = buffer_data_4[487:464];
    filter_input_1_2 = blur5x5_1_dout[487:464];
    current_RowCol_1 = {img_addr, 10'd59};
  end
  else if (detected_keypoint[1][59]) begin
    filter_input_1_0 = buffer_data_5[495:472];
    filter_input_1_1 = buffer_data_4[495:472];
    filter_input_1_2 = blur5x5_1_dout[495:472];
    current_RowCol_1 = {img_addr, 10'd60};
  end
  else if (detected_keypoint[1][60]) begin
    filter_input_1_0 = buffer_data_5[503:480];
    filter_input_1_1 = buffer_data_4[503:480];
    filter_input_1_2 = blur5x5_1_dout[503:480];
    current_RowCol_1 = {img_addr, 10'd61};
  end
  else if (detected_keypoint[1][61]) begin
    filter_input_1_0 = buffer_data_5[511:488];
    filter_input_1_1 = buffer_data_4[511:488];
    filter_input_1_2 = blur5x5_1_dout[511:488];
    current_RowCol_1 = {img_addr, 10'd62};
  end
  else if (detected_keypoint[1][62]) begin
    filter_input_1_0 = buffer_data_5[519:496];
    filter_input_1_1 = buffer_data_4[519:496];
    filter_input_1_2 = blur5x5_1_dout[519:496];
    current_RowCol_1 = {img_addr, 10'd63};
  end
  else if (detected_keypoint[1][63]) begin
    filter_input_1_0 = buffer_data_5[527:504];
    filter_input_1_1 = buffer_data_4[527:504];
    filter_input_1_2 = blur5x5_1_dout[527:504];
    current_RowCol_1 = {img_addr, 10'd64};
  end
  else if (detected_keypoint[1][64]) begin
    filter_input_1_0 = buffer_data_5[535:512];
    filter_input_1_1 = buffer_data_4[535:512];
    filter_input_1_2 = blur5x5_1_dout[535:512];
    current_RowCol_1 = {img_addr, 10'd65};
  end
  else if (detected_keypoint[1][65]) begin
    filter_input_1_0 = buffer_data_5[543:520];
    filter_input_1_1 = buffer_data_4[543:520];
    filter_input_1_2 = blur5x5_1_dout[543:520];
    current_RowCol_1 = {img_addr, 10'd66};
  end
  else if (detected_keypoint[1][66]) begin
    filter_input_1_0 = buffer_data_5[551:528];
    filter_input_1_1 = buffer_data_4[551:528];
    filter_input_1_2 = blur5x5_1_dout[551:528];
    current_RowCol_1 = {img_addr, 10'd67};
  end
  else if (detected_keypoint[1][67]) begin
    filter_input_1_0 = buffer_data_5[559:536];
    filter_input_1_1 = buffer_data_4[559:536];
    filter_input_1_2 = blur5x5_1_dout[559:536];
    current_RowCol_1 = {img_addr, 10'd68};
  end
  else if (detected_keypoint[1][68]) begin
    filter_input_1_0 = buffer_data_5[567:544];
    filter_input_1_1 = buffer_data_4[567:544];
    filter_input_1_2 = blur5x5_1_dout[567:544];
    current_RowCol_1 = {img_addr, 10'd69};
  end
  else if (detected_keypoint[1][69]) begin
    filter_input_1_0 = buffer_data_5[575:552];
    filter_input_1_1 = buffer_data_4[575:552];
    filter_input_1_2 = blur5x5_1_dout[575:552];
    current_RowCol_1 = {img_addr, 10'd70};
  end
  else if (detected_keypoint[1][70]) begin
    filter_input_1_0 = buffer_data_5[583:560];
    filter_input_1_1 = buffer_data_4[583:560];
    filter_input_1_2 = blur5x5_1_dout[583:560];
    current_RowCol_1 = {img_addr, 10'd71};
  end
  else if (detected_keypoint[1][71]) begin
    filter_input_1_0 = buffer_data_5[591:568];
    filter_input_1_1 = buffer_data_4[591:568];
    filter_input_1_2 = blur5x5_1_dout[591:568];
    current_RowCol_1 = {img_addr, 10'd72};
  end
  else if (detected_keypoint[1][72]) begin
    filter_input_1_0 = buffer_data_5[599:576];
    filter_input_1_1 = buffer_data_4[599:576];
    filter_input_1_2 = blur5x5_1_dout[599:576];
    current_RowCol_1 = {img_addr, 10'd73};
  end
  else if (detected_keypoint[1][73]) begin
    filter_input_1_0 = buffer_data_5[607:584];
    filter_input_1_1 = buffer_data_4[607:584];
    filter_input_1_2 = blur5x5_1_dout[607:584];
    current_RowCol_1 = {img_addr, 10'd74};
  end
  else if (detected_keypoint[1][74]) begin
    filter_input_1_0 = buffer_data_5[615:592];
    filter_input_1_1 = buffer_data_4[615:592];
    filter_input_1_2 = blur5x5_1_dout[615:592];
    current_RowCol_1 = {img_addr, 10'd75};
  end
  else if (detected_keypoint[1][75]) begin
    filter_input_1_0 = buffer_data_5[623:600];
    filter_input_1_1 = buffer_data_4[623:600];
    filter_input_1_2 = blur5x5_1_dout[623:600];
    current_RowCol_1 = {img_addr, 10'd76};
  end
  else if (detected_keypoint[1][76]) begin
    filter_input_1_0 = buffer_data_5[631:608];
    filter_input_1_1 = buffer_data_4[631:608];
    filter_input_1_2 = blur5x5_1_dout[631:608];
    current_RowCol_1 = {img_addr, 10'd77};
  end
  else if (detected_keypoint[1][77]) begin
    filter_input_1_0 = buffer_data_5[639:616];
    filter_input_1_1 = buffer_data_4[639:616];
    filter_input_1_2 = blur5x5_1_dout[639:616];
    current_RowCol_1 = {img_addr, 10'd78};
  end
  else if (detected_keypoint[1][78]) begin
    filter_input_1_0 = buffer_data_5[647:624];
    filter_input_1_1 = buffer_data_4[647:624];
    filter_input_1_2 = blur5x5_1_dout[647:624];
    current_RowCol_1 = {img_addr, 10'd79};
  end
  else if (detected_keypoint[1][79]) begin
    filter_input_1_0 = buffer_data_5[655:632];
    filter_input_1_1 = buffer_data_4[655:632];
    filter_input_1_2 = blur5x5_1_dout[655:632];
    current_RowCol_1 = {img_addr, 10'd80};
  end
  else if (detected_keypoint[1][80]) begin
    filter_input_1_0 = buffer_data_5[663:640];
    filter_input_1_1 = buffer_data_4[663:640];
    filter_input_1_2 = blur5x5_1_dout[663:640];
    current_RowCol_1 = {img_addr, 10'd81};
  end
  else if (detected_keypoint[1][81]) begin
    filter_input_1_0 = buffer_data_5[671:648];
    filter_input_1_1 = buffer_data_4[671:648];
    filter_input_1_2 = blur5x5_1_dout[671:648];
    current_RowCol_1 = {img_addr, 10'd82};
  end
  else if (detected_keypoint[1][82]) begin
    filter_input_1_0 = buffer_data_5[679:656];
    filter_input_1_1 = buffer_data_4[679:656];
    filter_input_1_2 = blur5x5_1_dout[679:656];
    current_RowCol_1 = {img_addr, 10'd83};
  end
  else if (detected_keypoint[1][83]) begin
    filter_input_1_0 = buffer_data_5[687:664];
    filter_input_1_1 = buffer_data_4[687:664];
    filter_input_1_2 = blur5x5_1_dout[687:664];
    current_RowCol_1 = {img_addr, 10'd84};
  end
  else if (detected_keypoint[1][84]) begin
    filter_input_1_0 = buffer_data_5[695:672];
    filter_input_1_1 = buffer_data_4[695:672];
    filter_input_1_2 = blur5x5_1_dout[695:672];
    current_RowCol_1 = {img_addr, 10'd85};
  end
  else if (detected_keypoint[1][85]) begin
    filter_input_1_0 = buffer_data_5[703:680];
    filter_input_1_1 = buffer_data_4[703:680];
    filter_input_1_2 = blur5x5_1_dout[703:680];
    current_RowCol_1 = {img_addr, 10'd86};
  end
  else if (detected_keypoint[1][86]) begin
    filter_input_1_0 = buffer_data_5[711:688];
    filter_input_1_1 = buffer_data_4[711:688];
    filter_input_1_2 = blur5x5_1_dout[711:688];
    current_RowCol_1 = {img_addr, 10'd87};
  end
  else if (detected_keypoint[1][87]) begin
    filter_input_1_0 = buffer_data_5[719:696];
    filter_input_1_1 = buffer_data_4[719:696];
    filter_input_1_2 = blur5x5_1_dout[719:696];
    current_RowCol_1 = {img_addr, 10'd88};
  end
  else if (detected_keypoint[1][88]) begin
    filter_input_1_0 = buffer_data_5[727:704];
    filter_input_1_1 = buffer_data_4[727:704];
    filter_input_1_2 = blur5x5_1_dout[727:704];
    current_RowCol_1 = {img_addr, 10'd89};
  end
  else if (detected_keypoint[1][89]) begin
    filter_input_1_0 = buffer_data_5[735:712];
    filter_input_1_1 = buffer_data_4[735:712];
    filter_input_1_2 = blur5x5_1_dout[735:712];
    current_RowCol_1 = {img_addr, 10'd90};
  end
  else if (detected_keypoint[1][90]) begin
    filter_input_1_0 = buffer_data_5[743:720];
    filter_input_1_1 = buffer_data_4[743:720];
    filter_input_1_2 = blur5x5_1_dout[743:720];
    current_RowCol_1 = {img_addr, 10'd91};
  end
  else if (detected_keypoint[1][91]) begin
    filter_input_1_0 = buffer_data_5[751:728];
    filter_input_1_1 = buffer_data_4[751:728];
    filter_input_1_2 = blur5x5_1_dout[751:728];
    current_RowCol_1 = {img_addr, 10'd92};
  end
  else if (detected_keypoint[1][92]) begin
    filter_input_1_0 = buffer_data_5[759:736];
    filter_input_1_1 = buffer_data_4[759:736];
    filter_input_1_2 = blur5x5_1_dout[759:736];
    current_RowCol_1 = {img_addr, 10'd93};
  end
  else if (detected_keypoint[1][93]) begin
    filter_input_1_0 = buffer_data_5[767:744];
    filter_input_1_1 = buffer_data_4[767:744];
    filter_input_1_2 = blur5x5_1_dout[767:744];
    current_RowCol_1 = {img_addr, 10'd94};
  end
  else if (detected_keypoint[1][94]) begin
    filter_input_1_0 = buffer_data_5[775:752];
    filter_input_1_1 = buffer_data_4[775:752];
    filter_input_1_2 = blur5x5_1_dout[775:752];
    current_RowCol_1 = {img_addr, 10'd95};
  end
  else if (detected_keypoint[1][95]) begin
    filter_input_1_0 = buffer_data_5[783:760];
    filter_input_1_1 = buffer_data_4[783:760];
    filter_input_1_2 = blur5x5_1_dout[783:760];
    current_RowCol_1 = {img_addr, 10'd96};
  end
  else if (detected_keypoint[1][96]) begin
    filter_input_1_0 = buffer_data_5[791:768];
    filter_input_1_1 = buffer_data_4[791:768];
    filter_input_1_2 = blur5x5_1_dout[791:768];
    current_RowCol_1 = {img_addr, 10'd97};
  end
  else if (detected_keypoint[1][97]) begin
    filter_input_1_0 = buffer_data_5[799:776];
    filter_input_1_1 = buffer_data_4[799:776];
    filter_input_1_2 = blur5x5_1_dout[799:776];
    current_RowCol_1 = {img_addr, 10'd98};
  end
  else if (detected_keypoint[1][98]) begin
    filter_input_1_0 = buffer_data_5[807:784];
    filter_input_1_1 = buffer_data_4[807:784];
    filter_input_1_2 = blur5x5_1_dout[807:784];
    current_RowCol_1 = {img_addr, 10'd99};
  end
  else if (detected_keypoint[1][99]) begin
    filter_input_1_0 = buffer_data_5[815:792];
    filter_input_1_1 = buffer_data_4[815:792];
    filter_input_1_2 = blur5x5_1_dout[815:792];
    current_RowCol_1 = {img_addr, 10'd100};
  end
  else if (detected_keypoint[1][100]) begin
    filter_input_1_0 = buffer_data_5[823:800];
    filter_input_1_1 = buffer_data_4[823:800];
    filter_input_1_2 = blur5x5_1_dout[823:800];
    current_RowCol_1 = {img_addr, 10'd101};
  end
  else if (detected_keypoint[1][101]) begin
    filter_input_1_0 = buffer_data_5[831:808];
    filter_input_1_1 = buffer_data_4[831:808];
    filter_input_1_2 = blur5x5_1_dout[831:808];
    current_RowCol_1 = {img_addr, 10'd102};
  end
  else if (detected_keypoint[1][102]) begin
    filter_input_1_0 = buffer_data_5[839:816];
    filter_input_1_1 = buffer_data_4[839:816];
    filter_input_1_2 = blur5x5_1_dout[839:816];
    current_RowCol_1 = {img_addr, 10'd103};
  end
  else if (detected_keypoint[1][103]) begin
    filter_input_1_0 = buffer_data_5[847:824];
    filter_input_1_1 = buffer_data_4[847:824];
    filter_input_1_2 = blur5x5_1_dout[847:824];
    current_RowCol_1 = {img_addr, 10'd104};
  end
  else if (detected_keypoint[1][104]) begin
    filter_input_1_0 = buffer_data_5[855:832];
    filter_input_1_1 = buffer_data_4[855:832];
    filter_input_1_2 = blur5x5_1_dout[855:832];
    current_RowCol_1 = {img_addr, 10'd105};
  end
  else if (detected_keypoint[1][105]) begin
    filter_input_1_0 = buffer_data_5[863:840];
    filter_input_1_1 = buffer_data_4[863:840];
    filter_input_1_2 = blur5x5_1_dout[863:840];
    current_RowCol_1 = {img_addr, 10'd106};
  end
  else if (detected_keypoint[1][106]) begin
    filter_input_1_0 = buffer_data_5[871:848];
    filter_input_1_1 = buffer_data_4[871:848];
    filter_input_1_2 = blur5x5_1_dout[871:848];
    current_RowCol_1 = {img_addr, 10'd107};
  end
  else if (detected_keypoint[1][107]) begin
    filter_input_1_0 = buffer_data_5[879:856];
    filter_input_1_1 = buffer_data_4[879:856];
    filter_input_1_2 = blur5x5_1_dout[879:856];
    current_RowCol_1 = {img_addr, 10'd108};
  end
  else if (detected_keypoint[1][108]) begin
    filter_input_1_0 = buffer_data_5[887:864];
    filter_input_1_1 = buffer_data_4[887:864];
    filter_input_1_2 = blur5x5_1_dout[887:864];
    current_RowCol_1 = {img_addr, 10'd109};
  end
  else if (detected_keypoint[1][109]) begin
    filter_input_1_0 = buffer_data_5[895:872];
    filter_input_1_1 = buffer_data_4[895:872];
    filter_input_1_2 = blur5x5_1_dout[895:872];
    current_RowCol_1 = {img_addr, 10'd110};
  end
  else if (detected_keypoint[1][110]) begin
    filter_input_1_0 = buffer_data_5[903:880];
    filter_input_1_1 = buffer_data_4[903:880];
    filter_input_1_2 = blur5x5_1_dout[903:880];
    current_RowCol_1 = {img_addr, 10'd111};
  end
  else if (detected_keypoint[1][111]) begin
    filter_input_1_0 = buffer_data_5[911:888];
    filter_input_1_1 = buffer_data_4[911:888];
    filter_input_1_2 = blur5x5_1_dout[911:888];
    current_RowCol_1 = {img_addr, 10'd112};
  end
  else if (detected_keypoint[1][112]) begin
    filter_input_1_0 = buffer_data_5[919:896];
    filter_input_1_1 = buffer_data_4[919:896];
    filter_input_1_2 = blur5x5_1_dout[919:896];
    current_RowCol_1 = {img_addr, 10'd113};
  end
  else if (detected_keypoint[1][113]) begin
    filter_input_1_0 = buffer_data_5[927:904];
    filter_input_1_1 = buffer_data_4[927:904];
    filter_input_1_2 = blur5x5_1_dout[927:904];
    current_RowCol_1 = {img_addr, 10'd114};
  end
  else if (detected_keypoint[1][114]) begin
    filter_input_1_0 = buffer_data_5[935:912];
    filter_input_1_1 = buffer_data_4[935:912];
    filter_input_1_2 = blur5x5_1_dout[935:912];
    current_RowCol_1 = {img_addr, 10'd115};
  end
  else if (detected_keypoint[1][115]) begin
    filter_input_1_0 = buffer_data_5[943:920];
    filter_input_1_1 = buffer_data_4[943:920];
    filter_input_1_2 = blur5x5_1_dout[943:920];
    current_RowCol_1 = {img_addr, 10'd116};
  end
  else if (detected_keypoint[1][116]) begin
    filter_input_1_0 = buffer_data_5[951:928];
    filter_input_1_1 = buffer_data_4[951:928];
    filter_input_1_2 = blur5x5_1_dout[951:928];
    current_RowCol_1 = {img_addr, 10'd117};
  end
  else if (detected_keypoint[1][117]) begin
    filter_input_1_0 = buffer_data_5[959:936];
    filter_input_1_1 = buffer_data_4[959:936];
    filter_input_1_2 = blur5x5_1_dout[959:936];
    current_RowCol_1 = {img_addr, 10'd118};
  end
  else if (detected_keypoint[1][118]) begin
    filter_input_1_0 = buffer_data_5[967:944];
    filter_input_1_1 = buffer_data_4[967:944];
    filter_input_1_2 = blur5x5_1_dout[967:944];
    current_RowCol_1 = {img_addr, 10'd119};
  end
  else if (detected_keypoint[1][119]) begin
    filter_input_1_0 = buffer_data_5[975:952];
    filter_input_1_1 = buffer_data_4[975:952];
    filter_input_1_2 = blur5x5_1_dout[975:952];
    current_RowCol_1 = {img_addr, 10'd120};
  end
  else if (detected_keypoint[1][120]) begin
    filter_input_1_0 = buffer_data_5[983:960];
    filter_input_1_1 = buffer_data_4[983:960];
    filter_input_1_2 = blur5x5_1_dout[983:960];
    current_RowCol_1 = {img_addr, 10'd121};
  end
  else if (detected_keypoint[1][121]) begin
    filter_input_1_0 = buffer_data_5[991:968];
    filter_input_1_1 = buffer_data_4[991:968];
    filter_input_1_2 = blur5x5_1_dout[991:968];
    current_RowCol_1 = {img_addr, 10'd122};
  end
  else if (detected_keypoint[1][122]) begin
    filter_input_1_0 = buffer_data_5[999:976];
    filter_input_1_1 = buffer_data_4[999:976];
    filter_input_1_2 = blur5x5_1_dout[999:976];
    current_RowCol_1 = {img_addr, 10'd123};
  end
  else if (detected_keypoint[1][123]) begin
    filter_input_1_0 = buffer_data_5[1007:984];
    filter_input_1_1 = buffer_data_4[1007:984];
    filter_input_1_2 = blur5x5_1_dout[1007:984];
    current_RowCol_1 = {img_addr, 10'd124};
  end
  else if (detected_keypoint[1][124]) begin
    filter_input_1_0 = buffer_data_5[1015:992];
    filter_input_1_1 = buffer_data_4[1015:992];
    filter_input_1_2 = blur5x5_1_dout[1015:992];
    current_RowCol_1 = {img_addr, 10'd125};
  end
  else if (detected_keypoint[1][125]) begin
    filter_input_1_0 = buffer_data_5[1023:1000];
    filter_input_1_1 = buffer_data_4[1023:1000];
    filter_input_1_2 = blur5x5_1_dout[1023:1000];
    current_RowCol_1 = {img_addr, 10'd126};
  end
  else if (detected_keypoint[1][126]) begin
    filter_input_1_0 = buffer_data_5[1031:1008];
    filter_input_1_1 = buffer_data_4[1031:1008];
    filter_input_1_2 = blur5x5_1_dout[1031:1008];
    current_RowCol_1 = {img_addr, 10'd127};
  end
  else if (detected_keypoint[1][127]) begin
    filter_input_1_0 = buffer_data_5[1039:1016];
    filter_input_1_1 = buffer_data_4[1039:1016];
    filter_input_1_2 = blur5x5_1_dout[1039:1016];
    current_RowCol_1 = {img_addr, 10'd128};
  end
  else if (detected_keypoint[1][128]) begin
    filter_input_1_0 = buffer_data_5[1047:1024];
    filter_input_1_1 = buffer_data_4[1047:1024];
    filter_input_1_2 = blur5x5_1_dout[1047:1024];
    current_RowCol_1 = {img_addr, 10'd129};
  end
  else if (detected_keypoint[1][129]) begin
    filter_input_1_0 = buffer_data_5[1055:1032];
    filter_input_1_1 = buffer_data_4[1055:1032];
    filter_input_1_2 = blur5x5_1_dout[1055:1032];
    current_RowCol_1 = {img_addr, 10'd130};
  end
  else if (detected_keypoint[1][130]) begin
    filter_input_1_0 = buffer_data_5[1063:1040];
    filter_input_1_1 = buffer_data_4[1063:1040];
    filter_input_1_2 = blur5x5_1_dout[1063:1040];
    current_RowCol_1 = {img_addr, 10'd131};
  end
  else if (detected_keypoint[1][131]) begin
    filter_input_1_0 = buffer_data_5[1071:1048];
    filter_input_1_1 = buffer_data_4[1071:1048];
    filter_input_1_2 = blur5x5_1_dout[1071:1048];
    current_RowCol_1 = {img_addr, 10'd132};
  end
  else if (detected_keypoint[1][132]) begin
    filter_input_1_0 = buffer_data_5[1079:1056];
    filter_input_1_1 = buffer_data_4[1079:1056];
    filter_input_1_2 = blur5x5_1_dout[1079:1056];
    current_RowCol_1 = {img_addr, 10'd133};
  end
  else if (detected_keypoint[1][133]) begin
    filter_input_1_0 = buffer_data_5[1087:1064];
    filter_input_1_1 = buffer_data_4[1087:1064];
    filter_input_1_2 = blur5x5_1_dout[1087:1064];
    current_RowCol_1 = {img_addr, 10'd134};
  end
  else if (detected_keypoint[1][134]) begin
    filter_input_1_0 = buffer_data_5[1095:1072];
    filter_input_1_1 = buffer_data_4[1095:1072];
    filter_input_1_2 = blur5x5_1_dout[1095:1072];
    current_RowCol_1 = {img_addr, 10'd135};
  end
  else if (detected_keypoint[1][135]) begin
    filter_input_1_0 = buffer_data_5[1103:1080];
    filter_input_1_1 = buffer_data_4[1103:1080];
    filter_input_1_2 = blur5x5_1_dout[1103:1080];
    current_RowCol_1 = {img_addr, 10'd136};
  end
  else if (detected_keypoint[1][136]) begin
    filter_input_1_0 = buffer_data_5[1111:1088];
    filter_input_1_1 = buffer_data_4[1111:1088];
    filter_input_1_2 = blur5x5_1_dout[1111:1088];
    current_RowCol_1 = {img_addr, 10'd137};
  end
  else if (detected_keypoint[1][137]) begin
    filter_input_1_0 = buffer_data_5[1119:1096];
    filter_input_1_1 = buffer_data_4[1119:1096];
    filter_input_1_2 = blur5x5_1_dout[1119:1096];
    current_RowCol_1 = {img_addr, 10'd138};
  end
  else if (detected_keypoint[1][138]) begin
    filter_input_1_0 = buffer_data_5[1127:1104];
    filter_input_1_1 = buffer_data_4[1127:1104];
    filter_input_1_2 = blur5x5_1_dout[1127:1104];
    current_RowCol_1 = {img_addr, 10'd139};
  end
  else if (detected_keypoint[1][139]) begin
    filter_input_1_0 = buffer_data_5[1135:1112];
    filter_input_1_1 = buffer_data_4[1135:1112];
    filter_input_1_2 = blur5x5_1_dout[1135:1112];
    current_RowCol_1 = {img_addr, 10'd140};
  end
  else if (detected_keypoint[1][140]) begin
    filter_input_1_0 = buffer_data_5[1143:1120];
    filter_input_1_1 = buffer_data_4[1143:1120];
    filter_input_1_2 = blur5x5_1_dout[1143:1120];
    current_RowCol_1 = {img_addr, 10'd141};
  end
  else if (detected_keypoint[1][141]) begin
    filter_input_1_0 = buffer_data_5[1151:1128];
    filter_input_1_1 = buffer_data_4[1151:1128];
    filter_input_1_2 = blur5x5_1_dout[1151:1128];
    current_RowCol_1 = {img_addr, 10'd142};
  end
  else if (detected_keypoint[1][142]) begin
    filter_input_1_0 = buffer_data_5[1159:1136];
    filter_input_1_1 = buffer_data_4[1159:1136];
    filter_input_1_2 = blur5x5_1_dout[1159:1136];
    current_RowCol_1 = {img_addr, 10'd143};
  end
  else if (detected_keypoint[1][143]) begin
    filter_input_1_0 = buffer_data_5[1167:1144];
    filter_input_1_1 = buffer_data_4[1167:1144];
    filter_input_1_2 = blur5x5_1_dout[1167:1144];
    current_RowCol_1 = {img_addr, 10'd144};
  end
  else if (detected_keypoint[1][144]) begin
    filter_input_1_0 = buffer_data_5[1175:1152];
    filter_input_1_1 = buffer_data_4[1175:1152];
    filter_input_1_2 = blur5x5_1_dout[1175:1152];
    current_RowCol_1 = {img_addr, 10'd145};
  end
  else if (detected_keypoint[1][145]) begin
    filter_input_1_0 = buffer_data_5[1183:1160];
    filter_input_1_1 = buffer_data_4[1183:1160];
    filter_input_1_2 = blur5x5_1_dout[1183:1160];
    current_RowCol_1 = {img_addr, 10'd146};
  end
  else if (detected_keypoint[1][146]) begin
    filter_input_1_0 = buffer_data_5[1191:1168];
    filter_input_1_1 = buffer_data_4[1191:1168];
    filter_input_1_2 = blur5x5_1_dout[1191:1168];
    current_RowCol_1 = {img_addr, 10'd147};
  end
  else if (detected_keypoint[1][147]) begin
    filter_input_1_0 = buffer_data_5[1199:1176];
    filter_input_1_1 = buffer_data_4[1199:1176];
    filter_input_1_2 = blur5x5_1_dout[1199:1176];
    current_RowCol_1 = {img_addr, 10'd148};
  end
  else if (detected_keypoint[1][148]) begin
    filter_input_1_0 = buffer_data_5[1207:1184];
    filter_input_1_1 = buffer_data_4[1207:1184];
    filter_input_1_2 = blur5x5_1_dout[1207:1184];
    current_RowCol_1 = {img_addr, 10'd149};
  end
  else if (detected_keypoint[1][149]) begin
    filter_input_1_0 = buffer_data_5[1215:1192];
    filter_input_1_1 = buffer_data_4[1215:1192];
    filter_input_1_2 = blur5x5_1_dout[1215:1192];
    current_RowCol_1 = {img_addr, 10'd150};
  end
  else if (detected_keypoint[1][150]) begin
    filter_input_1_0 = buffer_data_5[1223:1200];
    filter_input_1_1 = buffer_data_4[1223:1200];
    filter_input_1_2 = blur5x5_1_dout[1223:1200];
    current_RowCol_1 = {img_addr, 10'd151};
  end
  else if (detected_keypoint[1][151]) begin
    filter_input_1_0 = buffer_data_5[1231:1208];
    filter_input_1_1 = buffer_data_4[1231:1208];
    filter_input_1_2 = blur5x5_1_dout[1231:1208];
    current_RowCol_1 = {img_addr, 10'd152};
  end
  else if (detected_keypoint[1][152]) begin
    filter_input_1_0 = buffer_data_5[1239:1216];
    filter_input_1_1 = buffer_data_4[1239:1216];
    filter_input_1_2 = blur5x5_1_dout[1239:1216];
    current_RowCol_1 = {img_addr, 10'd153};
  end
  else if (detected_keypoint[1][153]) begin
    filter_input_1_0 = buffer_data_5[1247:1224];
    filter_input_1_1 = buffer_data_4[1247:1224];
    filter_input_1_2 = blur5x5_1_dout[1247:1224];
    current_RowCol_1 = {img_addr, 10'd154};
  end
  else if (detected_keypoint[1][154]) begin
    filter_input_1_0 = buffer_data_5[1255:1232];
    filter_input_1_1 = buffer_data_4[1255:1232];
    filter_input_1_2 = blur5x5_1_dout[1255:1232];
    current_RowCol_1 = {img_addr, 10'd155};
  end
  else if (detected_keypoint[1][155]) begin
    filter_input_1_0 = buffer_data_5[1263:1240];
    filter_input_1_1 = buffer_data_4[1263:1240];
    filter_input_1_2 = blur5x5_1_dout[1263:1240];
    current_RowCol_1 = {img_addr, 10'd156};
  end
  else if (detected_keypoint[1][156]) begin
    filter_input_1_0 = buffer_data_5[1271:1248];
    filter_input_1_1 = buffer_data_4[1271:1248];
    filter_input_1_2 = blur5x5_1_dout[1271:1248];
    current_RowCol_1 = {img_addr, 10'd157};
  end
  else if (detected_keypoint[1][157]) begin
    filter_input_1_0 = buffer_data_5[1279:1256];
    filter_input_1_1 = buffer_data_4[1279:1256];
    filter_input_1_2 = blur5x5_1_dout[1279:1256];
    current_RowCol_1 = {img_addr, 10'd158};
  end
  else if (detected_keypoint[1][158]) begin
    filter_input_1_0 = buffer_data_5[1287:1264];
    filter_input_1_1 = buffer_data_4[1287:1264];
    filter_input_1_2 = blur5x5_1_dout[1287:1264];
    current_RowCol_1 = {img_addr, 10'd159};
  end
  else if (detected_keypoint[1][159]) begin
    filter_input_1_0 = buffer_data_5[1295:1272];
    filter_input_1_1 = buffer_data_4[1295:1272];
    filter_input_1_2 = blur5x5_1_dout[1295:1272];
    current_RowCol_1 = {img_addr, 10'd160};
  end
  else if (detected_keypoint[1][160]) begin
    filter_input_1_0 = buffer_data_5[1303:1280];
    filter_input_1_1 = buffer_data_4[1303:1280];
    filter_input_1_2 = blur5x5_1_dout[1303:1280];
    current_RowCol_1 = {img_addr, 10'd161};
  end
  else if (detected_keypoint[1][161]) begin
    filter_input_1_0 = buffer_data_5[1311:1288];
    filter_input_1_1 = buffer_data_4[1311:1288];
    filter_input_1_2 = blur5x5_1_dout[1311:1288];
    current_RowCol_1 = {img_addr, 10'd162};
  end
  else if (detected_keypoint[1][162]) begin
    filter_input_1_0 = buffer_data_5[1319:1296];
    filter_input_1_1 = buffer_data_4[1319:1296];
    filter_input_1_2 = blur5x5_1_dout[1319:1296];
    current_RowCol_1 = {img_addr, 10'd163};
  end
  else if (detected_keypoint[1][163]) begin
    filter_input_1_0 = buffer_data_5[1327:1304];
    filter_input_1_1 = buffer_data_4[1327:1304];
    filter_input_1_2 = blur5x5_1_dout[1327:1304];
    current_RowCol_1 = {img_addr, 10'd164};
  end
  else if (detected_keypoint[1][164]) begin
    filter_input_1_0 = buffer_data_5[1335:1312];
    filter_input_1_1 = buffer_data_4[1335:1312];
    filter_input_1_2 = blur5x5_1_dout[1335:1312];
    current_RowCol_1 = {img_addr, 10'd165};
  end
  else if (detected_keypoint[1][165]) begin
    filter_input_1_0 = buffer_data_5[1343:1320];
    filter_input_1_1 = buffer_data_4[1343:1320];
    filter_input_1_2 = blur5x5_1_dout[1343:1320];
    current_RowCol_1 = {img_addr, 10'd166};
  end
  else if (detected_keypoint[1][166]) begin
    filter_input_1_0 = buffer_data_5[1351:1328];
    filter_input_1_1 = buffer_data_4[1351:1328];
    filter_input_1_2 = blur5x5_1_dout[1351:1328];
    current_RowCol_1 = {img_addr, 10'd167};
  end
  else if (detected_keypoint[1][167]) begin
    filter_input_1_0 = buffer_data_5[1359:1336];
    filter_input_1_1 = buffer_data_4[1359:1336];
    filter_input_1_2 = blur5x5_1_dout[1359:1336];
    current_RowCol_1 = {img_addr, 10'd168};
  end
  else if (detected_keypoint[1][168]) begin
    filter_input_1_0 = buffer_data_5[1367:1344];
    filter_input_1_1 = buffer_data_4[1367:1344];
    filter_input_1_2 = blur5x5_1_dout[1367:1344];
    current_RowCol_1 = {img_addr, 10'd169};
  end
  else if (detected_keypoint[1][169]) begin
    filter_input_1_0 = buffer_data_5[1375:1352];
    filter_input_1_1 = buffer_data_4[1375:1352];
    filter_input_1_2 = blur5x5_1_dout[1375:1352];
    current_RowCol_1 = {img_addr, 10'd170};
  end
  else if (detected_keypoint[1][170]) begin
    filter_input_1_0 = buffer_data_5[1383:1360];
    filter_input_1_1 = buffer_data_4[1383:1360];
    filter_input_1_2 = blur5x5_1_dout[1383:1360];
    current_RowCol_1 = {img_addr, 10'd171};
  end
  else if (detected_keypoint[1][171]) begin
    filter_input_1_0 = buffer_data_5[1391:1368];
    filter_input_1_1 = buffer_data_4[1391:1368];
    filter_input_1_2 = blur5x5_1_dout[1391:1368];
    current_RowCol_1 = {img_addr, 10'd172};
  end
  else if (detected_keypoint[1][172]) begin
    filter_input_1_0 = buffer_data_5[1399:1376];
    filter_input_1_1 = buffer_data_4[1399:1376];
    filter_input_1_2 = blur5x5_1_dout[1399:1376];
    current_RowCol_1 = {img_addr, 10'd173};
  end
  else if (detected_keypoint[1][173]) begin
    filter_input_1_0 = buffer_data_5[1407:1384];
    filter_input_1_1 = buffer_data_4[1407:1384];
    filter_input_1_2 = blur5x5_1_dout[1407:1384];
    current_RowCol_1 = {img_addr, 10'd174};
  end
  else if (detected_keypoint[1][174]) begin
    filter_input_1_0 = buffer_data_5[1415:1392];
    filter_input_1_1 = buffer_data_4[1415:1392];
    filter_input_1_2 = blur5x5_1_dout[1415:1392];
    current_RowCol_1 = {img_addr, 10'd175};
  end
  else if (detected_keypoint[1][175]) begin
    filter_input_1_0 = buffer_data_5[1423:1400];
    filter_input_1_1 = buffer_data_4[1423:1400];
    filter_input_1_2 = blur5x5_1_dout[1423:1400];
    current_RowCol_1 = {img_addr, 10'd176};
  end
  else if (detected_keypoint[1][176]) begin
    filter_input_1_0 = buffer_data_5[1431:1408];
    filter_input_1_1 = buffer_data_4[1431:1408];
    filter_input_1_2 = blur5x5_1_dout[1431:1408];
    current_RowCol_1 = {img_addr, 10'd177};
  end
  else if (detected_keypoint[1][177]) begin
    filter_input_1_0 = buffer_data_5[1439:1416];
    filter_input_1_1 = buffer_data_4[1439:1416];
    filter_input_1_2 = blur5x5_1_dout[1439:1416];
    current_RowCol_1 = {img_addr, 10'd178};
  end
  else if (detected_keypoint[1][178]) begin
    filter_input_1_0 = buffer_data_5[1447:1424];
    filter_input_1_1 = buffer_data_4[1447:1424];
    filter_input_1_2 = blur5x5_1_dout[1447:1424];
    current_RowCol_1 = {img_addr, 10'd179};
  end
  else if (detected_keypoint[1][179]) begin
    filter_input_1_0 = buffer_data_5[1455:1432];
    filter_input_1_1 = buffer_data_4[1455:1432];
    filter_input_1_2 = blur5x5_1_dout[1455:1432];
    current_RowCol_1 = {img_addr, 10'd180};
  end
  else if (detected_keypoint[1][180]) begin
    filter_input_1_0 = buffer_data_5[1463:1440];
    filter_input_1_1 = buffer_data_4[1463:1440];
    filter_input_1_2 = blur5x5_1_dout[1463:1440];
    current_RowCol_1 = {img_addr, 10'd181};
  end
  else if (detected_keypoint[1][181]) begin
    filter_input_1_0 = buffer_data_5[1471:1448];
    filter_input_1_1 = buffer_data_4[1471:1448];
    filter_input_1_2 = blur5x5_1_dout[1471:1448];
    current_RowCol_1 = {img_addr, 10'd182};
  end
  else if (detected_keypoint[1][182]) begin
    filter_input_1_0 = buffer_data_5[1479:1456];
    filter_input_1_1 = buffer_data_4[1479:1456];
    filter_input_1_2 = blur5x5_1_dout[1479:1456];
    current_RowCol_1 = {img_addr, 10'd183};
  end
  else if (detected_keypoint[1][183]) begin
    filter_input_1_0 = buffer_data_5[1487:1464];
    filter_input_1_1 = buffer_data_4[1487:1464];
    filter_input_1_2 = blur5x5_1_dout[1487:1464];
    current_RowCol_1 = {img_addr, 10'd184};
  end
  else if (detected_keypoint[1][184]) begin
    filter_input_1_0 = buffer_data_5[1495:1472];
    filter_input_1_1 = buffer_data_4[1495:1472];
    filter_input_1_2 = blur5x5_1_dout[1495:1472];
    current_RowCol_1 = {img_addr, 10'd185};
  end
  else if (detected_keypoint[1][185]) begin
    filter_input_1_0 = buffer_data_5[1503:1480];
    filter_input_1_1 = buffer_data_4[1503:1480];
    filter_input_1_2 = blur5x5_1_dout[1503:1480];
    current_RowCol_1 = {img_addr, 10'd186};
  end
  else if (detected_keypoint[1][186]) begin
    filter_input_1_0 = buffer_data_5[1511:1488];
    filter_input_1_1 = buffer_data_4[1511:1488];
    filter_input_1_2 = blur5x5_1_dout[1511:1488];
    current_RowCol_1 = {img_addr, 10'd187};
  end
  else if (detected_keypoint[1][187]) begin
    filter_input_1_0 = buffer_data_5[1519:1496];
    filter_input_1_1 = buffer_data_4[1519:1496];
    filter_input_1_2 = blur5x5_1_dout[1519:1496];
    current_RowCol_1 = {img_addr, 10'd188};
  end
  else if (detected_keypoint[1][188]) begin
    filter_input_1_0 = buffer_data_5[1527:1504];
    filter_input_1_1 = buffer_data_4[1527:1504];
    filter_input_1_2 = blur5x5_1_dout[1527:1504];
    current_RowCol_1 = {img_addr, 10'd189};
  end
  else if (detected_keypoint[1][189]) begin
    filter_input_1_0 = buffer_data_5[1535:1512];
    filter_input_1_1 = buffer_data_4[1535:1512];
    filter_input_1_2 = blur5x5_1_dout[1535:1512];
    current_RowCol_1 = {img_addr, 10'd190};
  end
  else if (detected_keypoint[1][190]) begin
    filter_input_1_0 = buffer_data_5[1543:1520];
    filter_input_1_1 = buffer_data_4[1543:1520];
    filter_input_1_2 = blur5x5_1_dout[1543:1520];
    current_RowCol_1 = {img_addr, 10'd191};
  end
  else if (detected_keypoint[1][191]) begin
    filter_input_1_0 = buffer_data_5[1551:1528];
    filter_input_1_1 = buffer_data_4[1551:1528];
    filter_input_1_2 = blur5x5_1_dout[1551:1528];
    current_RowCol_1 = {img_addr, 10'd192};
  end
  else if (detected_keypoint[1][192]) begin
    filter_input_1_0 = buffer_data_5[1559:1536];
    filter_input_1_1 = buffer_data_4[1559:1536];
    filter_input_1_2 = blur5x5_1_dout[1559:1536];
    current_RowCol_1 = {img_addr, 10'd193};
  end
  else if (detected_keypoint[1][193]) begin
    filter_input_1_0 = buffer_data_5[1567:1544];
    filter_input_1_1 = buffer_data_4[1567:1544];
    filter_input_1_2 = blur5x5_1_dout[1567:1544];
    current_RowCol_1 = {img_addr, 10'd194};
  end
  else if (detected_keypoint[1][194]) begin
    filter_input_1_0 = buffer_data_5[1575:1552];
    filter_input_1_1 = buffer_data_4[1575:1552];
    filter_input_1_2 = blur5x5_1_dout[1575:1552];
    current_RowCol_1 = {img_addr, 10'd195};
  end
  else if (detected_keypoint[1][195]) begin
    filter_input_1_0 = buffer_data_5[1583:1560];
    filter_input_1_1 = buffer_data_4[1583:1560];
    filter_input_1_2 = blur5x5_1_dout[1583:1560];
    current_RowCol_1 = {img_addr, 10'd196};
  end
  else if (detected_keypoint[1][196]) begin
    filter_input_1_0 = buffer_data_5[1591:1568];
    filter_input_1_1 = buffer_data_4[1591:1568];
    filter_input_1_2 = blur5x5_1_dout[1591:1568];
    current_RowCol_1 = {img_addr, 10'd197};
  end
  else if (detected_keypoint[1][197]) begin
    filter_input_1_0 = buffer_data_5[1599:1576];
    filter_input_1_1 = buffer_data_4[1599:1576];
    filter_input_1_2 = blur5x5_1_dout[1599:1576];
    current_RowCol_1 = {img_addr, 10'd198};
  end
  else if (detected_keypoint[1][198]) begin
    filter_input_1_0 = buffer_data_5[1607:1584];
    filter_input_1_1 = buffer_data_4[1607:1584];
    filter_input_1_2 = blur5x5_1_dout[1607:1584];
    current_RowCol_1 = {img_addr, 10'd199};
  end
  else if (detected_keypoint[1][199]) begin
    filter_input_1_0 = buffer_data_5[1615:1592];
    filter_input_1_1 = buffer_data_4[1615:1592];
    filter_input_1_2 = blur5x5_1_dout[1615:1592];
    current_RowCol_1 = {img_addr, 10'd200};
  end
  else if (detected_keypoint[1][200]) begin
    filter_input_1_0 = buffer_data_5[1623:1600];
    filter_input_1_1 = buffer_data_4[1623:1600];
    filter_input_1_2 = blur5x5_1_dout[1623:1600];
    current_RowCol_1 = {img_addr, 10'd201};
  end
  else if (detected_keypoint[1][201]) begin
    filter_input_1_0 = buffer_data_5[1631:1608];
    filter_input_1_1 = buffer_data_4[1631:1608];
    filter_input_1_2 = blur5x5_1_dout[1631:1608];
    current_RowCol_1 = {img_addr, 10'd202};
  end
  else if (detected_keypoint[1][202]) begin
    filter_input_1_0 = buffer_data_5[1639:1616];
    filter_input_1_1 = buffer_data_4[1639:1616];
    filter_input_1_2 = blur5x5_1_dout[1639:1616];
    current_RowCol_1 = {img_addr, 10'd203};
  end
  else if (detected_keypoint[1][203]) begin
    filter_input_1_0 = buffer_data_5[1647:1624];
    filter_input_1_1 = buffer_data_4[1647:1624];
    filter_input_1_2 = blur5x5_1_dout[1647:1624];
    current_RowCol_1 = {img_addr, 10'd204};
  end
  else if (detected_keypoint[1][204]) begin
    filter_input_1_0 = buffer_data_5[1655:1632];
    filter_input_1_1 = buffer_data_4[1655:1632];
    filter_input_1_2 = blur5x5_1_dout[1655:1632];
    current_RowCol_1 = {img_addr, 10'd205};
  end
  else if (detected_keypoint[1][205]) begin
    filter_input_1_0 = buffer_data_5[1663:1640];
    filter_input_1_1 = buffer_data_4[1663:1640];
    filter_input_1_2 = blur5x5_1_dout[1663:1640];
    current_RowCol_1 = {img_addr, 10'd206};
  end
  else if (detected_keypoint[1][206]) begin
    filter_input_1_0 = buffer_data_5[1671:1648];
    filter_input_1_1 = buffer_data_4[1671:1648];
    filter_input_1_2 = blur5x5_1_dout[1671:1648];
    current_RowCol_1 = {img_addr, 10'd207};
  end
  else if (detected_keypoint[1][207]) begin
    filter_input_1_0 = buffer_data_5[1679:1656];
    filter_input_1_1 = buffer_data_4[1679:1656];
    filter_input_1_2 = blur5x5_1_dout[1679:1656];
    current_RowCol_1 = {img_addr, 10'd208};
  end
  else if (detected_keypoint[1][208]) begin
    filter_input_1_0 = buffer_data_5[1687:1664];
    filter_input_1_1 = buffer_data_4[1687:1664];
    filter_input_1_2 = blur5x5_1_dout[1687:1664];
    current_RowCol_1 = {img_addr, 10'd209};
  end
  else if (detected_keypoint[1][209]) begin
    filter_input_1_0 = buffer_data_5[1695:1672];
    filter_input_1_1 = buffer_data_4[1695:1672];
    filter_input_1_2 = blur5x5_1_dout[1695:1672];
    current_RowCol_1 = {img_addr, 10'd210};
  end
  else if (detected_keypoint[1][210]) begin
    filter_input_1_0 = buffer_data_5[1703:1680];
    filter_input_1_1 = buffer_data_4[1703:1680];
    filter_input_1_2 = blur5x5_1_dout[1703:1680];
    current_RowCol_1 = {img_addr, 10'd211};
  end
  else if (detected_keypoint[1][211]) begin
    filter_input_1_0 = buffer_data_5[1711:1688];
    filter_input_1_1 = buffer_data_4[1711:1688];
    filter_input_1_2 = blur5x5_1_dout[1711:1688];
    current_RowCol_1 = {img_addr, 10'd212};
  end
  else if (detected_keypoint[1][212]) begin
    filter_input_1_0 = buffer_data_5[1719:1696];
    filter_input_1_1 = buffer_data_4[1719:1696];
    filter_input_1_2 = blur5x5_1_dout[1719:1696];
    current_RowCol_1 = {img_addr, 10'd213};
  end
  else if (detected_keypoint[1][213]) begin
    filter_input_1_0 = buffer_data_5[1727:1704];
    filter_input_1_1 = buffer_data_4[1727:1704];
    filter_input_1_2 = blur5x5_1_dout[1727:1704];
    current_RowCol_1 = {img_addr, 10'd214};
  end
  else if (detected_keypoint[1][214]) begin
    filter_input_1_0 = buffer_data_5[1735:1712];
    filter_input_1_1 = buffer_data_4[1735:1712];
    filter_input_1_2 = blur5x5_1_dout[1735:1712];
    current_RowCol_1 = {img_addr, 10'd215};
  end
  else if (detected_keypoint[1][215]) begin
    filter_input_1_0 = buffer_data_5[1743:1720];
    filter_input_1_1 = buffer_data_4[1743:1720];
    filter_input_1_2 = blur5x5_1_dout[1743:1720];
    current_RowCol_1 = {img_addr, 10'd216};
  end
  else if (detected_keypoint[1][216]) begin
    filter_input_1_0 = buffer_data_5[1751:1728];
    filter_input_1_1 = buffer_data_4[1751:1728];
    filter_input_1_2 = blur5x5_1_dout[1751:1728];
    current_RowCol_1 = {img_addr, 10'd217};
  end
  else if (detected_keypoint[1][217]) begin
    filter_input_1_0 = buffer_data_5[1759:1736];
    filter_input_1_1 = buffer_data_4[1759:1736];
    filter_input_1_2 = blur5x5_1_dout[1759:1736];
    current_RowCol_1 = {img_addr, 10'd218};
  end
  else if (detected_keypoint[1][218]) begin
    filter_input_1_0 = buffer_data_5[1767:1744];
    filter_input_1_1 = buffer_data_4[1767:1744];
    filter_input_1_2 = blur5x5_1_dout[1767:1744];
    current_RowCol_1 = {img_addr, 10'd219};
  end
  else if (detected_keypoint[1][219]) begin
    filter_input_1_0 = buffer_data_5[1775:1752];
    filter_input_1_1 = buffer_data_4[1775:1752];
    filter_input_1_2 = blur5x5_1_dout[1775:1752];
    current_RowCol_1 = {img_addr, 10'd220};
  end
  else if (detected_keypoint[1][220]) begin
    filter_input_1_0 = buffer_data_5[1783:1760];
    filter_input_1_1 = buffer_data_4[1783:1760];
    filter_input_1_2 = blur5x5_1_dout[1783:1760];
    current_RowCol_1 = {img_addr, 10'd221};
  end
  else if (detected_keypoint[1][221]) begin
    filter_input_1_0 = buffer_data_5[1791:1768];
    filter_input_1_1 = buffer_data_4[1791:1768];
    filter_input_1_2 = blur5x5_1_dout[1791:1768];
    current_RowCol_1 = {img_addr, 10'd222};
  end
  else if (detected_keypoint[1][222]) begin
    filter_input_1_0 = buffer_data_5[1799:1776];
    filter_input_1_1 = buffer_data_4[1799:1776];
    filter_input_1_2 = blur5x5_1_dout[1799:1776];
    current_RowCol_1 = {img_addr, 10'd223};
  end
  else if (detected_keypoint[1][223]) begin
    filter_input_1_0 = buffer_data_5[1807:1784];
    filter_input_1_1 = buffer_data_4[1807:1784];
    filter_input_1_2 = blur5x5_1_dout[1807:1784];
    current_RowCol_1 = {img_addr, 10'd224};
  end
  else if (detected_keypoint[1][224]) begin
    filter_input_1_0 = buffer_data_5[1815:1792];
    filter_input_1_1 = buffer_data_4[1815:1792];
    filter_input_1_2 = blur5x5_1_dout[1815:1792];
    current_RowCol_1 = {img_addr, 10'd225};
  end
  else if (detected_keypoint[1][225]) begin
    filter_input_1_0 = buffer_data_5[1823:1800];
    filter_input_1_1 = buffer_data_4[1823:1800];
    filter_input_1_2 = blur5x5_1_dout[1823:1800];
    current_RowCol_1 = {img_addr, 10'd226};
  end
  else if (detected_keypoint[1][226]) begin
    filter_input_1_0 = buffer_data_5[1831:1808];
    filter_input_1_1 = buffer_data_4[1831:1808];
    filter_input_1_2 = blur5x5_1_dout[1831:1808];
    current_RowCol_1 = {img_addr, 10'd227};
  end
  else if (detected_keypoint[1][227]) begin
    filter_input_1_0 = buffer_data_5[1839:1816];
    filter_input_1_1 = buffer_data_4[1839:1816];
    filter_input_1_2 = blur5x5_1_dout[1839:1816];
    current_RowCol_1 = {img_addr, 10'd228};
  end
  else if (detected_keypoint[1][228]) begin
    filter_input_1_0 = buffer_data_5[1847:1824];
    filter_input_1_1 = buffer_data_4[1847:1824];
    filter_input_1_2 = blur5x5_1_dout[1847:1824];
    current_RowCol_1 = {img_addr, 10'd229};
  end
  else if (detected_keypoint[1][229]) begin
    filter_input_1_0 = buffer_data_5[1855:1832];
    filter_input_1_1 = buffer_data_4[1855:1832];
    filter_input_1_2 = blur5x5_1_dout[1855:1832];
    current_RowCol_1 = {img_addr, 10'd230};
  end
  else if (detected_keypoint[1][230]) begin
    filter_input_1_0 = buffer_data_5[1863:1840];
    filter_input_1_1 = buffer_data_4[1863:1840];
    filter_input_1_2 = blur5x5_1_dout[1863:1840];
    current_RowCol_1 = {img_addr, 10'd231};
  end
  else if (detected_keypoint[1][231]) begin
    filter_input_1_0 = buffer_data_5[1871:1848];
    filter_input_1_1 = buffer_data_4[1871:1848];
    filter_input_1_2 = blur5x5_1_dout[1871:1848];
    current_RowCol_1 = {img_addr, 10'd232};
  end
  else if (detected_keypoint[1][232]) begin
    filter_input_1_0 = buffer_data_5[1879:1856];
    filter_input_1_1 = buffer_data_4[1879:1856];
    filter_input_1_2 = blur5x5_1_dout[1879:1856];
    current_RowCol_1 = {img_addr, 10'd233};
  end
  else if (detected_keypoint[1][233]) begin
    filter_input_1_0 = buffer_data_5[1887:1864];
    filter_input_1_1 = buffer_data_4[1887:1864];
    filter_input_1_2 = blur5x5_1_dout[1887:1864];
    current_RowCol_1 = {img_addr, 10'd234};
  end
  else if (detected_keypoint[1][234]) begin
    filter_input_1_0 = buffer_data_5[1895:1872];
    filter_input_1_1 = buffer_data_4[1895:1872];
    filter_input_1_2 = blur5x5_1_dout[1895:1872];
    current_RowCol_1 = {img_addr, 10'd235};
  end
  else if (detected_keypoint[1][235]) begin
    filter_input_1_0 = buffer_data_5[1903:1880];
    filter_input_1_1 = buffer_data_4[1903:1880];
    filter_input_1_2 = blur5x5_1_dout[1903:1880];
    current_RowCol_1 = {img_addr, 10'd236};
  end
  else if (detected_keypoint[1][236]) begin
    filter_input_1_0 = buffer_data_5[1911:1888];
    filter_input_1_1 = buffer_data_4[1911:1888];
    filter_input_1_2 = blur5x5_1_dout[1911:1888];
    current_RowCol_1 = {img_addr, 10'd237};
  end
  else if (detected_keypoint[1][237]) begin
    filter_input_1_0 = buffer_data_5[1919:1896];
    filter_input_1_1 = buffer_data_4[1919:1896];
    filter_input_1_2 = blur5x5_1_dout[1919:1896];
    current_RowCol_1 = {img_addr, 10'd238};
  end
  else if (detected_keypoint[1][238]) begin
    filter_input_1_0 = buffer_data_5[1927:1904];
    filter_input_1_1 = buffer_data_4[1927:1904];
    filter_input_1_2 = blur5x5_1_dout[1927:1904];
    current_RowCol_1 = {img_addr, 10'd239};
  end
  else if (detected_keypoint[1][239]) begin
    filter_input_1_0 = buffer_data_5[1935:1912];
    filter_input_1_1 = buffer_data_4[1935:1912];
    filter_input_1_2 = blur5x5_1_dout[1935:1912];
    current_RowCol_1 = {img_addr, 10'd240};
  end
  else if (detected_keypoint[1][240]) begin
    filter_input_1_0 = buffer_data_5[1943:1920];
    filter_input_1_1 = buffer_data_4[1943:1920];
    filter_input_1_2 = blur5x5_1_dout[1943:1920];
    current_RowCol_1 = {img_addr, 10'd241};
  end
  else if (detected_keypoint[1][241]) begin
    filter_input_1_0 = buffer_data_5[1951:1928];
    filter_input_1_1 = buffer_data_4[1951:1928];
    filter_input_1_2 = blur5x5_1_dout[1951:1928];
    current_RowCol_1 = {img_addr, 10'd242};
  end
  else if (detected_keypoint[1][242]) begin
    filter_input_1_0 = buffer_data_5[1959:1936];
    filter_input_1_1 = buffer_data_4[1959:1936];
    filter_input_1_2 = blur5x5_1_dout[1959:1936];
    current_RowCol_1 = {img_addr, 10'd243};
  end
  else if (detected_keypoint[1][243]) begin
    filter_input_1_0 = buffer_data_5[1967:1944];
    filter_input_1_1 = buffer_data_4[1967:1944];
    filter_input_1_2 = blur5x5_1_dout[1967:1944];
    current_RowCol_1 = {img_addr, 10'd244};
  end
  else if (detected_keypoint[1][244]) begin
    filter_input_1_0 = buffer_data_5[1975:1952];
    filter_input_1_1 = buffer_data_4[1975:1952];
    filter_input_1_2 = blur5x5_1_dout[1975:1952];
    current_RowCol_1 = {img_addr, 10'd245};
  end
  else if (detected_keypoint[1][245]) begin
    filter_input_1_0 = buffer_data_5[1983:1960];
    filter_input_1_1 = buffer_data_4[1983:1960];
    filter_input_1_2 = blur5x5_1_dout[1983:1960];
    current_RowCol_1 = {img_addr, 10'd246};
  end
  else if (detected_keypoint[1][246]) begin
    filter_input_1_0 = buffer_data_5[1991:1968];
    filter_input_1_1 = buffer_data_4[1991:1968];
    filter_input_1_2 = blur5x5_1_dout[1991:1968];
    current_RowCol_1 = {img_addr, 10'd247};
  end
  else if (detected_keypoint[1][247]) begin
    filter_input_1_0 = buffer_data_5[1999:1976];
    filter_input_1_1 = buffer_data_4[1999:1976];
    filter_input_1_2 = blur5x5_1_dout[1999:1976];
    current_RowCol_1 = {img_addr, 10'd248};
  end
  else if (detected_keypoint[1][248]) begin
    filter_input_1_0 = buffer_data_5[2007:1984];
    filter_input_1_1 = buffer_data_4[2007:1984];
    filter_input_1_2 = blur5x5_1_dout[2007:1984];
    current_RowCol_1 = {img_addr, 10'd249};
  end
  else if (detected_keypoint[1][249]) begin
    filter_input_1_0 = buffer_data_5[2015:1992];
    filter_input_1_1 = buffer_data_4[2015:1992];
    filter_input_1_2 = blur5x5_1_dout[2015:1992];
    current_RowCol_1 = {img_addr, 10'd250};
  end
  else if (detected_keypoint[1][250]) begin
    filter_input_1_0 = buffer_data_5[2023:2000];
    filter_input_1_1 = buffer_data_4[2023:2000];
    filter_input_1_2 = blur5x5_1_dout[2023:2000];
    current_RowCol_1 = {img_addr, 10'd251};
  end
  else if (detected_keypoint[1][251]) begin
    filter_input_1_0 = buffer_data_5[2031:2008];
    filter_input_1_1 = buffer_data_4[2031:2008];
    filter_input_1_2 = blur5x5_1_dout[2031:2008];
    current_RowCol_1 = {img_addr, 10'd252};
  end
  else if (detected_keypoint[1][252]) begin
    filter_input_1_0 = buffer_data_5[2039:2016];
    filter_input_1_1 = buffer_data_4[2039:2016];
    filter_input_1_2 = blur5x5_1_dout[2039:2016];
    current_RowCol_1 = {img_addr, 10'd253};
  end
  else if (detected_keypoint[1][253]) begin
    filter_input_1_0 = buffer_data_5[2047:2024];
    filter_input_1_1 = buffer_data_4[2047:2024];
    filter_input_1_2 = blur5x5_1_dout[2047:2024];
    current_RowCol_1 = {img_addr, 10'd254};
  end
  else if (detected_keypoint[1][254]) begin
    filter_input_1_0 = buffer_data_5[2055:2032];
    filter_input_1_1 = buffer_data_4[2055:2032];
    filter_input_1_2 = blur5x5_1_dout[2055:2032];
    current_RowCol_1 = {img_addr, 10'd255};
  end
  else if (detected_keypoint[1][255]) begin
    filter_input_1_0 = buffer_data_5[2063:2040];
    filter_input_1_1 = buffer_data_4[2063:2040];
    filter_input_1_2 = blur5x5_1_dout[2063:2040];
    current_RowCol_1 = {img_addr, 10'd256};
  end
  else if (detected_keypoint[1][256]) begin
    filter_input_1_0 = buffer_data_5[2071:2048];
    filter_input_1_1 = buffer_data_4[2071:2048];
    filter_input_1_2 = blur5x5_1_dout[2071:2048];
    current_RowCol_1 = {img_addr, 10'd257};
  end
  else if (detected_keypoint[1][257]) begin
    filter_input_1_0 = buffer_data_5[2079:2056];
    filter_input_1_1 = buffer_data_4[2079:2056];
    filter_input_1_2 = blur5x5_1_dout[2079:2056];
    current_RowCol_1 = {img_addr, 10'd258};
  end
  else if (detected_keypoint[1][258]) begin
    filter_input_1_0 = buffer_data_5[2087:2064];
    filter_input_1_1 = buffer_data_4[2087:2064];
    filter_input_1_2 = blur5x5_1_dout[2087:2064];
    current_RowCol_1 = {img_addr, 10'd259};
  end
  else if (detected_keypoint[1][259]) begin
    filter_input_1_0 = buffer_data_5[2095:2072];
    filter_input_1_1 = buffer_data_4[2095:2072];
    filter_input_1_2 = blur5x5_1_dout[2095:2072];
    current_RowCol_1 = {img_addr, 10'd260};
  end
  else if (detected_keypoint[1][260]) begin
    filter_input_1_0 = buffer_data_5[2103:2080];
    filter_input_1_1 = buffer_data_4[2103:2080];
    filter_input_1_2 = blur5x5_1_dout[2103:2080];
    current_RowCol_1 = {img_addr, 10'd261};
  end
  else if (detected_keypoint[1][261]) begin
    filter_input_1_0 = buffer_data_5[2111:2088];
    filter_input_1_1 = buffer_data_4[2111:2088];
    filter_input_1_2 = blur5x5_1_dout[2111:2088];
    current_RowCol_1 = {img_addr, 10'd262};
  end
  else if (detected_keypoint[1][262]) begin
    filter_input_1_0 = buffer_data_5[2119:2096];
    filter_input_1_1 = buffer_data_4[2119:2096];
    filter_input_1_2 = blur5x5_1_dout[2119:2096];
    current_RowCol_1 = {img_addr, 10'd263};
  end
  else if (detected_keypoint[1][263]) begin
    filter_input_1_0 = buffer_data_5[2127:2104];
    filter_input_1_1 = buffer_data_4[2127:2104];
    filter_input_1_2 = blur5x5_1_dout[2127:2104];
    current_RowCol_1 = {img_addr, 10'd264};
  end
  else if (detected_keypoint[1][264]) begin
    filter_input_1_0 = buffer_data_5[2135:2112];
    filter_input_1_1 = buffer_data_4[2135:2112];
    filter_input_1_2 = blur5x5_1_dout[2135:2112];
    current_RowCol_1 = {img_addr, 10'd265};
  end
  else if (detected_keypoint[1][265]) begin
    filter_input_1_0 = buffer_data_5[2143:2120];
    filter_input_1_1 = buffer_data_4[2143:2120];
    filter_input_1_2 = blur5x5_1_dout[2143:2120];
    current_RowCol_1 = {img_addr, 10'd266};
  end
  else if (detected_keypoint[1][266]) begin
    filter_input_1_0 = buffer_data_5[2151:2128];
    filter_input_1_1 = buffer_data_4[2151:2128];
    filter_input_1_2 = blur5x5_1_dout[2151:2128];
    current_RowCol_1 = {img_addr, 10'd267};
  end
  else if (detected_keypoint[1][267]) begin
    filter_input_1_0 = buffer_data_5[2159:2136];
    filter_input_1_1 = buffer_data_4[2159:2136];
    filter_input_1_2 = blur5x5_1_dout[2159:2136];
    current_RowCol_1 = {img_addr, 10'd268};
  end
  else if (detected_keypoint[1][268]) begin
    filter_input_1_0 = buffer_data_5[2167:2144];
    filter_input_1_1 = buffer_data_4[2167:2144];
    filter_input_1_2 = blur5x5_1_dout[2167:2144];
    current_RowCol_1 = {img_addr, 10'd269};
  end
  else if (detected_keypoint[1][269]) begin
    filter_input_1_0 = buffer_data_5[2175:2152];
    filter_input_1_1 = buffer_data_4[2175:2152];
    filter_input_1_2 = blur5x5_1_dout[2175:2152];
    current_RowCol_1 = {img_addr, 10'd270};
  end
  else if (detected_keypoint[1][270]) begin
    filter_input_1_0 = buffer_data_5[2183:2160];
    filter_input_1_1 = buffer_data_4[2183:2160];
    filter_input_1_2 = blur5x5_1_dout[2183:2160];
    current_RowCol_1 = {img_addr, 10'd271};
  end
  else if (detected_keypoint[1][271]) begin
    filter_input_1_0 = buffer_data_5[2191:2168];
    filter_input_1_1 = buffer_data_4[2191:2168];
    filter_input_1_2 = blur5x5_1_dout[2191:2168];
    current_RowCol_1 = {img_addr, 10'd272};
  end
  else if (detected_keypoint[1][272]) begin
    filter_input_1_0 = buffer_data_5[2199:2176];
    filter_input_1_1 = buffer_data_4[2199:2176];
    filter_input_1_2 = blur5x5_1_dout[2199:2176];
    current_RowCol_1 = {img_addr, 10'd273};
  end
  else if (detected_keypoint[1][273]) begin
    filter_input_1_0 = buffer_data_5[2207:2184];
    filter_input_1_1 = buffer_data_4[2207:2184];
    filter_input_1_2 = blur5x5_1_dout[2207:2184];
    current_RowCol_1 = {img_addr, 10'd274};
  end
  else if (detected_keypoint[1][274]) begin
    filter_input_1_0 = buffer_data_5[2215:2192];
    filter_input_1_1 = buffer_data_4[2215:2192];
    filter_input_1_2 = blur5x5_1_dout[2215:2192];
    current_RowCol_1 = {img_addr, 10'd275};
  end
  else if (detected_keypoint[1][275]) begin
    filter_input_1_0 = buffer_data_5[2223:2200];
    filter_input_1_1 = buffer_data_4[2223:2200];
    filter_input_1_2 = blur5x5_1_dout[2223:2200];
    current_RowCol_1 = {img_addr, 10'd276};
  end
  else if (detected_keypoint[1][276]) begin
    filter_input_1_0 = buffer_data_5[2231:2208];
    filter_input_1_1 = buffer_data_4[2231:2208];
    filter_input_1_2 = blur5x5_1_dout[2231:2208];
    current_RowCol_1 = {img_addr, 10'd277};
  end
  else if (detected_keypoint[1][277]) begin
    filter_input_1_0 = buffer_data_5[2239:2216];
    filter_input_1_1 = buffer_data_4[2239:2216];
    filter_input_1_2 = blur5x5_1_dout[2239:2216];
    current_RowCol_1 = {img_addr, 10'd278};
  end
  else if (detected_keypoint[1][278]) begin
    filter_input_1_0 = buffer_data_5[2247:2224];
    filter_input_1_1 = buffer_data_4[2247:2224];
    filter_input_1_2 = blur5x5_1_dout[2247:2224];
    current_RowCol_1 = {img_addr, 10'd279};
  end
  else if (detected_keypoint[1][279]) begin
    filter_input_1_0 = buffer_data_5[2255:2232];
    filter_input_1_1 = buffer_data_4[2255:2232];
    filter_input_1_2 = blur5x5_1_dout[2255:2232];
    current_RowCol_1 = {img_addr, 10'd280};
  end
  else if (detected_keypoint[1][280]) begin
    filter_input_1_0 = buffer_data_5[2263:2240];
    filter_input_1_1 = buffer_data_4[2263:2240];
    filter_input_1_2 = blur5x5_1_dout[2263:2240];
    current_RowCol_1 = {img_addr, 10'd281};
  end
  else if (detected_keypoint[1][281]) begin
    filter_input_1_0 = buffer_data_5[2271:2248];
    filter_input_1_1 = buffer_data_4[2271:2248];
    filter_input_1_2 = blur5x5_1_dout[2271:2248];
    current_RowCol_1 = {img_addr, 10'd282};
  end
  else if (detected_keypoint[1][282]) begin
    filter_input_1_0 = buffer_data_5[2279:2256];
    filter_input_1_1 = buffer_data_4[2279:2256];
    filter_input_1_2 = blur5x5_1_dout[2279:2256];
    current_RowCol_1 = {img_addr, 10'd283};
  end
  else if (detected_keypoint[1][283]) begin
    filter_input_1_0 = buffer_data_5[2287:2264];
    filter_input_1_1 = buffer_data_4[2287:2264];
    filter_input_1_2 = blur5x5_1_dout[2287:2264];
    current_RowCol_1 = {img_addr, 10'd284};
  end
  else if (detected_keypoint[1][284]) begin
    filter_input_1_0 = buffer_data_5[2295:2272];
    filter_input_1_1 = buffer_data_4[2295:2272];
    filter_input_1_2 = blur5x5_1_dout[2295:2272];
    current_RowCol_1 = {img_addr, 10'd285};
  end
  else if (detected_keypoint[1][285]) begin
    filter_input_1_0 = buffer_data_5[2303:2280];
    filter_input_1_1 = buffer_data_4[2303:2280];
    filter_input_1_2 = blur5x5_1_dout[2303:2280];
    current_RowCol_1 = {img_addr, 10'd286};
  end
  else if (detected_keypoint[1][286]) begin
    filter_input_1_0 = buffer_data_5[2311:2288];
    filter_input_1_1 = buffer_data_4[2311:2288];
    filter_input_1_2 = blur5x5_1_dout[2311:2288];
    current_RowCol_1 = {img_addr, 10'd287};
  end
  else if (detected_keypoint[1][287]) begin
    filter_input_1_0 = buffer_data_5[2319:2296];
    filter_input_1_1 = buffer_data_4[2319:2296];
    filter_input_1_2 = blur5x5_1_dout[2319:2296];
    current_RowCol_1 = {img_addr, 10'd288};
  end
  else if (detected_keypoint[1][288]) begin
    filter_input_1_0 = buffer_data_5[2327:2304];
    filter_input_1_1 = buffer_data_4[2327:2304];
    filter_input_1_2 = blur5x5_1_dout[2327:2304];
    current_RowCol_1 = {img_addr, 10'd289};
  end
  else if (detected_keypoint[1][289]) begin
    filter_input_1_0 = buffer_data_5[2335:2312];
    filter_input_1_1 = buffer_data_4[2335:2312];
    filter_input_1_2 = blur5x5_1_dout[2335:2312];
    current_RowCol_1 = {img_addr, 10'd290};
  end
  else if (detected_keypoint[1][290]) begin
    filter_input_1_0 = buffer_data_5[2343:2320];
    filter_input_1_1 = buffer_data_4[2343:2320];
    filter_input_1_2 = blur5x5_1_dout[2343:2320];
    current_RowCol_1 = {img_addr, 10'd291};
  end
  else if (detected_keypoint[1][291]) begin
    filter_input_1_0 = buffer_data_5[2351:2328];
    filter_input_1_1 = buffer_data_4[2351:2328];
    filter_input_1_2 = blur5x5_1_dout[2351:2328];
    current_RowCol_1 = {img_addr, 10'd292};
  end
  else if (detected_keypoint[1][292]) begin
    filter_input_1_0 = buffer_data_5[2359:2336];
    filter_input_1_1 = buffer_data_4[2359:2336];
    filter_input_1_2 = blur5x5_1_dout[2359:2336];
    current_RowCol_1 = {img_addr, 10'd293};
  end
  else if (detected_keypoint[1][293]) begin
    filter_input_1_0 = buffer_data_5[2367:2344];
    filter_input_1_1 = buffer_data_4[2367:2344];
    filter_input_1_2 = blur5x5_1_dout[2367:2344];
    current_RowCol_1 = {img_addr, 10'd294};
  end
  else if (detected_keypoint[1][294]) begin
    filter_input_1_0 = buffer_data_5[2375:2352];
    filter_input_1_1 = buffer_data_4[2375:2352];
    filter_input_1_2 = blur5x5_1_dout[2375:2352];
    current_RowCol_1 = {img_addr, 10'd295};
  end
  else if (detected_keypoint[1][295]) begin
    filter_input_1_0 = buffer_data_5[2383:2360];
    filter_input_1_1 = buffer_data_4[2383:2360];
    filter_input_1_2 = blur5x5_1_dout[2383:2360];
    current_RowCol_1 = {img_addr, 10'd296};
  end
  else if (detected_keypoint[1][296]) begin
    filter_input_1_0 = buffer_data_5[2391:2368];
    filter_input_1_1 = buffer_data_4[2391:2368];
    filter_input_1_2 = blur5x5_1_dout[2391:2368];
    current_RowCol_1 = {img_addr, 10'd297};
  end
  else if (detected_keypoint[1][297]) begin
    filter_input_1_0 = buffer_data_5[2399:2376];
    filter_input_1_1 = buffer_data_4[2399:2376];
    filter_input_1_2 = blur5x5_1_dout[2399:2376];
    current_RowCol_1 = {img_addr, 10'd298};
  end
  else if (detected_keypoint[1][298]) begin
    filter_input_1_0 = buffer_data_5[2407:2384];
    filter_input_1_1 = buffer_data_4[2407:2384];
    filter_input_1_2 = blur5x5_1_dout[2407:2384];
    current_RowCol_1 = {img_addr, 10'd299};
  end
  else if (detected_keypoint[1][299]) begin
    filter_input_1_0 = buffer_data_5[2415:2392];
    filter_input_1_1 = buffer_data_4[2415:2392];
    filter_input_1_2 = blur5x5_1_dout[2415:2392];
    current_RowCol_1 = {img_addr, 10'd300};
  end
  else if (detected_keypoint[1][300]) begin
    filter_input_1_0 = buffer_data_5[2423:2400];
    filter_input_1_1 = buffer_data_4[2423:2400];
    filter_input_1_2 = blur5x5_1_dout[2423:2400];
    current_RowCol_1 = {img_addr, 10'd301};
  end
  else if (detected_keypoint[1][301]) begin
    filter_input_1_0 = buffer_data_5[2431:2408];
    filter_input_1_1 = buffer_data_4[2431:2408];
    filter_input_1_2 = blur5x5_1_dout[2431:2408];
    current_RowCol_1 = {img_addr, 10'd302};
  end
  else if (detected_keypoint[1][302]) begin
    filter_input_1_0 = buffer_data_5[2439:2416];
    filter_input_1_1 = buffer_data_4[2439:2416];
    filter_input_1_2 = blur5x5_1_dout[2439:2416];
    current_RowCol_1 = {img_addr, 10'd303};
  end
  else if (detected_keypoint[1][303]) begin
    filter_input_1_0 = buffer_data_5[2447:2424];
    filter_input_1_1 = buffer_data_4[2447:2424];
    filter_input_1_2 = blur5x5_1_dout[2447:2424];
    current_RowCol_1 = {img_addr, 10'd304};
  end
  else if (detected_keypoint[1][304]) begin
    filter_input_1_0 = buffer_data_5[2455:2432];
    filter_input_1_1 = buffer_data_4[2455:2432];
    filter_input_1_2 = blur5x5_1_dout[2455:2432];
    current_RowCol_1 = {img_addr, 10'd305};
  end
  else if (detected_keypoint[1][305]) begin
    filter_input_1_0 = buffer_data_5[2463:2440];
    filter_input_1_1 = buffer_data_4[2463:2440];
    filter_input_1_2 = blur5x5_1_dout[2463:2440];
    current_RowCol_1 = {img_addr, 10'd306};
  end
  else if (detected_keypoint[1][306]) begin
    filter_input_1_0 = buffer_data_5[2471:2448];
    filter_input_1_1 = buffer_data_4[2471:2448];
    filter_input_1_2 = blur5x5_1_dout[2471:2448];
    current_RowCol_1 = {img_addr, 10'd307};
  end
  else if (detected_keypoint[1][307]) begin
    filter_input_1_0 = buffer_data_5[2479:2456];
    filter_input_1_1 = buffer_data_4[2479:2456];
    filter_input_1_2 = blur5x5_1_dout[2479:2456];
    current_RowCol_1 = {img_addr, 10'd308};
  end
  else if (detected_keypoint[1][308]) begin
    filter_input_1_0 = buffer_data_5[2487:2464];
    filter_input_1_1 = buffer_data_4[2487:2464];
    filter_input_1_2 = blur5x5_1_dout[2487:2464];
    current_RowCol_1 = {img_addr, 10'd309};
  end
  else if (detected_keypoint[1][309]) begin
    filter_input_1_0 = buffer_data_5[2495:2472];
    filter_input_1_1 = buffer_data_4[2495:2472];
    filter_input_1_2 = blur5x5_1_dout[2495:2472];
    current_RowCol_1 = {img_addr, 10'd310};
  end
  else if (detected_keypoint[1][310]) begin
    filter_input_1_0 = buffer_data_5[2503:2480];
    filter_input_1_1 = buffer_data_4[2503:2480];
    filter_input_1_2 = blur5x5_1_dout[2503:2480];
    current_RowCol_1 = {img_addr, 10'd311};
  end
  else if (detected_keypoint[1][311]) begin
    filter_input_1_0 = buffer_data_5[2511:2488];
    filter_input_1_1 = buffer_data_4[2511:2488];
    filter_input_1_2 = blur5x5_1_dout[2511:2488];
    current_RowCol_1 = {img_addr, 10'd312};
  end
  else if (detected_keypoint[1][312]) begin
    filter_input_1_0 = buffer_data_5[2519:2496];
    filter_input_1_1 = buffer_data_4[2519:2496];
    filter_input_1_2 = blur5x5_1_dout[2519:2496];
    current_RowCol_1 = {img_addr, 10'd313};
  end
  else if (detected_keypoint[1][313]) begin
    filter_input_1_0 = buffer_data_5[2527:2504];
    filter_input_1_1 = buffer_data_4[2527:2504];
    filter_input_1_2 = blur5x5_1_dout[2527:2504];
    current_RowCol_1 = {img_addr, 10'd314};
  end
  else if (detected_keypoint[1][314]) begin
    filter_input_1_0 = buffer_data_5[2535:2512];
    filter_input_1_1 = buffer_data_4[2535:2512];
    filter_input_1_2 = blur5x5_1_dout[2535:2512];
    current_RowCol_1 = {img_addr, 10'd315};
  end
  else if (detected_keypoint[1][315]) begin
    filter_input_1_0 = buffer_data_5[2543:2520];
    filter_input_1_1 = buffer_data_4[2543:2520];
    filter_input_1_2 = blur5x5_1_dout[2543:2520];
    current_RowCol_1 = {img_addr, 10'd316};
  end
  else if (detected_keypoint[1][316]) begin
    filter_input_1_0 = buffer_data_5[2551:2528];
    filter_input_1_1 = buffer_data_4[2551:2528];
    filter_input_1_2 = blur5x5_1_dout[2551:2528];
    current_RowCol_1 = {img_addr, 10'd317};
  end
  else if (detected_keypoint[1][317]) begin
    filter_input_1_0 = buffer_data_5[2559:2536];
    filter_input_1_1 = buffer_data_4[2559:2536];
    filter_input_1_2 = blur5x5_1_dout[2559:2536];
    current_RowCol_1 = {img_addr, 10'd318};
  end
  else if (detected_keypoint[1][318]) begin
    filter_input_1_0 = buffer_data_5[2567:2544];
    filter_input_1_1 = buffer_data_4[2567:2544];
    filter_input_1_2 = blur5x5_1_dout[2567:2544];
    current_RowCol_1 = {img_addr, 10'd319};
  end
  else if (detected_keypoint[1][319]) begin
    filter_input_1_0 = buffer_data_5[2575:2552];
    filter_input_1_1 = buffer_data_4[2575:2552];
    filter_input_1_2 = blur5x5_1_dout[2575:2552];
    current_RowCol_1 = {img_addr, 10'd320};
  end
  else if (detected_keypoint[1][320]) begin
    filter_input_1_0 = buffer_data_5[2583:2560];
    filter_input_1_1 = buffer_data_4[2583:2560];
    filter_input_1_2 = blur5x5_1_dout[2583:2560];
    current_RowCol_1 = {img_addr, 10'd321};
  end
  else if (detected_keypoint[1][321]) begin
    filter_input_1_0 = buffer_data_5[2591:2568];
    filter_input_1_1 = buffer_data_4[2591:2568];
    filter_input_1_2 = blur5x5_1_dout[2591:2568];
    current_RowCol_1 = {img_addr, 10'd322};
  end
  else if (detected_keypoint[1][322]) begin
    filter_input_1_0 = buffer_data_5[2599:2576];
    filter_input_1_1 = buffer_data_4[2599:2576];
    filter_input_1_2 = blur5x5_1_dout[2599:2576];
    current_RowCol_1 = {img_addr, 10'd323};
  end
  else if (detected_keypoint[1][323]) begin
    filter_input_1_0 = buffer_data_5[2607:2584];
    filter_input_1_1 = buffer_data_4[2607:2584];
    filter_input_1_2 = blur5x5_1_dout[2607:2584];
    current_RowCol_1 = {img_addr, 10'd324};
  end
  else if (detected_keypoint[1][324]) begin
    filter_input_1_0 = buffer_data_5[2615:2592];
    filter_input_1_1 = buffer_data_4[2615:2592];
    filter_input_1_2 = blur5x5_1_dout[2615:2592];
    current_RowCol_1 = {img_addr, 10'd325};
  end
  else if (detected_keypoint[1][325]) begin
    filter_input_1_0 = buffer_data_5[2623:2600];
    filter_input_1_1 = buffer_data_4[2623:2600];
    filter_input_1_2 = blur5x5_1_dout[2623:2600];
    current_RowCol_1 = {img_addr, 10'd326};
  end
  else if (detected_keypoint[1][326]) begin
    filter_input_1_0 = buffer_data_5[2631:2608];
    filter_input_1_1 = buffer_data_4[2631:2608];
    filter_input_1_2 = blur5x5_1_dout[2631:2608];
    current_RowCol_1 = {img_addr, 10'd327};
  end
  else if (detected_keypoint[1][327]) begin
    filter_input_1_0 = buffer_data_5[2639:2616];
    filter_input_1_1 = buffer_data_4[2639:2616];
    filter_input_1_2 = blur5x5_1_dout[2639:2616];
    current_RowCol_1 = {img_addr, 10'd328};
  end
  else if (detected_keypoint[1][328]) begin
    filter_input_1_0 = buffer_data_5[2647:2624];
    filter_input_1_1 = buffer_data_4[2647:2624];
    filter_input_1_2 = blur5x5_1_dout[2647:2624];
    current_RowCol_1 = {img_addr, 10'd329};
  end
  else if (detected_keypoint[1][329]) begin
    filter_input_1_0 = buffer_data_5[2655:2632];
    filter_input_1_1 = buffer_data_4[2655:2632];
    filter_input_1_2 = blur5x5_1_dout[2655:2632];
    current_RowCol_1 = {img_addr, 10'd330};
  end
  else if (detected_keypoint[1][330]) begin
    filter_input_1_0 = buffer_data_5[2663:2640];
    filter_input_1_1 = buffer_data_4[2663:2640];
    filter_input_1_2 = blur5x5_1_dout[2663:2640];
    current_RowCol_1 = {img_addr, 10'd331};
  end
  else if (detected_keypoint[1][331]) begin
    filter_input_1_0 = buffer_data_5[2671:2648];
    filter_input_1_1 = buffer_data_4[2671:2648];
    filter_input_1_2 = blur5x5_1_dout[2671:2648];
    current_RowCol_1 = {img_addr, 10'd332};
  end
  else if (detected_keypoint[1][332]) begin
    filter_input_1_0 = buffer_data_5[2679:2656];
    filter_input_1_1 = buffer_data_4[2679:2656];
    filter_input_1_2 = blur5x5_1_dout[2679:2656];
    current_RowCol_1 = {img_addr, 10'd333};
  end
  else if (detected_keypoint[1][333]) begin
    filter_input_1_0 = buffer_data_5[2687:2664];
    filter_input_1_1 = buffer_data_4[2687:2664];
    filter_input_1_2 = blur5x5_1_dout[2687:2664];
    current_RowCol_1 = {img_addr, 10'd334};
  end
  else if (detected_keypoint[1][334]) begin
    filter_input_1_0 = buffer_data_5[2695:2672];
    filter_input_1_1 = buffer_data_4[2695:2672];
    filter_input_1_2 = blur5x5_1_dout[2695:2672];
    current_RowCol_1 = {img_addr, 10'd335};
  end
  else if (detected_keypoint[1][335]) begin
    filter_input_1_0 = buffer_data_5[2703:2680];
    filter_input_1_1 = buffer_data_4[2703:2680];
    filter_input_1_2 = blur5x5_1_dout[2703:2680];
    current_RowCol_1 = {img_addr, 10'd336};
  end
  else if (detected_keypoint[1][336]) begin
    filter_input_1_0 = buffer_data_5[2711:2688];
    filter_input_1_1 = buffer_data_4[2711:2688];
    filter_input_1_2 = blur5x5_1_dout[2711:2688];
    current_RowCol_1 = {img_addr, 10'd337};
  end
  else if (detected_keypoint[1][337]) begin
    filter_input_1_0 = buffer_data_5[2719:2696];
    filter_input_1_1 = buffer_data_4[2719:2696];
    filter_input_1_2 = blur5x5_1_dout[2719:2696];
    current_RowCol_1 = {img_addr, 10'd338};
  end
  else if (detected_keypoint[1][338]) begin
    filter_input_1_0 = buffer_data_5[2727:2704];
    filter_input_1_1 = buffer_data_4[2727:2704];
    filter_input_1_2 = blur5x5_1_dout[2727:2704];
    current_RowCol_1 = {img_addr, 10'd339};
  end
  else if (detected_keypoint[1][339]) begin
    filter_input_1_0 = buffer_data_5[2735:2712];
    filter_input_1_1 = buffer_data_4[2735:2712];
    filter_input_1_2 = blur5x5_1_dout[2735:2712];
    current_RowCol_1 = {img_addr, 10'd340};
  end
  else if (detected_keypoint[1][340]) begin
    filter_input_1_0 = buffer_data_5[2743:2720];
    filter_input_1_1 = buffer_data_4[2743:2720];
    filter_input_1_2 = blur5x5_1_dout[2743:2720];
    current_RowCol_1 = {img_addr, 10'd341};
  end
  else if (detected_keypoint[1][341]) begin
    filter_input_1_0 = buffer_data_5[2751:2728];
    filter_input_1_1 = buffer_data_4[2751:2728];
    filter_input_1_2 = blur5x5_1_dout[2751:2728];
    current_RowCol_1 = {img_addr, 10'd342};
  end
  else if (detected_keypoint[1][342]) begin
    filter_input_1_0 = buffer_data_5[2759:2736];
    filter_input_1_1 = buffer_data_4[2759:2736];
    filter_input_1_2 = blur5x5_1_dout[2759:2736];
    current_RowCol_1 = {img_addr, 10'd343};
  end
  else if (detected_keypoint[1][343]) begin
    filter_input_1_0 = buffer_data_5[2767:2744];
    filter_input_1_1 = buffer_data_4[2767:2744];
    filter_input_1_2 = blur5x5_1_dout[2767:2744];
    current_RowCol_1 = {img_addr, 10'd344};
  end
  else if (detected_keypoint[1][344]) begin
    filter_input_1_0 = buffer_data_5[2775:2752];
    filter_input_1_1 = buffer_data_4[2775:2752];
    filter_input_1_2 = blur5x5_1_dout[2775:2752];
    current_RowCol_1 = {img_addr, 10'd345};
  end
  else if (detected_keypoint[1][345]) begin
    filter_input_1_0 = buffer_data_5[2783:2760];
    filter_input_1_1 = buffer_data_4[2783:2760];
    filter_input_1_2 = blur5x5_1_dout[2783:2760];
    current_RowCol_1 = {img_addr, 10'd346};
  end
  else if (detected_keypoint[1][346]) begin
    filter_input_1_0 = buffer_data_5[2791:2768];
    filter_input_1_1 = buffer_data_4[2791:2768];
    filter_input_1_2 = blur5x5_1_dout[2791:2768];
    current_RowCol_1 = {img_addr, 10'd347};
  end
  else if (detected_keypoint[1][347]) begin
    filter_input_1_0 = buffer_data_5[2799:2776];
    filter_input_1_1 = buffer_data_4[2799:2776];
    filter_input_1_2 = blur5x5_1_dout[2799:2776];
    current_RowCol_1 = {img_addr, 10'd348};
  end
  else if (detected_keypoint[1][348]) begin
    filter_input_1_0 = buffer_data_5[2807:2784];
    filter_input_1_1 = buffer_data_4[2807:2784];
    filter_input_1_2 = blur5x5_1_dout[2807:2784];
    current_RowCol_1 = {img_addr, 10'd349};
  end
  else if (detected_keypoint[1][349]) begin
    filter_input_1_0 = buffer_data_5[2815:2792];
    filter_input_1_1 = buffer_data_4[2815:2792];
    filter_input_1_2 = blur5x5_1_dout[2815:2792];
    current_RowCol_1 = {img_addr, 10'd350};
  end
  else if (detected_keypoint[1][350]) begin
    filter_input_1_0 = buffer_data_5[2823:2800];
    filter_input_1_1 = buffer_data_4[2823:2800];
    filter_input_1_2 = blur5x5_1_dout[2823:2800];
    current_RowCol_1 = {img_addr, 10'd351};
  end
  else if (detected_keypoint[1][351]) begin
    filter_input_1_0 = buffer_data_5[2831:2808];
    filter_input_1_1 = buffer_data_4[2831:2808];
    filter_input_1_2 = blur5x5_1_dout[2831:2808];
    current_RowCol_1 = {img_addr, 10'd352};
  end
  else if (detected_keypoint[1][352]) begin
    filter_input_1_0 = buffer_data_5[2839:2816];
    filter_input_1_1 = buffer_data_4[2839:2816];
    filter_input_1_2 = blur5x5_1_dout[2839:2816];
    current_RowCol_1 = {img_addr, 10'd353};
  end
  else if (detected_keypoint[1][353]) begin
    filter_input_1_0 = buffer_data_5[2847:2824];
    filter_input_1_1 = buffer_data_4[2847:2824];
    filter_input_1_2 = blur5x5_1_dout[2847:2824];
    current_RowCol_1 = {img_addr, 10'd354};
  end
  else if (detected_keypoint[1][354]) begin
    filter_input_1_0 = buffer_data_5[2855:2832];
    filter_input_1_1 = buffer_data_4[2855:2832];
    filter_input_1_2 = blur5x5_1_dout[2855:2832];
    current_RowCol_1 = {img_addr, 10'd355};
  end
  else if (detected_keypoint[1][355]) begin
    filter_input_1_0 = buffer_data_5[2863:2840];
    filter_input_1_1 = buffer_data_4[2863:2840];
    filter_input_1_2 = blur5x5_1_dout[2863:2840];
    current_RowCol_1 = {img_addr, 10'd356};
  end
  else if (detected_keypoint[1][356]) begin
    filter_input_1_0 = buffer_data_5[2871:2848];
    filter_input_1_1 = buffer_data_4[2871:2848];
    filter_input_1_2 = blur5x5_1_dout[2871:2848];
    current_RowCol_1 = {img_addr, 10'd357};
  end
  else if (detected_keypoint[1][357]) begin
    filter_input_1_0 = buffer_data_5[2879:2856];
    filter_input_1_1 = buffer_data_4[2879:2856];
    filter_input_1_2 = blur5x5_1_dout[2879:2856];
    current_RowCol_1 = {img_addr, 10'd358};
  end
  else if (detected_keypoint[1][358]) begin
    filter_input_1_0 = buffer_data_5[2887:2864];
    filter_input_1_1 = buffer_data_4[2887:2864];
    filter_input_1_2 = blur5x5_1_dout[2887:2864];
    current_RowCol_1 = {img_addr, 10'd359};
  end
  else if (detected_keypoint[1][359]) begin
    filter_input_1_0 = buffer_data_5[2895:2872];
    filter_input_1_1 = buffer_data_4[2895:2872];
    filter_input_1_2 = blur5x5_1_dout[2895:2872];
    current_RowCol_1 = {img_addr, 10'd360};
  end
  else if (detected_keypoint[1][360]) begin
    filter_input_1_0 = buffer_data_5[2903:2880];
    filter_input_1_1 = buffer_data_4[2903:2880];
    filter_input_1_2 = blur5x5_1_dout[2903:2880];
    current_RowCol_1 = {img_addr, 10'd361};
  end
  else if (detected_keypoint[1][361]) begin
    filter_input_1_0 = buffer_data_5[2911:2888];
    filter_input_1_1 = buffer_data_4[2911:2888];
    filter_input_1_2 = blur5x5_1_dout[2911:2888];
    current_RowCol_1 = {img_addr, 10'd362};
  end
  else if (detected_keypoint[1][362]) begin
    filter_input_1_0 = buffer_data_5[2919:2896];
    filter_input_1_1 = buffer_data_4[2919:2896];
    filter_input_1_2 = blur5x5_1_dout[2919:2896];
    current_RowCol_1 = {img_addr, 10'd363};
  end
  else if (detected_keypoint[1][363]) begin
    filter_input_1_0 = buffer_data_5[2927:2904];
    filter_input_1_1 = buffer_data_4[2927:2904];
    filter_input_1_2 = blur5x5_1_dout[2927:2904];
    current_RowCol_1 = {img_addr, 10'd364};
  end
  else if (detected_keypoint[1][364]) begin
    filter_input_1_0 = buffer_data_5[2935:2912];
    filter_input_1_1 = buffer_data_4[2935:2912];
    filter_input_1_2 = blur5x5_1_dout[2935:2912];
    current_RowCol_1 = {img_addr, 10'd365};
  end
  else if (detected_keypoint[1][365]) begin
    filter_input_1_0 = buffer_data_5[2943:2920];
    filter_input_1_1 = buffer_data_4[2943:2920];
    filter_input_1_2 = blur5x5_1_dout[2943:2920];
    current_RowCol_1 = {img_addr, 10'd366};
  end
  else if (detected_keypoint[1][366]) begin
    filter_input_1_0 = buffer_data_5[2951:2928];
    filter_input_1_1 = buffer_data_4[2951:2928];
    filter_input_1_2 = blur5x5_1_dout[2951:2928];
    current_RowCol_1 = {img_addr, 10'd367};
  end
  else if (detected_keypoint[1][367]) begin
    filter_input_1_0 = buffer_data_5[2959:2936];
    filter_input_1_1 = buffer_data_4[2959:2936];
    filter_input_1_2 = blur5x5_1_dout[2959:2936];
    current_RowCol_1 = {img_addr, 10'd368};
  end
  else if (detected_keypoint[1][368]) begin
    filter_input_1_0 = buffer_data_5[2967:2944];
    filter_input_1_1 = buffer_data_4[2967:2944];
    filter_input_1_2 = blur5x5_1_dout[2967:2944];
    current_RowCol_1 = {img_addr, 10'd369};
  end
  else if (detected_keypoint[1][369]) begin
    filter_input_1_0 = buffer_data_5[2975:2952];
    filter_input_1_1 = buffer_data_4[2975:2952];
    filter_input_1_2 = blur5x5_1_dout[2975:2952];
    current_RowCol_1 = {img_addr, 10'd370};
  end
  else if (detected_keypoint[1][370]) begin
    filter_input_1_0 = buffer_data_5[2983:2960];
    filter_input_1_1 = buffer_data_4[2983:2960];
    filter_input_1_2 = blur5x5_1_dout[2983:2960];
    current_RowCol_1 = {img_addr, 10'd371};
  end
  else if (detected_keypoint[1][371]) begin
    filter_input_1_0 = buffer_data_5[2991:2968];
    filter_input_1_1 = buffer_data_4[2991:2968];
    filter_input_1_2 = blur5x5_1_dout[2991:2968];
    current_RowCol_1 = {img_addr, 10'd372};
  end
  else if (detected_keypoint[1][372]) begin
    filter_input_1_0 = buffer_data_5[2999:2976];
    filter_input_1_1 = buffer_data_4[2999:2976];
    filter_input_1_2 = blur5x5_1_dout[2999:2976];
    current_RowCol_1 = {img_addr, 10'd373};
  end
  else if (detected_keypoint[1][373]) begin
    filter_input_1_0 = buffer_data_5[3007:2984];
    filter_input_1_1 = buffer_data_4[3007:2984];
    filter_input_1_2 = blur5x5_1_dout[3007:2984];
    current_RowCol_1 = {img_addr, 10'd374};
  end
  else if (detected_keypoint[1][374]) begin
    filter_input_1_0 = buffer_data_5[3015:2992];
    filter_input_1_1 = buffer_data_4[3015:2992];
    filter_input_1_2 = blur5x5_1_dout[3015:2992];
    current_RowCol_1 = {img_addr, 10'd375};
  end
  else if (detected_keypoint[1][375]) begin
    filter_input_1_0 = buffer_data_5[3023:3000];
    filter_input_1_1 = buffer_data_4[3023:3000];
    filter_input_1_2 = blur5x5_1_dout[3023:3000];
    current_RowCol_1 = {img_addr, 10'd376};
  end
  else if (detected_keypoint[1][376]) begin
    filter_input_1_0 = buffer_data_5[3031:3008];
    filter_input_1_1 = buffer_data_4[3031:3008];
    filter_input_1_2 = blur5x5_1_dout[3031:3008];
    current_RowCol_1 = {img_addr, 10'd377};
  end
  else if (detected_keypoint[1][377]) begin
    filter_input_1_0 = buffer_data_5[3039:3016];
    filter_input_1_1 = buffer_data_4[3039:3016];
    filter_input_1_2 = blur5x5_1_dout[3039:3016];
    current_RowCol_1 = {img_addr, 10'd378};
  end
  else if (detected_keypoint[1][378]) begin
    filter_input_1_0 = buffer_data_5[3047:3024];
    filter_input_1_1 = buffer_data_4[3047:3024];
    filter_input_1_2 = blur5x5_1_dout[3047:3024];
    current_RowCol_1 = {img_addr, 10'd379};
  end
  else if (detected_keypoint[1][379]) begin
    filter_input_1_0 = buffer_data_5[3055:3032];
    filter_input_1_1 = buffer_data_4[3055:3032];
    filter_input_1_2 = blur5x5_1_dout[3055:3032];
    current_RowCol_1 = {img_addr, 10'd380};
  end
  else if (detected_keypoint[1][380]) begin
    filter_input_1_0 = buffer_data_5[3063:3040];
    filter_input_1_1 = buffer_data_4[3063:3040];
    filter_input_1_2 = blur5x5_1_dout[3063:3040];
    current_RowCol_1 = {img_addr, 10'd381};
  end
  else if (detected_keypoint[1][381]) begin
    filter_input_1_0 = buffer_data_5[3071:3048];
    filter_input_1_1 = buffer_data_4[3071:3048];
    filter_input_1_2 = blur5x5_1_dout[3071:3048];
    current_RowCol_1 = {img_addr, 10'd382};
  end
  else if (detected_keypoint[1][382]) begin
    filter_input_1_0 = buffer_data_5[3079:3056];
    filter_input_1_1 = buffer_data_4[3079:3056];
    filter_input_1_2 = blur5x5_1_dout[3079:3056];
    current_RowCol_1 = {img_addr, 10'd383};
  end
  else if (detected_keypoint[1][383]) begin
    filter_input_1_0 = buffer_data_5[3087:3064];
    filter_input_1_1 = buffer_data_4[3087:3064];
    filter_input_1_2 = blur5x5_1_dout[3087:3064];
    current_RowCol_1 = {img_addr, 10'd384};
  end
  else if (detected_keypoint[1][384]) begin
    filter_input_1_0 = buffer_data_5[3095:3072];
    filter_input_1_1 = buffer_data_4[3095:3072];
    filter_input_1_2 = blur5x5_1_dout[3095:3072];
    current_RowCol_1 = {img_addr, 10'd385};
  end
  else if (detected_keypoint[1][385]) begin
    filter_input_1_0 = buffer_data_5[3103:3080];
    filter_input_1_1 = buffer_data_4[3103:3080];
    filter_input_1_2 = blur5x5_1_dout[3103:3080];
    current_RowCol_1 = {img_addr, 10'd386};
  end
  else if (detected_keypoint[1][386]) begin
    filter_input_1_0 = buffer_data_5[3111:3088];
    filter_input_1_1 = buffer_data_4[3111:3088];
    filter_input_1_2 = blur5x5_1_dout[3111:3088];
    current_RowCol_1 = {img_addr, 10'd387};
  end
  else if (detected_keypoint[1][387]) begin
    filter_input_1_0 = buffer_data_5[3119:3096];
    filter_input_1_1 = buffer_data_4[3119:3096];
    filter_input_1_2 = blur5x5_1_dout[3119:3096];
    current_RowCol_1 = {img_addr, 10'd388};
  end
  else if (detected_keypoint[1][388]) begin
    filter_input_1_0 = buffer_data_5[3127:3104];
    filter_input_1_1 = buffer_data_4[3127:3104];
    filter_input_1_2 = blur5x5_1_dout[3127:3104];
    current_RowCol_1 = {img_addr, 10'd389};
  end
  else if (detected_keypoint[1][389]) begin
    filter_input_1_0 = buffer_data_5[3135:3112];
    filter_input_1_1 = buffer_data_4[3135:3112];
    filter_input_1_2 = blur5x5_1_dout[3135:3112];
    current_RowCol_1 = {img_addr, 10'd390};
  end
  else if (detected_keypoint[1][390]) begin
    filter_input_1_0 = buffer_data_5[3143:3120];
    filter_input_1_1 = buffer_data_4[3143:3120];
    filter_input_1_2 = blur5x5_1_dout[3143:3120];
    current_RowCol_1 = {img_addr, 10'd391};
  end
  else if (detected_keypoint[1][391]) begin
    filter_input_1_0 = buffer_data_5[3151:3128];
    filter_input_1_1 = buffer_data_4[3151:3128];
    filter_input_1_2 = blur5x5_1_dout[3151:3128];
    current_RowCol_1 = {img_addr, 10'd392};
  end
  else if (detected_keypoint[1][392]) begin
    filter_input_1_0 = buffer_data_5[3159:3136];
    filter_input_1_1 = buffer_data_4[3159:3136];
    filter_input_1_2 = blur5x5_1_dout[3159:3136];
    current_RowCol_1 = {img_addr, 10'd393};
  end
  else if (detected_keypoint[1][393]) begin
    filter_input_1_0 = buffer_data_5[3167:3144];
    filter_input_1_1 = buffer_data_4[3167:3144];
    filter_input_1_2 = blur5x5_1_dout[3167:3144];
    current_RowCol_1 = {img_addr, 10'd394};
  end
  else if (detected_keypoint[1][394]) begin
    filter_input_1_0 = buffer_data_5[3175:3152];
    filter_input_1_1 = buffer_data_4[3175:3152];
    filter_input_1_2 = blur5x5_1_dout[3175:3152];
    current_RowCol_1 = {img_addr, 10'd395};
  end
  else if (detected_keypoint[1][395]) begin
    filter_input_1_0 = buffer_data_5[3183:3160];
    filter_input_1_1 = buffer_data_4[3183:3160];
    filter_input_1_2 = blur5x5_1_dout[3183:3160];
    current_RowCol_1 = {img_addr, 10'd396};
  end
  else if (detected_keypoint[1][396]) begin
    filter_input_1_0 = buffer_data_5[3191:3168];
    filter_input_1_1 = buffer_data_4[3191:3168];
    filter_input_1_2 = blur5x5_1_dout[3191:3168];
    current_RowCol_1 = {img_addr, 10'd397};
  end
  else if (detected_keypoint[1][397]) begin
    filter_input_1_0 = buffer_data_5[3199:3176];
    filter_input_1_1 = buffer_data_4[3199:3176];
    filter_input_1_2 = blur5x5_1_dout[3199:3176];
    current_RowCol_1 = {img_addr, 10'd398};
  end
  else if (detected_keypoint[1][398]) begin
    filter_input_1_0 = buffer_data_5[3207:3184];
    filter_input_1_1 = buffer_data_4[3207:3184];
    filter_input_1_2 = blur5x5_1_dout[3207:3184];
    current_RowCol_1 = {img_addr, 10'd399};
  end
  else if (detected_keypoint[1][399]) begin
    filter_input_1_0 = buffer_data_5[3215:3192];
    filter_input_1_1 = buffer_data_4[3215:3192];
    filter_input_1_2 = blur5x5_1_dout[3215:3192];
    current_RowCol_1 = {img_addr, 10'd400};
  end
  else if (detected_keypoint[1][400]) begin
    filter_input_1_0 = buffer_data_5[3223:3200];
    filter_input_1_1 = buffer_data_4[3223:3200];
    filter_input_1_2 = blur5x5_1_dout[3223:3200];
    current_RowCol_1 = {img_addr, 10'd401};
  end
  else if (detected_keypoint[1][401]) begin
    filter_input_1_0 = buffer_data_5[3231:3208];
    filter_input_1_1 = buffer_data_4[3231:3208];
    filter_input_1_2 = blur5x5_1_dout[3231:3208];
    current_RowCol_1 = {img_addr, 10'd402};
  end
  else if (detected_keypoint[1][402]) begin
    filter_input_1_0 = buffer_data_5[3239:3216];
    filter_input_1_1 = buffer_data_4[3239:3216];
    filter_input_1_2 = blur5x5_1_dout[3239:3216];
    current_RowCol_1 = {img_addr, 10'd403};
  end
  else if (detected_keypoint[1][403]) begin
    filter_input_1_0 = buffer_data_5[3247:3224];
    filter_input_1_1 = buffer_data_4[3247:3224];
    filter_input_1_2 = blur5x5_1_dout[3247:3224];
    current_RowCol_1 = {img_addr, 10'd404};
  end
  else if (detected_keypoint[1][404]) begin
    filter_input_1_0 = buffer_data_5[3255:3232];
    filter_input_1_1 = buffer_data_4[3255:3232];
    filter_input_1_2 = blur5x5_1_dout[3255:3232];
    current_RowCol_1 = {img_addr, 10'd405};
  end
  else if (detected_keypoint[1][405]) begin
    filter_input_1_0 = buffer_data_5[3263:3240];
    filter_input_1_1 = buffer_data_4[3263:3240];
    filter_input_1_2 = blur5x5_1_dout[3263:3240];
    current_RowCol_1 = {img_addr, 10'd406};
  end
  else if (detected_keypoint[1][406]) begin
    filter_input_1_0 = buffer_data_5[3271:3248];
    filter_input_1_1 = buffer_data_4[3271:3248];
    filter_input_1_2 = blur5x5_1_dout[3271:3248];
    current_RowCol_1 = {img_addr, 10'd407};
  end
  else if (detected_keypoint[1][407]) begin
    filter_input_1_0 = buffer_data_5[3279:3256];
    filter_input_1_1 = buffer_data_4[3279:3256];
    filter_input_1_2 = blur5x5_1_dout[3279:3256];
    current_RowCol_1 = {img_addr, 10'd408};
  end
  else if (detected_keypoint[1][408]) begin
    filter_input_1_0 = buffer_data_5[3287:3264];
    filter_input_1_1 = buffer_data_4[3287:3264];
    filter_input_1_2 = blur5x5_1_dout[3287:3264];
    current_RowCol_1 = {img_addr, 10'd409};
  end
  else if (detected_keypoint[1][409]) begin
    filter_input_1_0 = buffer_data_5[3295:3272];
    filter_input_1_1 = buffer_data_4[3295:3272];
    filter_input_1_2 = blur5x5_1_dout[3295:3272];
    current_RowCol_1 = {img_addr, 10'd410};
  end
  else if (detected_keypoint[1][410]) begin
    filter_input_1_0 = buffer_data_5[3303:3280];
    filter_input_1_1 = buffer_data_4[3303:3280];
    filter_input_1_2 = blur5x5_1_dout[3303:3280];
    current_RowCol_1 = {img_addr, 10'd411};
  end
  else if (detected_keypoint[1][411]) begin
    filter_input_1_0 = buffer_data_5[3311:3288];
    filter_input_1_1 = buffer_data_4[3311:3288];
    filter_input_1_2 = blur5x5_1_dout[3311:3288];
    current_RowCol_1 = {img_addr, 10'd412};
  end
  else if (detected_keypoint[1][412]) begin
    filter_input_1_0 = buffer_data_5[3319:3296];
    filter_input_1_1 = buffer_data_4[3319:3296];
    filter_input_1_2 = blur5x5_1_dout[3319:3296];
    current_RowCol_1 = {img_addr, 10'd413};
  end
  else if (detected_keypoint[1][413]) begin
    filter_input_1_0 = buffer_data_5[3327:3304];
    filter_input_1_1 = buffer_data_4[3327:3304];
    filter_input_1_2 = blur5x5_1_dout[3327:3304];
    current_RowCol_1 = {img_addr, 10'd414};
  end
  else if (detected_keypoint[1][414]) begin
    filter_input_1_0 = buffer_data_5[3335:3312];
    filter_input_1_1 = buffer_data_4[3335:3312];
    filter_input_1_2 = blur5x5_1_dout[3335:3312];
    current_RowCol_1 = {img_addr, 10'd415};
  end
  else if (detected_keypoint[1][415]) begin
    filter_input_1_0 = buffer_data_5[3343:3320];
    filter_input_1_1 = buffer_data_4[3343:3320];
    filter_input_1_2 = blur5x5_1_dout[3343:3320];
    current_RowCol_1 = {img_addr, 10'd416};
  end
  else if (detected_keypoint[1][416]) begin
    filter_input_1_0 = buffer_data_5[3351:3328];
    filter_input_1_1 = buffer_data_4[3351:3328];
    filter_input_1_2 = blur5x5_1_dout[3351:3328];
    current_RowCol_1 = {img_addr, 10'd417};
  end
  else if (detected_keypoint[1][417]) begin
    filter_input_1_0 = buffer_data_5[3359:3336];
    filter_input_1_1 = buffer_data_4[3359:3336];
    filter_input_1_2 = blur5x5_1_dout[3359:3336];
    current_RowCol_1 = {img_addr, 10'd418};
  end
  else if (detected_keypoint[1][418]) begin
    filter_input_1_0 = buffer_data_5[3367:3344];
    filter_input_1_1 = buffer_data_4[3367:3344];
    filter_input_1_2 = blur5x5_1_dout[3367:3344];
    current_RowCol_1 = {img_addr, 10'd419};
  end
  else if (detected_keypoint[1][419]) begin
    filter_input_1_0 = buffer_data_5[3375:3352];
    filter_input_1_1 = buffer_data_4[3375:3352];
    filter_input_1_2 = blur5x5_1_dout[3375:3352];
    current_RowCol_1 = {img_addr, 10'd420};
  end
  else if (detected_keypoint[1][420]) begin
    filter_input_1_0 = buffer_data_5[3383:3360];
    filter_input_1_1 = buffer_data_4[3383:3360];
    filter_input_1_2 = blur5x5_1_dout[3383:3360];
    current_RowCol_1 = {img_addr, 10'd421};
  end
  else if (detected_keypoint[1][421]) begin
    filter_input_1_0 = buffer_data_5[3391:3368];
    filter_input_1_1 = buffer_data_4[3391:3368];
    filter_input_1_2 = blur5x5_1_dout[3391:3368];
    current_RowCol_1 = {img_addr, 10'd422};
  end
  else if (detected_keypoint[1][422]) begin
    filter_input_1_0 = buffer_data_5[3399:3376];
    filter_input_1_1 = buffer_data_4[3399:3376];
    filter_input_1_2 = blur5x5_1_dout[3399:3376];
    current_RowCol_1 = {img_addr, 10'd423};
  end
  else if (detected_keypoint[1][423]) begin
    filter_input_1_0 = buffer_data_5[3407:3384];
    filter_input_1_1 = buffer_data_4[3407:3384];
    filter_input_1_2 = blur5x5_1_dout[3407:3384];
    current_RowCol_1 = {img_addr, 10'd424};
  end
  else if (detected_keypoint[1][424]) begin
    filter_input_1_0 = buffer_data_5[3415:3392];
    filter_input_1_1 = buffer_data_4[3415:3392];
    filter_input_1_2 = blur5x5_1_dout[3415:3392];
    current_RowCol_1 = {img_addr, 10'd425};
  end
  else if (detected_keypoint[1][425]) begin
    filter_input_1_0 = buffer_data_5[3423:3400];
    filter_input_1_1 = buffer_data_4[3423:3400];
    filter_input_1_2 = blur5x5_1_dout[3423:3400];
    current_RowCol_1 = {img_addr, 10'd426};
  end
  else if (detected_keypoint[1][426]) begin
    filter_input_1_0 = buffer_data_5[3431:3408];
    filter_input_1_1 = buffer_data_4[3431:3408];
    filter_input_1_2 = blur5x5_1_dout[3431:3408];
    current_RowCol_1 = {img_addr, 10'd427};
  end
  else if (detected_keypoint[1][427]) begin
    filter_input_1_0 = buffer_data_5[3439:3416];
    filter_input_1_1 = buffer_data_4[3439:3416];
    filter_input_1_2 = blur5x5_1_dout[3439:3416];
    current_RowCol_1 = {img_addr, 10'd428};
  end
  else if (detected_keypoint[1][428]) begin
    filter_input_1_0 = buffer_data_5[3447:3424];
    filter_input_1_1 = buffer_data_4[3447:3424];
    filter_input_1_2 = blur5x5_1_dout[3447:3424];
    current_RowCol_1 = {img_addr, 10'd429};
  end
  else if (detected_keypoint[1][429]) begin
    filter_input_1_0 = buffer_data_5[3455:3432];
    filter_input_1_1 = buffer_data_4[3455:3432];
    filter_input_1_2 = blur5x5_1_dout[3455:3432];
    current_RowCol_1 = {img_addr, 10'd430};
  end
  else if (detected_keypoint[1][430]) begin
    filter_input_1_0 = buffer_data_5[3463:3440];
    filter_input_1_1 = buffer_data_4[3463:3440];
    filter_input_1_2 = blur5x5_1_dout[3463:3440];
    current_RowCol_1 = {img_addr, 10'd431};
  end
  else if (detected_keypoint[1][431]) begin
    filter_input_1_0 = buffer_data_5[3471:3448];
    filter_input_1_1 = buffer_data_4[3471:3448];
    filter_input_1_2 = blur5x5_1_dout[3471:3448];
    current_RowCol_1 = {img_addr, 10'd432};
  end
  else if (detected_keypoint[1][432]) begin
    filter_input_1_0 = buffer_data_5[3479:3456];
    filter_input_1_1 = buffer_data_4[3479:3456];
    filter_input_1_2 = blur5x5_1_dout[3479:3456];
    current_RowCol_1 = {img_addr, 10'd433};
  end
  else if (detected_keypoint[1][433]) begin
    filter_input_1_0 = buffer_data_5[3487:3464];
    filter_input_1_1 = buffer_data_4[3487:3464];
    filter_input_1_2 = blur5x5_1_dout[3487:3464];
    current_RowCol_1 = {img_addr, 10'd434};
  end
  else if (detected_keypoint[1][434]) begin
    filter_input_1_0 = buffer_data_5[3495:3472];
    filter_input_1_1 = buffer_data_4[3495:3472];
    filter_input_1_2 = blur5x5_1_dout[3495:3472];
    current_RowCol_1 = {img_addr, 10'd435};
  end
  else if (detected_keypoint[1][435]) begin
    filter_input_1_0 = buffer_data_5[3503:3480];
    filter_input_1_1 = buffer_data_4[3503:3480];
    filter_input_1_2 = blur5x5_1_dout[3503:3480];
    current_RowCol_1 = {img_addr, 10'd436};
  end
  else if (detected_keypoint[1][436]) begin
    filter_input_1_0 = buffer_data_5[3511:3488];
    filter_input_1_1 = buffer_data_4[3511:3488];
    filter_input_1_2 = blur5x5_1_dout[3511:3488];
    current_RowCol_1 = {img_addr, 10'd437};
  end
  else if (detected_keypoint[1][437]) begin
    filter_input_1_0 = buffer_data_5[3519:3496];
    filter_input_1_1 = buffer_data_4[3519:3496];
    filter_input_1_2 = blur5x5_1_dout[3519:3496];
    current_RowCol_1 = {img_addr, 10'd438};
  end
  else if (detected_keypoint[1][438]) begin
    filter_input_1_0 = buffer_data_5[3527:3504];
    filter_input_1_1 = buffer_data_4[3527:3504];
    filter_input_1_2 = blur5x5_1_dout[3527:3504];
    current_RowCol_1 = {img_addr, 10'd439};
  end
  else if (detected_keypoint[1][439]) begin
    filter_input_1_0 = buffer_data_5[3535:3512];
    filter_input_1_1 = buffer_data_4[3535:3512];
    filter_input_1_2 = blur5x5_1_dout[3535:3512];
    current_RowCol_1 = {img_addr, 10'd440};
  end
  else if (detected_keypoint[1][440]) begin
    filter_input_1_0 = buffer_data_5[3543:3520];
    filter_input_1_1 = buffer_data_4[3543:3520];
    filter_input_1_2 = blur5x5_1_dout[3543:3520];
    current_RowCol_1 = {img_addr, 10'd441};
  end
  else if (detected_keypoint[1][441]) begin
    filter_input_1_0 = buffer_data_5[3551:3528];
    filter_input_1_1 = buffer_data_4[3551:3528];
    filter_input_1_2 = blur5x5_1_dout[3551:3528];
    current_RowCol_1 = {img_addr, 10'd442};
  end
  else if (detected_keypoint[1][442]) begin
    filter_input_1_0 = buffer_data_5[3559:3536];
    filter_input_1_1 = buffer_data_4[3559:3536];
    filter_input_1_2 = blur5x5_1_dout[3559:3536];
    current_RowCol_1 = {img_addr, 10'd443};
  end
  else if (detected_keypoint[1][443]) begin
    filter_input_1_0 = buffer_data_5[3567:3544];
    filter_input_1_1 = buffer_data_4[3567:3544];
    filter_input_1_2 = blur5x5_1_dout[3567:3544];
    current_RowCol_1 = {img_addr, 10'd444};
  end
  else if (detected_keypoint[1][444]) begin
    filter_input_1_0 = buffer_data_5[3575:3552];
    filter_input_1_1 = buffer_data_4[3575:3552];
    filter_input_1_2 = blur5x5_1_dout[3575:3552];
    current_RowCol_1 = {img_addr, 10'd445};
  end
  else if (detected_keypoint[1][445]) begin
    filter_input_1_0 = buffer_data_5[3583:3560];
    filter_input_1_1 = buffer_data_4[3583:3560];
    filter_input_1_2 = blur5x5_1_dout[3583:3560];
    current_RowCol_1 = {img_addr, 10'd446};
  end
  else if (detected_keypoint[1][446]) begin
    filter_input_1_0 = buffer_data_5[3591:3568];
    filter_input_1_1 = buffer_data_4[3591:3568];
    filter_input_1_2 = blur5x5_1_dout[3591:3568];
    current_RowCol_1 = {img_addr, 10'd447};
  end
  else if (detected_keypoint[1][447]) begin
    filter_input_1_0 = buffer_data_5[3599:3576];
    filter_input_1_1 = buffer_data_4[3599:3576];
    filter_input_1_2 = blur5x5_1_dout[3599:3576];
    current_RowCol_1 = {img_addr, 10'd448};
  end
  else if (detected_keypoint[1][448]) begin
    filter_input_1_0 = buffer_data_5[3607:3584];
    filter_input_1_1 = buffer_data_4[3607:3584];
    filter_input_1_2 = blur5x5_1_dout[3607:3584];
    current_RowCol_1 = {img_addr, 10'd449};
  end
  else if (detected_keypoint[1][449]) begin
    filter_input_1_0 = buffer_data_5[3615:3592];
    filter_input_1_1 = buffer_data_4[3615:3592];
    filter_input_1_2 = blur5x5_1_dout[3615:3592];
    current_RowCol_1 = {img_addr, 10'd450};
  end
  else if (detected_keypoint[1][450]) begin
    filter_input_1_0 = buffer_data_5[3623:3600];
    filter_input_1_1 = buffer_data_4[3623:3600];
    filter_input_1_2 = blur5x5_1_dout[3623:3600];
    current_RowCol_1 = {img_addr, 10'd451};
  end
  else if (detected_keypoint[1][451]) begin
    filter_input_1_0 = buffer_data_5[3631:3608];
    filter_input_1_1 = buffer_data_4[3631:3608];
    filter_input_1_2 = blur5x5_1_dout[3631:3608];
    current_RowCol_1 = {img_addr, 10'd452};
  end
  else if (detected_keypoint[1][452]) begin
    filter_input_1_0 = buffer_data_5[3639:3616];
    filter_input_1_1 = buffer_data_4[3639:3616];
    filter_input_1_2 = blur5x5_1_dout[3639:3616];
    current_RowCol_1 = {img_addr, 10'd453};
  end
  else if (detected_keypoint[1][453]) begin
    filter_input_1_0 = buffer_data_5[3647:3624];
    filter_input_1_1 = buffer_data_4[3647:3624];
    filter_input_1_2 = blur5x5_1_dout[3647:3624];
    current_RowCol_1 = {img_addr, 10'd454};
  end
  else if (detected_keypoint[1][454]) begin
    filter_input_1_0 = buffer_data_5[3655:3632];
    filter_input_1_1 = buffer_data_4[3655:3632];
    filter_input_1_2 = blur5x5_1_dout[3655:3632];
    current_RowCol_1 = {img_addr, 10'd455};
  end
  else if (detected_keypoint[1][455]) begin
    filter_input_1_0 = buffer_data_5[3663:3640];
    filter_input_1_1 = buffer_data_4[3663:3640];
    filter_input_1_2 = blur5x5_1_dout[3663:3640];
    current_RowCol_1 = {img_addr, 10'd456};
  end
  else if (detected_keypoint[1][456]) begin
    filter_input_1_0 = buffer_data_5[3671:3648];
    filter_input_1_1 = buffer_data_4[3671:3648];
    filter_input_1_2 = blur5x5_1_dout[3671:3648];
    current_RowCol_1 = {img_addr, 10'd457};
  end
  else if (detected_keypoint[1][457]) begin
    filter_input_1_0 = buffer_data_5[3679:3656];
    filter_input_1_1 = buffer_data_4[3679:3656];
    filter_input_1_2 = blur5x5_1_dout[3679:3656];
    current_RowCol_1 = {img_addr, 10'd458};
  end
  else if (detected_keypoint[1][458]) begin
    filter_input_1_0 = buffer_data_5[3687:3664];
    filter_input_1_1 = buffer_data_4[3687:3664];
    filter_input_1_2 = blur5x5_1_dout[3687:3664];
    current_RowCol_1 = {img_addr, 10'd459};
  end
  else if (detected_keypoint[1][459]) begin
    filter_input_1_0 = buffer_data_5[3695:3672];
    filter_input_1_1 = buffer_data_4[3695:3672];
    filter_input_1_2 = blur5x5_1_dout[3695:3672];
    current_RowCol_1 = {img_addr, 10'd460};
  end
  else if (detected_keypoint[1][460]) begin
    filter_input_1_0 = buffer_data_5[3703:3680];
    filter_input_1_1 = buffer_data_4[3703:3680];
    filter_input_1_2 = blur5x5_1_dout[3703:3680];
    current_RowCol_1 = {img_addr, 10'd461};
  end
  else if (detected_keypoint[1][461]) begin
    filter_input_1_0 = buffer_data_5[3711:3688];
    filter_input_1_1 = buffer_data_4[3711:3688];
    filter_input_1_2 = blur5x5_1_dout[3711:3688];
    current_RowCol_1 = {img_addr, 10'd462};
  end
  else if (detected_keypoint[1][462]) begin
    filter_input_1_0 = buffer_data_5[3719:3696];
    filter_input_1_1 = buffer_data_4[3719:3696];
    filter_input_1_2 = blur5x5_1_dout[3719:3696];
    current_RowCol_1 = {img_addr, 10'd463};
  end
  else if (detected_keypoint[1][463]) begin
    filter_input_1_0 = buffer_data_5[3727:3704];
    filter_input_1_1 = buffer_data_4[3727:3704];
    filter_input_1_2 = blur5x5_1_dout[3727:3704];
    current_RowCol_1 = {img_addr, 10'd464};
  end
  else if (detected_keypoint[1][464]) begin
    filter_input_1_0 = buffer_data_5[3735:3712];
    filter_input_1_1 = buffer_data_4[3735:3712];
    filter_input_1_2 = blur5x5_1_dout[3735:3712];
    current_RowCol_1 = {img_addr, 10'd465};
  end
  else if (detected_keypoint[1][465]) begin
    filter_input_1_0 = buffer_data_5[3743:3720];
    filter_input_1_1 = buffer_data_4[3743:3720];
    filter_input_1_2 = blur5x5_1_dout[3743:3720];
    current_RowCol_1 = {img_addr, 10'd466};
  end
  else if (detected_keypoint[1][466]) begin
    filter_input_1_0 = buffer_data_5[3751:3728];
    filter_input_1_1 = buffer_data_4[3751:3728];
    filter_input_1_2 = blur5x5_1_dout[3751:3728];
    current_RowCol_1 = {img_addr, 10'd467};
  end
  else if (detected_keypoint[1][467]) begin
    filter_input_1_0 = buffer_data_5[3759:3736];
    filter_input_1_1 = buffer_data_4[3759:3736];
    filter_input_1_2 = blur5x5_1_dout[3759:3736];
    current_RowCol_1 = {img_addr, 10'd468};
  end
  else if (detected_keypoint[1][468]) begin
    filter_input_1_0 = buffer_data_5[3767:3744];
    filter_input_1_1 = buffer_data_4[3767:3744];
    filter_input_1_2 = blur5x5_1_dout[3767:3744];
    current_RowCol_1 = {img_addr, 10'd469};
  end
  else if (detected_keypoint[1][469]) begin
    filter_input_1_0 = buffer_data_5[3775:3752];
    filter_input_1_1 = buffer_data_4[3775:3752];
    filter_input_1_2 = blur5x5_1_dout[3775:3752];
    current_RowCol_1 = {img_addr, 10'd470};
  end
  else if (detected_keypoint[1][470]) begin
    filter_input_1_0 = buffer_data_5[3783:3760];
    filter_input_1_1 = buffer_data_4[3783:3760];
    filter_input_1_2 = blur5x5_1_dout[3783:3760];
    current_RowCol_1 = {img_addr, 10'd471};
  end
  else if (detected_keypoint[1][471]) begin
    filter_input_1_0 = buffer_data_5[3791:3768];
    filter_input_1_1 = buffer_data_4[3791:3768];
    filter_input_1_2 = blur5x5_1_dout[3791:3768];
    current_RowCol_1 = {img_addr, 10'd472};
  end
  else if (detected_keypoint[1][472]) begin
    filter_input_1_0 = buffer_data_5[3799:3776];
    filter_input_1_1 = buffer_data_4[3799:3776];
    filter_input_1_2 = blur5x5_1_dout[3799:3776];
    current_RowCol_1 = {img_addr, 10'd473};
  end
  else if (detected_keypoint[1][473]) begin
    filter_input_1_0 = buffer_data_5[3807:3784];
    filter_input_1_1 = buffer_data_4[3807:3784];
    filter_input_1_2 = blur5x5_1_dout[3807:3784];
    current_RowCol_1 = {img_addr, 10'd474};
  end
  else if (detected_keypoint[1][474]) begin
    filter_input_1_0 = buffer_data_5[3815:3792];
    filter_input_1_1 = buffer_data_4[3815:3792];
    filter_input_1_2 = blur5x5_1_dout[3815:3792];
    current_RowCol_1 = {img_addr, 10'd475};
  end
  else if (detected_keypoint[1][475]) begin
    filter_input_1_0 = buffer_data_5[3823:3800];
    filter_input_1_1 = buffer_data_4[3823:3800];
    filter_input_1_2 = blur5x5_1_dout[3823:3800];
    current_RowCol_1 = {img_addr, 10'd476};
  end
  else if (detected_keypoint[1][476]) begin
    filter_input_1_0 = buffer_data_5[3831:3808];
    filter_input_1_1 = buffer_data_4[3831:3808];
    filter_input_1_2 = blur5x5_1_dout[3831:3808];
    current_RowCol_1 = {img_addr, 10'd477};
  end
  else if (detected_keypoint[1][477]) begin
    filter_input_1_0 = buffer_data_5[3839:3816];
    filter_input_1_1 = buffer_data_4[3839:3816];
    filter_input_1_2 = blur5x5_1_dout[3839:3816];
    current_RowCol_1 = {img_addr, 10'd478};
  end
  else if (detected_keypoint[1][478]) begin
    filter_input_1_0 = buffer_data_5[3847:3824];
    filter_input_1_1 = buffer_data_4[3847:3824];
    filter_input_1_2 = blur5x5_1_dout[3847:3824];
    current_RowCol_1 = {img_addr, 10'd479};
  end
  else if (detected_keypoint[1][479]) begin
    filter_input_1_0 = buffer_data_5[3855:3832];
    filter_input_1_1 = buffer_data_4[3855:3832];
    filter_input_1_2 = blur5x5_1_dout[3855:3832];
    current_RowCol_1 = {img_addr, 10'd480};
  end
  else if (detected_keypoint[1][480]) begin
    filter_input_1_0 = buffer_data_5[3863:3840];
    filter_input_1_1 = buffer_data_4[3863:3840];
    filter_input_1_2 = blur5x5_1_dout[3863:3840];
    current_RowCol_1 = {img_addr, 10'd481};
  end
  else if (detected_keypoint[1][481]) begin
    filter_input_1_0 = buffer_data_5[3871:3848];
    filter_input_1_1 = buffer_data_4[3871:3848];
    filter_input_1_2 = blur5x5_1_dout[3871:3848];
    current_RowCol_1 = {img_addr, 10'd482};
  end
  else if (detected_keypoint[1][482]) begin
    filter_input_1_0 = buffer_data_5[3879:3856];
    filter_input_1_1 = buffer_data_4[3879:3856];
    filter_input_1_2 = blur5x5_1_dout[3879:3856];
    current_RowCol_1 = {img_addr, 10'd483};
  end
  else if (detected_keypoint[1][483]) begin
    filter_input_1_0 = buffer_data_5[3887:3864];
    filter_input_1_1 = buffer_data_4[3887:3864];
    filter_input_1_2 = blur5x5_1_dout[3887:3864];
    current_RowCol_1 = {img_addr, 10'd484};
  end
  else if (detected_keypoint[1][484]) begin
    filter_input_1_0 = buffer_data_5[3895:3872];
    filter_input_1_1 = buffer_data_4[3895:3872];
    filter_input_1_2 = blur5x5_1_dout[3895:3872];
    current_RowCol_1 = {img_addr, 10'd485};
  end
  else if (detected_keypoint[1][485]) begin
    filter_input_1_0 = buffer_data_5[3903:3880];
    filter_input_1_1 = buffer_data_4[3903:3880];
    filter_input_1_2 = blur5x5_1_dout[3903:3880];
    current_RowCol_1 = {img_addr, 10'd486};
  end
  else if (detected_keypoint[1][486]) begin
    filter_input_1_0 = buffer_data_5[3911:3888];
    filter_input_1_1 = buffer_data_4[3911:3888];
    filter_input_1_2 = blur5x5_1_dout[3911:3888];
    current_RowCol_1 = {img_addr, 10'd487};
  end
  else if (detected_keypoint[1][487]) begin
    filter_input_1_0 = buffer_data_5[3919:3896];
    filter_input_1_1 = buffer_data_4[3919:3896];
    filter_input_1_2 = blur5x5_1_dout[3919:3896];
    current_RowCol_1 = {img_addr, 10'd488};
  end
  else if (detected_keypoint[1][488]) begin
    filter_input_1_0 = buffer_data_5[3927:3904];
    filter_input_1_1 = buffer_data_4[3927:3904];
    filter_input_1_2 = blur5x5_1_dout[3927:3904];
    current_RowCol_1 = {img_addr, 10'd489};
  end
  else if (detected_keypoint[1][489]) begin
    filter_input_1_0 = buffer_data_5[3935:3912];
    filter_input_1_1 = buffer_data_4[3935:3912];
    filter_input_1_2 = blur5x5_1_dout[3935:3912];
    current_RowCol_1 = {img_addr, 10'd490};
  end
  else if (detected_keypoint[1][490]) begin
    filter_input_1_0 = buffer_data_5[3943:3920];
    filter_input_1_1 = buffer_data_4[3943:3920];
    filter_input_1_2 = blur5x5_1_dout[3943:3920];
    current_RowCol_1 = {img_addr, 10'd491};
  end
  else if (detected_keypoint[1][491]) begin
    filter_input_1_0 = buffer_data_5[3951:3928];
    filter_input_1_1 = buffer_data_4[3951:3928];
    filter_input_1_2 = blur5x5_1_dout[3951:3928];
    current_RowCol_1 = {img_addr, 10'd492};
  end
  else if (detected_keypoint[1][492]) begin
    filter_input_1_0 = buffer_data_5[3959:3936];
    filter_input_1_1 = buffer_data_4[3959:3936];
    filter_input_1_2 = blur5x5_1_dout[3959:3936];
    current_RowCol_1 = {img_addr, 10'd493};
  end
  else if (detected_keypoint[1][493]) begin
    filter_input_1_0 = buffer_data_5[3967:3944];
    filter_input_1_1 = buffer_data_4[3967:3944];
    filter_input_1_2 = blur5x5_1_dout[3967:3944];
    current_RowCol_1 = {img_addr, 10'd494};
  end
  else if (detected_keypoint[1][494]) begin
    filter_input_1_0 = buffer_data_5[3975:3952];
    filter_input_1_1 = buffer_data_4[3975:3952];
    filter_input_1_2 = blur5x5_1_dout[3975:3952];
    current_RowCol_1 = {img_addr, 10'd495};
  end
  else if (detected_keypoint[1][495]) begin
    filter_input_1_0 = buffer_data_5[3983:3960];
    filter_input_1_1 = buffer_data_4[3983:3960];
    filter_input_1_2 = blur5x5_1_dout[3983:3960];
    current_RowCol_1 = {img_addr, 10'd496};
  end
  else if (detected_keypoint[1][496]) begin
    filter_input_1_0 = buffer_data_5[3991:3968];
    filter_input_1_1 = buffer_data_4[3991:3968];
    filter_input_1_2 = blur5x5_1_dout[3991:3968];
    current_RowCol_1 = {img_addr, 10'd497};
  end
  else if (detected_keypoint[1][497]) begin
    filter_input_1_0 = buffer_data_5[3999:3976];
    filter_input_1_1 = buffer_data_4[3999:3976];
    filter_input_1_2 = blur5x5_1_dout[3999:3976];
    current_RowCol_1 = {img_addr, 10'd498};
  end
  else if (detected_keypoint[1][498]) begin
    filter_input_1_0 = buffer_data_5[4007:3984];
    filter_input_1_1 = buffer_data_4[4007:3984];
    filter_input_1_2 = blur5x5_1_dout[4007:3984];
    current_RowCol_1 = {img_addr, 10'd499};
  end
  else if (detected_keypoint[1][499]) begin
    filter_input_1_0 = buffer_data_5[4015:3992];
    filter_input_1_1 = buffer_data_4[4015:3992];
    filter_input_1_2 = blur5x5_1_dout[4015:3992];
    current_RowCol_1 = {img_addr, 10'd500};
  end
  else if (detected_keypoint[1][500]) begin
    filter_input_1_0 = buffer_data_5[4023:4000];
    filter_input_1_1 = buffer_data_4[4023:4000];
    filter_input_1_2 = blur5x5_1_dout[4023:4000];
    current_RowCol_1 = {img_addr, 10'd501};
  end
  else if (detected_keypoint[1][501]) begin
    filter_input_1_0 = buffer_data_5[4031:4008];
    filter_input_1_1 = buffer_data_4[4031:4008];
    filter_input_1_2 = blur5x5_1_dout[4031:4008];
    current_RowCol_1 = {img_addr, 10'd502};
  end
  else if (detected_keypoint[1][502]) begin
    filter_input_1_0 = buffer_data_5[4039:4016];
    filter_input_1_1 = buffer_data_4[4039:4016];
    filter_input_1_2 = blur5x5_1_dout[4039:4016];
    current_RowCol_1 = {img_addr, 10'd503};
  end
  else if (detected_keypoint[1][503]) begin
    filter_input_1_0 = buffer_data_5[4047:4024];
    filter_input_1_1 = buffer_data_4[4047:4024];
    filter_input_1_2 = blur5x5_1_dout[4047:4024];
    current_RowCol_1 = {img_addr, 10'd504};
  end
  else if (detected_keypoint[1][504]) begin
    filter_input_1_0 = buffer_data_5[4055:4032];
    filter_input_1_1 = buffer_data_4[4055:4032];
    filter_input_1_2 = blur5x5_1_dout[4055:4032];
    current_RowCol_1 = {img_addr, 10'd505};
  end
  else if (detected_keypoint[1][505]) begin
    filter_input_1_0 = buffer_data_5[4063:4040];
    filter_input_1_1 = buffer_data_4[4063:4040];
    filter_input_1_2 = blur5x5_1_dout[4063:4040];
    current_RowCol_1 = {img_addr, 10'd506};
  end
  else if (detected_keypoint[1][506]) begin
    filter_input_1_0 = buffer_data_5[4071:4048];
    filter_input_1_1 = buffer_data_4[4071:4048];
    filter_input_1_2 = blur5x5_1_dout[4071:4048];
    current_RowCol_1 = {img_addr, 10'd507};
  end
  else if (detected_keypoint[1][507]) begin
    filter_input_1_0 = buffer_data_5[4079:4056];
    filter_input_1_1 = buffer_data_4[4079:4056];
    filter_input_1_2 = blur5x5_1_dout[4079:4056];
    current_RowCol_1 = {img_addr, 10'd508};
  end
  else if (detected_keypoint[1][508]) begin
    filter_input_1_0 = buffer_data_5[4087:4064];
    filter_input_1_1 = buffer_data_4[4087:4064];
    filter_input_1_2 = blur5x5_1_dout[4087:4064];
    current_RowCol_1 = {img_addr, 10'd509};
  end
  else if (detected_keypoint[1][509]) begin
    filter_input_1_0 = buffer_data_5[4095:4072];
    filter_input_1_1 = buffer_data_4[4095:4072];
    filter_input_1_2 = blur5x5_1_dout[4095:4072];
    current_RowCol_1 = {img_addr, 10'd510};
  end
  else if (detected_keypoint[1][510]) begin
    filter_input_1_0 = buffer_data_5[4103:4080];
    filter_input_1_1 = buffer_data_4[4103:4080];
    filter_input_1_2 = blur5x5_1_dout[4103:4080];
    current_RowCol_1 = {img_addr, 10'd511};
  end
  else if (detected_keypoint[1][511]) begin
    filter_input_1_0 = buffer_data_5[4111:4088];
    filter_input_1_1 = buffer_data_4[4111:4088];
    filter_input_1_2 = blur5x5_1_dout[4111:4088];
    current_RowCol_1 = {img_addr, 10'd512};
  end
  else if (detected_keypoint[1][512]) begin
    filter_input_1_0 = buffer_data_5[4119:4096];
    filter_input_1_1 = buffer_data_4[4119:4096];
    filter_input_1_2 = blur5x5_1_dout[4119:4096];
    current_RowCol_1 = {img_addr, 10'd513};
  end
  else if (detected_keypoint[1][513]) begin
    filter_input_1_0 = buffer_data_5[4127:4104];
    filter_input_1_1 = buffer_data_4[4127:4104];
    filter_input_1_2 = blur5x5_1_dout[4127:4104];
    current_RowCol_1 = {img_addr, 10'd514};
  end
  else if (detected_keypoint[1][514]) begin
    filter_input_1_0 = buffer_data_5[4135:4112];
    filter_input_1_1 = buffer_data_4[4135:4112];
    filter_input_1_2 = blur5x5_1_dout[4135:4112];
    current_RowCol_1 = {img_addr, 10'd515};
  end
  else if (detected_keypoint[1][515]) begin
    filter_input_1_0 = buffer_data_5[4143:4120];
    filter_input_1_1 = buffer_data_4[4143:4120];
    filter_input_1_2 = blur5x5_1_dout[4143:4120];
    current_RowCol_1 = {img_addr, 10'd516};
  end
  else if (detected_keypoint[1][516]) begin
    filter_input_1_0 = buffer_data_5[4151:4128];
    filter_input_1_1 = buffer_data_4[4151:4128];
    filter_input_1_2 = blur5x5_1_dout[4151:4128];
    current_RowCol_1 = {img_addr, 10'd517};
  end
  else if (detected_keypoint[1][517]) begin
    filter_input_1_0 = buffer_data_5[4159:4136];
    filter_input_1_1 = buffer_data_4[4159:4136];
    filter_input_1_2 = blur5x5_1_dout[4159:4136];
    current_RowCol_1 = {img_addr, 10'd518};
  end
  else if (detected_keypoint[1][518]) begin
    filter_input_1_0 = buffer_data_5[4167:4144];
    filter_input_1_1 = buffer_data_4[4167:4144];
    filter_input_1_2 = blur5x5_1_dout[4167:4144];
    current_RowCol_1 = {img_addr, 10'd519};
  end
  else if (detected_keypoint[1][519]) begin
    filter_input_1_0 = buffer_data_5[4175:4152];
    filter_input_1_1 = buffer_data_4[4175:4152];
    filter_input_1_2 = blur5x5_1_dout[4175:4152];
    current_RowCol_1 = {img_addr, 10'd520};
  end
  else if (detected_keypoint[1][520]) begin
    filter_input_1_0 = buffer_data_5[4183:4160];
    filter_input_1_1 = buffer_data_4[4183:4160];
    filter_input_1_2 = blur5x5_1_dout[4183:4160];
    current_RowCol_1 = {img_addr, 10'd521};
  end
  else if (detected_keypoint[1][521]) begin
    filter_input_1_0 = buffer_data_5[4191:4168];
    filter_input_1_1 = buffer_data_4[4191:4168];
    filter_input_1_2 = blur5x5_1_dout[4191:4168];
    current_RowCol_1 = {img_addr, 10'd522};
  end
  else if (detected_keypoint[1][522]) begin
    filter_input_1_0 = buffer_data_5[4199:4176];
    filter_input_1_1 = buffer_data_4[4199:4176];
    filter_input_1_2 = blur5x5_1_dout[4199:4176];
    current_RowCol_1 = {img_addr, 10'd523};
  end
  else if (detected_keypoint[1][523]) begin
    filter_input_1_0 = buffer_data_5[4207:4184];
    filter_input_1_1 = buffer_data_4[4207:4184];
    filter_input_1_2 = blur5x5_1_dout[4207:4184];
    current_RowCol_1 = {img_addr, 10'd524};
  end
  else if (detected_keypoint[1][524]) begin
    filter_input_1_0 = buffer_data_5[4215:4192];
    filter_input_1_1 = buffer_data_4[4215:4192];
    filter_input_1_2 = blur5x5_1_dout[4215:4192];
    current_RowCol_1 = {img_addr, 10'd525};
  end
  else if (detected_keypoint[1][525]) begin
    filter_input_1_0 = buffer_data_5[4223:4200];
    filter_input_1_1 = buffer_data_4[4223:4200];
    filter_input_1_2 = blur5x5_1_dout[4223:4200];
    current_RowCol_1 = {img_addr, 10'd526};
  end
  else if (detected_keypoint[1][526]) begin
    filter_input_1_0 = buffer_data_5[4231:4208];
    filter_input_1_1 = buffer_data_4[4231:4208];
    filter_input_1_2 = blur5x5_1_dout[4231:4208];
    current_RowCol_1 = {img_addr, 10'd527};
  end
  else if (detected_keypoint[1][527]) begin
    filter_input_1_0 = buffer_data_5[4239:4216];
    filter_input_1_1 = buffer_data_4[4239:4216];
    filter_input_1_2 = blur5x5_1_dout[4239:4216];
    current_RowCol_1 = {img_addr, 10'd528};
  end
  else if (detected_keypoint[1][528]) begin
    filter_input_1_0 = buffer_data_5[4247:4224];
    filter_input_1_1 = buffer_data_4[4247:4224];
    filter_input_1_2 = blur5x5_1_dout[4247:4224];
    current_RowCol_1 = {img_addr, 10'd529};
  end
  else if (detected_keypoint[1][529]) begin
    filter_input_1_0 = buffer_data_5[4255:4232];
    filter_input_1_1 = buffer_data_4[4255:4232];
    filter_input_1_2 = blur5x5_1_dout[4255:4232];
    current_RowCol_1 = {img_addr, 10'd530};
  end
  else if (detected_keypoint[1][530]) begin
    filter_input_1_0 = buffer_data_5[4263:4240];
    filter_input_1_1 = buffer_data_4[4263:4240];
    filter_input_1_2 = blur5x5_1_dout[4263:4240];
    current_RowCol_1 = {img_addr, 10'd531};
  end
  else if (detected_keypoint[1][531]) begin
    filter_input_1_0 = buffer_data_5[4271:4248];
    filter_input_1_1 = buffer_data_4[4271:4248];
    filter_input_1_2 = blur5x5_1_dout[4271:4248];
    current_RowCol_1 = {img_addr, 10'd532};
  end
  else if (detected_keypoint[1][532]) begin
    filter_input_1_0 = buffer_data_5[4279:4256];
    filter_input_1_1 = buffer_data_4[4279:4256];
    filter_input_1_2 = blur5x5_1_dout[4279:4256];
    current_RowCol_1 = {img_addr, 10'd533};
  end
  else if (detected_keypoint[1][533]) begin
    filter_input_1_0 = buffer_data_5[4287:4264];
    filter_input_1_1 = buffer_data_4[4287:4264];
    filter_input_1_2 = blur5x5_1_dout[4287:4264];
    current_RowCol_1 = {img_addr, 10'd534};
  end
  else if (detected_keypoint[1][534]) begin
    filter_input_1_0 = buffer_data_5[4295:4272];
    filter_input_1_1 = buffer_data_4[4295:4272];
    filter_input_1_2 = blur5x5_1_dout[4295:4272];
    current_RowCol_1 = {img_addr, 10'd535};
  end
  else if (detected_keypoint[1][535]) begin
    filter_input_1_0 = buffer_data_5[4303:4280];
    filter_input_1_1 = buffer_data_4[4303:4280];
    filter_input_1_2 = blur5x5_1_dout[4303:4280];
    current_RowCol_1 = {img_addr, 10'd536};
  end
  else if (detected_keypoint[1][536]) begin
    filter_input_1_0 = buffer_data_5[4311:4288];
    filter_input_1_1 = buffer_data_4[4311:4288];
    filter_input_1_2 = blur5x5_1_dout[4311:4288];
    current_RowCol_1 = {img_addr, 10'd537};
  end
  else if (detected_keypoint[1][537]) begin
    filter_input_1_0 = buffer_data_5[4319:4296];
    filter_input_1_1 = buffer_data_4[4319:4296];
    filter_input_1_2 = blur5x5_1_dout[4319:4296];
    current_RowCol_1 = {img_addr, 10'd538};
  end
  else if (detected_keypoint[1][538]) begin
    filter_input_1_0 = buffer_data_5[4327:4304];
    filter_input_1_1 = buffer_data_4[4327:4304];
    filter_input_1_2 = blur5x5_1_dout[4327:4304];
    current_RowCol_1 = {img_addr, 10'd539};
  end
  else if (detected_keypoint[1][539]) begin
    filter_input_1_0 = buffer_data_5[4335:4312];
    filter_input_1_1 = buffer_data_4[4335:4312];
    filter_input_1_2 = blur5x5_1_dout[4335:4312];
    current_RowCol_1 = {img_addr, 10'd540};
  end
  else if (detected_keypoint[1][540]) begin
    filter_input_1_0 = buffer_data_5[4343:4320];
    filter_input_1_1 = buffer_data_4[4343:4320];
    filter_input_1_2 = blur5x5_1_dout[4343:4320];
    current_RowCol_1 = {img_addr, 10'd541};
  end
  else if (detected_keypoint[1][541]) begin
    filter_input_1_0 = buffer_data_5[4351:4328];
    filter_input_1_1 = buffer_data_4[4351:4328];
    filter_input_1_2 = blur5x5_1_dout[4351:4328];
    current_RowCol_1 = {img_addr, 10'd542};
  end
  else if (detected_keypoint[1][542]) begin
    filter_input_1_0 = buffer_data_5[4359:4336];
    filter_input_1_1 = buffer_data_4[4359:4336];
    filter_input_1_2 = blur5x5_1_dout[4359:4336];
    current_RowCol_1 = {img_addr, 10'd543};
  end
  else if (detected_keypoint[1][543]) begin
    filter_input_1_0 = buffer_data_5[4367:4344];
    filter_input_1_1 = buffer_data_4[4367:4344];
    filter_input_1_2 = blur5x5_1_dout[4367:4344];
    current_RowCol_1 = {img_addr, 10'd544};
  end
  else if (detected_keypoint[1][544]) begin
    filter_input_1_0 = buffer_data_5[4375:4352];
    filter_input_1_1 = buffer_data_4[4375:4352];
    filter_input_1_2 = blur5x5_1_dout[4375:4352];
    current_RowCol_1 = {img_addr, 10'd545};
  end
  else if (detected_keypoint[1][545]) begin
    filter_input_1_0 = buffer_data_5[4383:4360];
    filter_input_1_1 = buffer_data_4[4383:4360];
    filter_input_1_2 = blur5x5_1_dout[4383:4360];
    current_RowCol_1 = {img_addr, 10'd546};
  end
  else if (detected_keypoint[1][546]) begin
    filter_input_1_0 = buffer_data_5[4391:4368];
    filter_input_1_1 = buffer_data_4[4391:4368];
    filter_input_1_2 = blur5x5_1_dout[4391:4368];
    current_RowCol_1 = {img_addr, 10'd547};
  end
  else if (detected_keypoint[1][547]) begin
    filter_input_1_0 = buffer_data_5[4399:4376];
    filter_input_1_1 = buffer_data_4[4399:4376];
    filter_input_1_2 = blur5x5_1_dout[4399:4376];
    current_RowCol_1 = {img_addr, 10'd548};
  end
  else if (detected_keypoint[1][548]) begin
    filter_input_1_0 = buffer_data_5[4407:4384];
    filter_input_1_1 = buffer_data_4[4407:4384];
    filter_input_1_2 = blur5x5_1_dout[4407:4384];
    current_RowCol_1 = {img_addr, 10'd549};
  end
  else if (detected_keypoint[1][549]) begin
    filter_input_1_0 = buffer_data_5[4415:4392];
    filter_input_1_1 = buffer_data_4[4415:4392];
    filter_input_1_2 = blur5x5_1_dout[4415:4392];
    current_RowCol_1 = {img_addr, 10'd550};
  end
  else if (detected_keypoint[1][550]) begin
    filter_input_1_0 = buffer_data_5[4423:4400];
    filter_input_1_1 = buffer_data_4[4423:4400];
    filter_input_1_2 = blur5x5_1_dout[4423:4400];
    current_RowCol_1 = {img_addr, 10'd551};
  end
  else if (detected_keypoint[1][551]) begin
    filter_input_1_0 = buffer_data_5[4431:4408];
    filter_input_1_1 = buffer_data_4[4431:4408];
    filter_input_1_2 = blur5x5_1_dout[4431:4408];
    current_RowCol_1 = {img_addr, 10'd552};
  end
  else if (detected_keypoint[1][552]) begin
    filter_input_1_0 = buffer_data_5[4439:4416];
    filter_input_1_1 = buffer_data_4[4439:4416];
    filter_input_1_2 = blur5x5_1_dout[4439:4416];
    current_RowCol_1 = {img_addr, 10'd553};
  end
  else if (detected_keypoint[1][553]) begin
    filter_input_1_0 = buffer_data_5[4447:4424];
    filter_input_1_1 = buffer_data_4[4447:4424];
    filter_input_1_2 = blur5x5_1_dout[4447:4424];
    current_RowCol_1 = {img_addr, 10'd554};
  end
  else if (detected_keypoint[1][554]) begin
    filter_input_1_0 = buffer_data_5[4455:4432];
    filter_input_1_1 = buffer_data_4[4455:4432];
    filter_input_1_2 = blur5x5_1_dout[4455:4432];
    current_RowCol_1 = {img_addr, 10'd555};
  end
  else if (detected_keypoint[1][555]) begin
    filter_input_1_0 = buffer_data_5[4463:4440];
    filter_input_1_1 = buffer_data_4[4463:4440];
    filter_input_1_2 = blur5x5_1_dout[4463:4440];
    current_RowCol_1 = {img_addr, 10'd556};
  end
  else if (detected_keypoint[1][556]) begin
    filter_input_1_0 = buffer_data_5[4471:4448];
    filter_input_1_1 = buffer_data_4[4471:4448];
    filter_input_1_2 = blur5x5_1_dout[4471:4448];
    current_RowCol_1 = {img_addr, 10'd557};
  end
  else if (detected_keypoint[1][557]) begin
    filter_input_1_0 = buffer_data_5[4479:4456];
    filter_input_1_1 = buffer_data_4[4479:4456];
    filter_input_1_2 = blur5x5_1_dout[4479:4456];
    current_RowCol_1 = {img_addr, 10'd558};
  end
  else if (detected_keypoint[1][558]) begin
    filter_input_1_0 = buffer_data_5[4487:4464];
    filter_input_1_1 = buffer_data_4[4487:4464];
    filter_input_1_2 = blur5x5_1_dout[4487:4464];
    current_RowCol_1 = {img_addr, 10'd559};
  end
  else if (detected_keypoint[1][559]) begin
    filter_input_1_0 = buffer_data_5[4495:4472];
    filter_input_1_1 = buffer_data_4[4495:4472];
    filter_input_1_2 = blur5x5_1_dout[4495:4472];
    current_RowCol_1 = {img_addr, 10'd560};
  end
  else if (detected_keypoint[1][560]) begin
    filter_input_1_0 = buffer_data_5[4503:4480];
    filter_input_1_1 = buffer_data_4[4503:4480];
    filter_input_1_2 = blur5x5_1_dout[4503:4480];
    current_RowCol_1 = {img_addr, 10'd561};
  end
  else if (detected_keypoint[1][561]) begin
    filter_input_1_0 = buffer_data_5[4511:4488];
    filter_input_1_1 = buffer_data_4[4511:4488];
    filter_input_1_2 = blur5x5_1_dout[4511:4488];
    current_RowCol_1 = {img_addr, 10'd562};
  end
  else if (detected_keypoint[1][562]) begin
    filter_input_1_0 = buffer_data_5[4519:4496];
    filter_input_1_1 = buffer_data_4[4519:4496];
    filter_input_1_2 = blur5x5_1_dout[4519:4496];
    current_RowCol_1 = {img_addr, 10'd563};
  end
  else if (detected_keypoint[1][563]) begin
    filter_input_1_0 = buffer_data_5[4527:4504];
    filter_input_1_1 = buffer_data_4[4527:4504];
    filter_input_1_2 = blur5x5_1_dout[4527:4504];
    current_RowCol_1 = {img_addr, 10'd564};
  end
  else if (detected_keypoint[1][564]) begin
    filter_input_1_0 = buffer_data_5[4535:4512];
    filter_input_1_1 = buffer_data_4[4535:4512];
    filter_input_1_2 = blur5x5_1_dout[4535:4512];
    current_RowCol_1 = {img_addr, 10'd565};
  end
  else if (detected_keypoint[1][565]) begin
    filter_input_1_0 = buffer_data_5[4543:4520];
    filter_input_1_1 = buffer_data_4[4543:4520];
    filter_input_1_2 = blur5x5_1_dout[4543:4520];
    current_RowCol_1 = {img_addr, 10'd566};
  end
  else if (detected_keypoint[1][566]) begin
    filter_input_1_0 = buffer_data_5[4551:4528];
    filter_input_1_1 = buffer_data_4[4551:4528];
    filter_input_1_2 = blur5x5_1_dout[4551:4528];
    current_RowCol_1 = {img_addr, 10'd567};
  end
  else if (detected_keypoint[1][567]) begin
    filter_input_1_0 = buffer_data_5[4559:4536];
    filter_input_1_1 = buffer_data_4[4559:4536];
    filter_input_1_2 = blur5x5_1_dout[4559:4536];
    current_RowCol_1 = {img_addr, 10'd568};
  end
  else if (detected_keypoint[1][568]) begin
    filter_input_1_0 = buffer_data_5[4567:4544];
    filter_input_1_1 = buffer_data_4[4567:4544];
    filter_input_1_2 = blur5x5_1_dout[4567:4544];
    current_RowCol_1 = {img_addr, 10'd569};
  end
  else if (detected_keypoint[1][569]) begin
    filter_input_1_0 = buffer_data_5[4575:4552];
    filter_input_1_1 = buffer_data_4[4575:4552];
    filter_input_1_2 = blur5x5_1_dout[4575:4552];
    current_RowCol_1 = {img_addr, 10'd570};
  end
  else if (detected_keypoint[1][570]) begin
    filter_input_1_0 = buffer_data_5[4583:4560];
    filter_input_1_1 = buffer_data_4[4583:4560];
    filter_input_1_2 = blur5x5_1_dout[4583:4560];
    current_RowCol_1 = {img_addr, 10'd571};
  end
  else if (detected_keypoint[1][571]) begin
    filter_input_1_0 = buffer_data_5[4591:4568];
    filter_input_1_1 = buffer_data_4[4591:4568];
    filter_input_1_2 = blur5x5_1_dout[4591:4568];
    current_RowCol_1 = {img_addr, 10'd572};
  end
  else if (detected_keypoint[1][572]) begin
    filter_input_1_0 = buffer_data_5[4599:4576];
    filter_input_1_1 = buffer_data_4[4599:4576];
    filter_input_1_2 = blur5x5_1_dout[4599:4576];
    current_RowCol_1 = {img_addr, 10'd573};
  end
  else if (detected_keypoint[1][573]) begin
    filter_input_1_0 = buffer_data_5[4607:4584];
    filter_input_1_1 = buffer_data_4[4607:4584];
    filter_input_1_2 = blur5x5_1_dout[4607:4584];
    current_RowCol_1 = {img_addr, 10'd574};
  end
  else if (detected_keypoint[1][574]) begin
    filter_input_1_0 = buffer_data_5[4615:4592];
    filter_input_1_1 = buffer_data_4[4615:4592];
    filter_input_1_2 = blur5x5_1_dout[4615:4592];
    current_RowCol_1 = {img_addr, 10'd575};
  end
  else if (detected_keypoint[1][575]) begin
    filter_input_1_0 = buffer_data_5[4623:4600];
    filter_input_1_1 = buffer_data_4[4623:4600];
    filter_input_1_2 = blur5x5_1_dout[4623:4600];
    current_RowCol_1 = {img_addr, 10'd576};
  end
  else if (detected_keypoint[1][576]) begin
    filter_input_1_0 = buffer_data_5[4631:4608];
    filter_input_1_1 = buffer_data_4[4631:4608];
    filter_input_1_2 = blur5x5_1_dout[4631:4608];
    current_RowCol_1 = {img_addr, 10'd577};
  end
  else if (detected_keypoint[1][577]) begin
    filter_input_1_0 = buffer_data_5[4639:4616];
    filter_input_1_1 = buffer_data_4[4639:4616];
    filter_input_1_2 = blur5x5_1_dout[4639:4616];
    current_RowCol_1 = {img_addr, 10'd578};
  end
  else if (detected_keypoint[1][578]) begin
    filter_input_1_0 = buffer_data_5[4647:4624];
    filter_input_1_1 = buffer_data_4[4647:4624];
    filter_input_1_2 = blur5x5_1_dout[4647:4624];
    current_RowCol_1 = {img_addr, 10'd579};
  end
  else if (detected_keypoint[1][579]) begin
    filter_input_1_0 = buffer_data_5[4655:4632];
    filter_input_1_1 = buffer_data_4[4655:4632];
    filter_input_1_2 = blur5x5_1_dout[4655:4632];
    current_RowCol_1 = {img_addr, 10'd580};
  end
  else if (detected_keypoint[1][580]) begin
    filter_input_1_0 = buffer_data_5[4663:4640];
    filter_input_1_1 = buffer_data_4[4663:4640];
    filter_input_1_2 = blur5x5_1_dout[4663:4640];
    current_RowCol_1 = {img_addr, 10'd581};
  end
  else if (detected_keypoint[1][581]) begin
    filter_input_1_0 = buffer_data_5[4671:4648];
    filter_input_1_1 = buffer_data_4[4671:4648];
    filter_input_1_2 = blur5x5_1_dout[4671:4648];
    current_RowCol_1 = {img_addr, 10'd582};
  end
  else if (detected_keypoint[1][582]) begin
    filter_input_1_0 = buffer_data_5[4679:4656];
    filter_input_1_1 = buffer_data_4[4679:4656];
    filter_input_1_2 = blur5x5_1_dout[4679:4656];
    current_RowCol_1 = {img_addr, 10'd583};
  end
  else if (detected_keypoint[1][583]) begin
    filter_input_1_0 = buffer_data_5[4687:4664];
    filter_input_1_1 = buffer_data_4[4687:4664];
    filter_input_1_2 = blur5x5_1_dout[4687:4664];
    current_RowCol_1 = {img_addr, 10'd584};
  end
  else if (detected_keypoint[1][584]) begin
    filter_input_1_0 = buffer_data_5[4695:4672];
    filter_input_1_1 = buffer_data_4[4695:4672];
    filter_input_1_2 = blur5x5_1_dout[4695:4672];
    current_RowCol_1 = {img_addr, 10'd585};
  end
  else if (detected_keypoint[1][585]) begin
    filter_input_1_0 = buffer_data_5[4703:4680];
    filter_input_1_1 = buffer_data_4[4703:4680];
    filter_input_1_2 = blur5x5_1_dout[4703:4680];
    current_RowCol_1 = {img_addr, 10'd586};
  end
  else if (detected_keypoint[1][586]) begin
    filter_input_1_0 = buffer_data_5[4711:4688];
    filter_input_1_1 = buffer_data_4[4711:4688];
    filter_input_1_2 = blur5x5_1_dout[4711:4688];
    current_RowCol_1 = {img_addr, 10'd587};
  end
  else if (detected_keypoint[1][587]) begin
    filter_input_1_0 = buffer_data_5[4719:4696];
    filter_input_1_1 = buffer_data_4[4719:4696];
    filter_input_1_2 = blur5x5_1_dout[4719:4696];
    current_RowCol_1 = {img_addr, 10'd588};
  end
  else if (detected_keypoint[1][588]) begin
    filter_input_1_0 = buffer_data_5[4727:4704];
    filter_input_1_1 = buffer_data_4[4727:4704];
    filter_input_1_2 = blur5x5_1_dout[4727:4704];
    current_RowCol_1 = {img_addr, 10'd589};
  end
  else if (detected_keypoint[1][589]) begin
    filter_input_1_0 = buffer_data_5[4735:4712];
    filter_input_1_1 = buffer_data_4[4735:4712];
    filter_input_1_2 = blur5x5_1_dout[4735:4712];
    current_RowCol_1 = {img_addr, 10'd590};
  end
  else if (detected_keypoint[1][590]) begin
    filter_input_1_0 = buffer_data_5[4743:4720];
    filter_input_1_1 = buffer_data_4[4743:4720];
    filter_input_1_2 = blur5x5_1_dout[4743:4720];
    current_RowCol_1 = {img_addr, 10'd591};
  end
  else if (detected_keypoint[1][591]) begin
    filter_input_1_0 = buffer_data_5[4751:4728];
    filter_input_1_1 = buffer_data_4[4751:4728];
    filter_input_1_2 = blur5x5_1_dout[4751:4728];
    current_RowCol_1 = {img_addr, 10'd592};
  end
  else if (detected_keypoint[1][592]) begin
    filter_input_1_0 = buffer_data_5[4759:4736];
    filter_input_1_1 = buffer_data_4[4759:4736];
    filter_input_1_2 = blur5x5_1_dout[4759:4736];
    current_RowCol_1 = {img_addr, 10'd593};
  end
  else if (detected_keypoint[1][593]) begin
    filter_input_1_0 = buffer_data_5[4767:4744];
    filter_input_1_1 = buffer_data_4[4767:4744];
    filter_input_1_2 = blur5x5_1_dout[4767:4744];
    current_RowCol_1 = {img_addr, 10'd594};
  end
  else if (detected_keypoint[1][594]) begin
    filter_input_1_0 = buffer_data_5[4775:4752];
    filter_input_1_1 = buffer_data_4[4775:4752];
    filter_input_1_2 = blur5x5_1_dout[4775:4752];
    current_RowCol_1 = {img_addr, 10'd595};
  end
  else if (detected_keypoint[1][595]) begin
    filter_input_1_0 = buffer_data_5[4783:4760];
    filter_input_1_1 = buffer_data_4[4783:4760];
    filter_input_1_2 = blur5x5_1_dout[4783:4760];
    current_RowCol_1 = {img_addr, 10'd596};
  end
  else if (detected_keypoint[1][596]) begin
    filter_input_1_0 = buffer_data_5[4791:4768];
    filter_input_1_1 = buffer_data_4[4791:4768];
    filter_input_1_2 = blur5x5_1_dout[4791:4768];
    current_RowCol_1 = {img_addr, 10'd597};
  end
  else if (detected_keypoint[1][597]) begin
    filter_input_1_0 = buffer_data_5[4799:4776];
    filter_input_1_1 = buffer_data_4[4799:4776];
    filter_input_1_2 = blur5x5_1_dout[4799:4776];
    current_RowCol_1 = {img_addr, 10'd598};
  end
  else if (detected_keypoint[1][598]) begin
    filter_input_1_0 = buffer_data_5[4807:4784];
    filter_input_1_1 = buffer_data_4[4807:4784];
    filter_input_1_2 = blur5x5_1_dout[4807:4784];
    current_RowCol_1 = {img_addr, 10'd599};
  end
  else if (detected_keypoint[1][599]) begin
    filter_input_1_0 = buffer_data_5[4815:4792];
    filter_input_1_1 = buffer_data_4[4815:4792];
    filter_input_1_2 = blur5x5_1_dout[4815:4792];
    current_RowCol_1 = {img_addr, 10'd600};
  end
  else if (detected_keypoint[1][600]) begin
    filter_input_1_0 = buffer_data_5[4823:4800];
    filter_input_1_1 = buffer_data_4[4823:4800];
    filter_input_1_2 = blur5x5_1_dout[4823:4800];
    current_RowCol_1 = {img_addr, 10'd601};
  end
  else if (detected_keypoint[1][601]) begin
    filter_input_1_0 = buffer_data_5[4831:4808];
    filter_input_1_1 = buffer_data_4[4831:4808];
    filter_input_1_2 = blur5x5_1_dout[4831:4808];
    current_RowCol_1 = {img_addr, 10'd602};
  end
  else if (detected_keypoint[1][602]) begin
    filter_input_1_0 = buffer_data_5[4839:4816];
    filter_input_1_1 = buffer_data_4[4839:4816];
    filter_input_1_2 = blur5x5_1_dout[4839:4816];
    current_RowCol_1 = {img_addr, 10'd603};
  end
  else if (detected_keypoint[1][603]) begin
    filter_input_1_0 = buffer_data_5[4847:4824];
    filter_input_1_1 = buffer_data_4[4847:4824];
    filter_input_1_2 = blur5x5_1_dout[4847:4824];
    current_RowCol_1 = {img_addr, 10'd604};
  end
  else if (detected_keypoint[1][604]) begin
    filter_input_1_0 = buffer_data_5[4855:4832];
    filter_input_1_1 = buffer_data_4[4855:4832];
    filter_input_1_2 = blur5x5_1_dout[4855:4832];
    current_RowCol_1 = {img_addr, 10'd605};
  end
  else if (detected_keypoint[1][605]) begin
    filter_input_1_0 = buffer_data_5[4863:4840];
    filter_input_1_1 = buffer_data_4[4863:4840];
    filter_input_1_2 = blur5x5_1_dout[4863:4840];
    current_RowCol_1 = {img_addr, 10'd606};
  end
  else if (detected_keypoint[1][606]) begin
    filter_input_1_0 = buffer_data_5[4871:4848];
    filter_input_1_1 = buffer_data_4[4871:4848];
    filter_input_1_2 = blur5x5_1_dout[4871:4848];
    current_RowCol_1 = {img_addr, 10'd607};
  end
  else if (detected_keypoint[1][607]) begin
    filter_input_1_0 = buffer_data_5[4879:4856];
    filter_input_1_1 = buffer_data_4[4879:4856];
    filter_input_1_2 = blur5x5_1_dout[4879:4856];
    current_RowCol_1 = {img_addr, 10'd608};
  end
  else if (detected_keypoint[1][608]) begin
    filter_input_1_0 = buffer_data_5[4887:4864];
    filter_input_1_1 = buffer_data_4[4887:4864];
    filter_input_1_2 = blur5x5_1_dout[4887:4864];
    current_RowCol_1 = {img_addr, 10'd609};
  end
  else if (detected_keypoint[1][609]) begin
    filter_input_1_0 = buffer_data_5[4895:4872];
    filter_input_1_1 = buffer_data_4[4895:4872];
    filter_input_1_2 = blur5x5_1_dout[4895:4872];
    current_RowCol_1 = {img_addr, 10'd610};
  end
  else if (detected_keypoint[1][610]) begin
    filter_input_1_0 = buffer_data_5[4903:4880];
    filter_input_1_1 = buffer_data_4[4903:4880];
    filter_input_1_2 = blur5x5_1_dout[4903:4880];
    current_RowCol_1 = {img_addr, 10'd611};
  end
  else if (detected_keypoint[1][611]) begin
    filter_input_1_0 = buffer_data_5[4911:4888];
    filter_input_1_1 = buffer_data_4[4911:4888];
    filter_input_1_2 = blur5x5_1_dout[4911:4888];
    current_RowCol_1 = {img_addr, 10'd612};
  end
  else if (detected_keypoint[1][612]) begin
    filter_input_1_0 = buffer_data_5[4919:4896];
    filter_input_1_1 = buffer_data_4[4919:4896];
    filter_input_1_2 = blur5x5_1_dout[4919:4896];
    current_RowCol_1 = {img_addr, 10'd613};
  end
  else if (detected_keypoint[1][613]) begin
    filter_input_1_0 = buffer_data_5[4927:4904];
    filter_input_1_1 = buffer_data_4[4927:4904];
    filter_input_1_2 = blur5x5_1_dout[4927:4904];
    current_RowCol_1 = {img_addr, 10'd614};
  end
  else if (detected_keypoint[1][614]) begin
    filter_input_1_0 = buffer_data_5[4935:4912];
    filter_input_1_1 = buffer_data_4[4935:4912];
    filter_input_1_2 = blur5x5_1_dout[4935:4912];
    current_RowCol_1 = {img_addr, 10'd615};
  end
  else if (detected_keypoint[1][615]) begin
    filter_input_1_0 = buffer_data_5[4943:4920];
    filter_input_1_1 = buffer_data_4[4943:4920];
    filter_input_1_2 = blur5x5_1_dout[4943:4920];
    current_RowCol_1 = {img_addr, 10'd616};
  end
  else if (detected_keypoint[1][616]) begin
    filter_input_1_0 = buffer_data_5[4951:4928];
    filter_input_1_1 = buffer_data_4[4951:4928];
    filter_input_1_2 = blur5x5_1_dout[4951:4928];
    current_RowCol_1 = {img_addr, 10'd617};
  end
  else if (detected_keypoint[1][617]) begin
    filter_input_1_0 = buffer_data_5[4959:4936];
    filter_input_1_1 = buffer_data_4[4959:4936];
    filter_input_1_2 = blur5x5_1_dout[4959:4936];
    current_RowCol_1 = {img_addr, 10'd618};
  end
  else if (detected_keypoint[1][618]) begin
    filter_input_1_0 = buffer_data_5[4967:4944];
    filter_input_1_1 = buffer_data_4[4967:4944];
    filter_input_1_2 = blur5x5_1_dout[4967:4944];
    current_RowCol_1 = {img_addr, 10'd619};
  end
  else if (detected_keypoint[1][619]) begin
    filter_input_1_0 = buffer_data_5[4975:4952];
    filter_input_1_1 = buffer_data_4[4975:4952];
    filter_input_1_2 = blur5x5_1_dout[4975:4952];
    current_RowCol_1 = {img_addr, 10'd620};
  end
  else if (detected_keypoint[1][620]) begin
    filter_input_1_0 = buffer_data_5[4983:4960];
    filter_input_1_1 = buffer_data_4[4983:4960];
    filter_input_1_2 = blur5x5_1_dout[4983:4960];
    current_RowCol_1 = {img_addr, 10'd621};
  end
  else if (detected_keypoint[1][621]) begin
    filter_input_1_0 = buffer_data_5[4991:4968];
    filter_input_1_1 = buffer_data_4[4991:4968];
    filter_input_1_2 = blur5x5_1_dout[4991:4968];
    current_RowCol_1 = {img_addr, 10'd622};
  end
  else if (detected_keypoint[1][622]) begin
    filter_input_1_0 = buffer_data_5[4999:4976];
    filter_input_1_1 = buffer_data_4[4999:4976];
    filter_input_1_2 = blur5x5_1_dout[4999:4976];
    current_RowCol_1 = {img_addr, 10'd623};
  end
  else if (detected_keypoint[1][623]) begin
    filter_input_1_0 = buffer_data_5[5007:4984];
    filter_input_1_1 = buffer_data_4[5007:4984];
    filter_input_1_2 = blur5x5_1_dout[5007:4984];
    current_RowCol_1 = {img_addr, 10'd624};
  end
  else if (detected_keypoint[1][624]) begin
    filter_input_1_0 = buffer_data_5[5015:4992];
    filter_input_1_1 = buffer_data_4[5015:4992];
    filter_input_1_2 = blur5x5_1_dout[5015:4992];
    current_RowCol_1 = {img_addr, 10'd625};
  end
  else if (detected_keypoint[1][625]) begin
    filter_input_1_0 = buffer_data_5[5023:5000];
    filter_input_1_1 = buffer_data_4[5023:5000];
    filter_input_1_2 = blur5x5_1_dout[5023:5000];
    current_RowCol_1 = {img_addr, 10'd626};
  end
  else if (detected_keypoint[1][626]) begin
    filter_input_1_0 = buffer_data_5[5031:5008];
    filter_input_1_1 = buffer_data_4[5031:5008];
    filter_input_1_2 = blur5x5_1_dout[5031:5008];
    current_RowCol_1 = {img_addr, 10'd627};
  end
  else if (detected_keypoint[1][627]) begin
    filter_input_1_0 = buffer_data_5[5039:5016];
    filter_input_1_1 = buffer_data_4[5039:5016];
    filter_input_1_2 = blur5x5_1_dout[5039:5016];
    current_RowCol_1 = {img_addr, 10'd628};
  end
  else if (detected_keypoint[1][628]) begin
    filter_input_1_0 = buffer_data_5[5047:5024];
    filter_input_1_1 = buffer_data_4[5047:5024];
    filter_input_1_2 = blur5x5_1_dout[5047:5024];
    current_RowCol_1 = {img_addr, 10'd629};
  end
  else if (detected_keypoint[1][629]) begin
    filter_input_1_0 = buffer_data_5[5055:5032];
    filter_input_1_1 = buffer_data_4[5055:5032];
    filter_input_1_2 = blur5x5_1_dout[5055:5032];
    current_RowCol_1 = {img_addr, 10'd630};
  end
  else if (detected_keypoint[1][630]) begin
    filter_input_1_0 = buffer_data_5[5063:5040];
    filter_input_1_1 = buffer_data_4[5063:5040];
    filter_input_1_2 = blur5x5_1_dout[5063:5040];
    current_RowCol_1 = {img_addr, 10'd631};
  end
  else if (detected_keypoint[1][631]) begin
    filter_input_1_0 = buffer_data_5[5071:5048];
    filter_input_1_1 = buffer_data_4[5071:5048];
    filter_input_1_2 = blur5x5_1_dout[5071:5048];
    current_RowCol_1 = {img_addr, 10'd632};
  end
  else if (detected_keypoint[1][632]) begin
    filter_input_1_0 = buffer_data_5[5079:5056];
    filter_input_1_1 = buffer_data_4[5079:5056];
    filter_input_1_2 = blur5x5_1_dout[5079:5056];
    current_RowCol_1 = {img_addr, 10'd633};
  end
  else if (detected_keypoint[1][633]) begin
    filter_input_1_0 = buffer_data_5[5087:5064];
    filter_input_1_1 = buffer_data_4[5087:5064];
    filter_input_1_2 = blur5x5_1_dout[5087:5064];
    current_RowCol_1 = {img_addr, 10'd634};
  end
  else if (detected_keypoint[1][634]) begin
    filter_input_1_0 = buffer_data_5[5095:5072];
    filter_input_1_1 = buffer_data_4[5095:5072];
    filter_input_1_2 = blur5x5_1_dout[5095:5072];
    current_RowCol_1 = {img_addr, 10'd635};
  end
  else if (detected_keypoint[1][635]) begin
    filter_input_1_0 = buffer_data_5[5103:5080];
    filter_input_1_1 = buffer_data_4[5103:5080];
    filter_input_1_2 = blur5x5_1_dout[5103:5080];
    current_RowCol_1 = {img_addr, 10'd636};
  end
  else if (detected_keypoint[1][636]) begin
    filter_input_1_0 = buffer_data_5[5111:5088];
    filter_input_1_1 = buffer_data_4[5111:5088];
    filter_input_1_2 = blur5x5_1_dout[5111:5088];
    current_RowCol_1 = {img_addr, 10'd637};
  end
  else if (detected_keypoint[1][637]) begin
    filter_input_1_0 = buffer_data_5[5119:5096];
    filter_input_1_1 = buffer_data_4[5119:5096];
    filter_input_1_2 = blur5x5_1_dout[5119:5096];
    current_RowCol_1 = {img_addr, 10'd638};
  end
  else begin
    filter_input_1_0 = 'd0;
    filter_input_1_1 = 'd0;
    filter_input_1_2 = 'd0;
    current_RowCol_1 = 'd0;
  end

endmodule