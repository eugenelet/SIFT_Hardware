module Gaussian_Blur_5x5_1(
  clk,
  rst_n,
  buffer_data_0,
  buffer_data_1,
  buffer_data_2,
  buffer_data_3,
  buffer_data_4,
  current_state,
  blur_din
);

input                 clk;
input                 rst_n;
input         [3:0]   current_state;
input       [5119:0]   buffer_data_0;
input       [5119:0]   buffer_data_1;
input       [5119:0]   buffer_data_2;
input       [5119:0]   buffer_data_3;
input       [5119:0]   buffer_data_4;
output reg  [5119:0]  blur_din;

parameter ST_IDLE        = 0,
          ST_READY       = 1,/*Idle 1 state for SRAM to get READY*/
          ST_GAUSSIAN_0  = 2,
          ST_GAUSSIAN_1  = 3,
          ST_GAUSSIAN_2  = 4,
          ST_GAUSSIAN_3  = 5,
          ST_GAUSSIAN_4  = 6,
          ST_GAUSSIAN_5  = 7,
          ST_GAUSSIAN_6  = 8,
          ST_GAUSSIAN_7  = 9,
          ST_GAUSSIAN_8  = 10,
          ST_GAUSSIAN_9  = 11;

reg       [159:0]  G_Kernel_5x5[0:2];
always @(posedge clk) begin
  if (!rst_n) begin
    G_Kernel_5x5[0][31:0]  <= 32'h07E31AF6; //18'b000001111110001100;//'d030809;
    G_Kernel_5x5[0][63:32] <= 32'h0983EB80; //18'b000010011000001111;//'d037169;
    G_Kernel_5x5[0][95:64] <= 32'h0A212B91; //18'b000010100010000100;//'d039568;
    G_Kernel_5x5[0][127:96] <= 32'h0983EB80; //18'b000010011000001111;//'d037169;
    G_Kernel_5x5[0][159:128] <= 32'h07E31AF6; //18'b000001111110001100;//'d030809;
    G_Kernel_5x5[1][31:0]  <= 32'h0983EB80; //18'b000010011000001111;//'d037169;
    G_Kernel_5x5[1][63:32] <= 32'h0B7AC7A0; //18'b000010110111101011;//'d044842;
    G_Kernel_5x5[1][95:64] <= 32'h0C387DF7; //18'b000011000011100001;//'d047737;
    G_Kernel_5x5[1][127:96] <= 32'h0B7AC7A0; //18'b000010110111101011;//'d044842;
    G_Kernel_5x5[1][159:128] <= 32'h0983EB80; //18'b000010011000001111;//'d037169;
    G_Kernel_5x5[2][31:0]  <= 32'h0A212B91; //18'b000010100010000100;//'d039568;
    G_Kernel_5x5[2][63:32] <= 32'h0C387DF7; //18'b000011000011100001;//'d047737;
    G_Kernel_5x5[2][95:64] <= 32'h0D02737E; //18'b000011010000001001;//'d050818;
    G_Kernel_5x5[2][127:96] <= 32'h0C387DF7; //18'b000011000011100001;//'d047737;
    G_Kernel_5x5[2][159:128] <= 32'h0A212B91; //18'b000010100010000100;//'d039568;
  end
end

reg    [39:0]    layer0[0:63]; //wire
reg    [39:0]    layer1[0:63]; //wire
reg    [39:0]    layer2[0:63]; //wire
reg    [39:0]    layer3[0:63]; //wire
reg    [39:0]    layer4[0:63]; //wire
always @(*) begin
  case(current_state)
    ST_GAUSSIAN_0: begin
        layer0[0][7:0] = 0;
        layer0[0][15:8] = 0;
        layer0[0][23:16] = buffer_data_4[7:0];
        layer0[0][31:24] = buffer_data_4[15:8];
        layer0[0][39:32] = buffer_data_4[23:16];
        layer1[0][7:0] = 0;
        layer1[0][15:8] = 0;
        layer1[0][23:16] = buffer_data_3[7:0];
        layer1[0][31:24] = buffer_data_3[15:8];
        layer1[0][39:32] = buffer_data_3[23:16];
        layer2[0][7:0] = 0;
        layer2[0][15:8] = 0;
        layer2[0][23:16] = buffer_data_2[7:0];
        layer2[0][31:24] = buffer_data_2[15:8];
        layer2[0][39:32] = buffer_data_2[23:16];
        layer3[0][7:0] = 0;
        layer3[0][15:8] = 0;
        layer3[0][23:16] = buffer_data_1[7:0];
        layer3[0][31:24] = buffer_data_1[15:8];
        layer3[0][39:32] = buffer_data_1[23:16];
        layer4[0][7:0] = 0;
        layer4[0][15:8] = 0;
        layer4[0][23:16] = buffer_data_0[7:0];
        layer4[0][31:24] = buffer_data_0[15:8];
        layer4[0][39:32] = buffer_data_0[23:16];
        layer0[1][7:0] = 0;
        layer0[1][15:8] = buffer_data_4[7:0];
        layer0[1][23:16] = buffer_data_4[15:8];
        layer0[1][31:24] = buffer_data_4[23:16];
        layer0[1][39:32] = buffer_data_4[31:24];
        layer1[1][7:0] = 0;
        layer1[1][15:8] = buffer_data_3[7:0];
        layer1[1][23:16] = buffer_data_3[15:8];
        layer1[1][31:24] = buffer_data_3[23:16];
        layer1[1][39:32] = buffer_data_3[31:24];
        layer2[1][7:0] = 0;
        layer2[1][15:8] = buffer_data_2[7:0];
        layer2[1][23:16] = buffer_data_2[15:8];
        layer2[1][31:24] = buffer_data_2[23:16];
        layer2[1][39:32] = buffer_data_2[31:24];
        layer3[1][7:0] = 0;
        layer3[1][15:8] = buffer_data_1[7:0];
        layer3[1][23:16] = buffer_data_1[15:8];
        layer3[1][31:24] = buffer_data_1[23:16];
        layer3[1][39:32] = buffer_data_1[31:24];
        layer4[1][7:0] = 0;
        layer4[1][15:8] = buffer_data_0[7:0];
        layer4[1][23:16] = buffer_data_0[15:8];
        layer4[1][31:24] = buffer_data_0[23:16];
        layer4[1][39:32] = buffer_data_0[31:24];
        layer0[2][7:0] = buffer_data_4[7:0];
        layer0[2][15:8] = buffer_data_4[15:8];
        layer0[2][23:16] = buffer_data_4[23:16];
        layer0[2][31:24] = buffer_data_4[31:24];
        layer0[2][39:32] = buffer_data_4[39:32];
        layer1[2][7:0] = buffer_data_3[7:0];
        layer1[2][15:8] = buffer_data_3[15:8];
        layer1[2][23:16] = buffer_data_3[23:16];
        layer1[2][31:24] = buffer_data_3[31:24];
        layer1[2][39:32] = buffer_data_3[39:32];
        layer2[2][7:0] = buffer_data_2[7:0];
        layer2[2][15:8] = buffer_data_2[15:8];
        layer2[2][23:16] = buffer_data_2[23:16];
        layer2[2][31:24] = buffer_data_2[31:24];
        layer2[2][39:32] = buffer_data_2[39:32];
        layer3[2][7:0] = buffer_data_1[7:0];
        layer3[2][15:8] = buffer_data_1[15:8];
        layer3[2][23:16] = buffer_data_1[23:16];
        layer3[2][31:24] = buffer_data_1[31:24];
        layer3[2][39:32] = buffer_data_1[39:32];
        layer4[2][7:0] = buffer_data_0[7:0];
        layer4[2][15:8] = buffer_data_0[15:8];
        layer4[2][23:16] = buffer_data_0[23:16];
        layer4[2][31:24] = buffer_data_0[31:24];
        layer4[2][39:32] = buffer_data_0[39:32];
        layer0[3][7:0] = buffer_data_4[15:8];
        layer0[3][15:8] = buffer_data_4[23:16];
        layer0[3][23:16] = buffer_data_4[31:24];
        layer0[3][31:24] = buffer_data_4[39:32];
        layer0[3][39:32] = buffer_data_4[47:40];
        layer1[3][7:0] = buffer_data_3[15:8];
        layer1[3][15:8] = buffer_data_3[23:16];
        layer1[3][23:16] = buffer_data_3[31:24];
        layer1[3][31:24] = buffer_data_3[39:32];
        layer1[3][39:32] = buffer_data_3[47:40];
        layer2[3][7:0] = buffer_data_2[15:8];
        layer2[3][15:8] = buffer_data_2[23:16];
        layer2[3][23:16] = buffer_data_2[31:24];
        layer2[3][31:24] = buffer_data_2[39:32];
        layer2[3][39:32] = buffer_data_2[47:40];
        layer3[3][7:0] = buffer_data_1[15:8];
        layer3[3][15:8] = buffer_data_1[23:16];
        layer3[3][23:16] = buffer_data_1[31:24];
        layer3[3][31:24] = buffer_data_1[39:32];
        layer3[3][39:32] = buffer_data_1[47:40];
        layer4[3][7:0] = buffer_data_0[15:8];
        layer4[3][15:8] = buffer_data_0[23:16];
        layer4[3][23:16] = buffer_data_0[31:24];
        layer4[3][31:24] = buffer_data_0[39:32];
        layer4[3][39:32] = buffer_data_0[47:40];
        layer0[4][7:0] = buffer_data_4[23:16];
        layer0[4][15:8] = buffer_data_4[31:24];
        layer0[4][23:16] = buffer_data_4[39:32];
        layer0[4][31:24] = buffer_data_4[47:40];
        layer0[4][39:32] = buffer_data_4[55:48];
        layer1[4][7:0] = buffer_data_3[23:16];
        layer1[4][15:8] = buffer_data_3[31:24];
        layer1[4][23:16] = buffer_data_3[39:32];
        layer1[4][31:24] = buffer_data_3[47:40];
        layer1[4][39:32] = buffer_data_3[55:48];
        layer2[4][7:0] = buffer_data_2[23:16];
        layer2[4][15:8] = buffer_data_2[31:24];
        layer2[4][23:16] = buffer_data_2[39:32];
        layer2[4][31:24] = buffer_data_2[47:40];
        layer2[4][39:32] = buffer_data_2[55:48];
        layer3[4][7:0] = buffer_data_1[23:16];
        layer3[4][15:8] = buffer_data_1[31:24];
        layer3[4][23:16] = buffer_data_1[39:32];
        layer3[4][31:24] = buffer_data_1[47:40];
        layer3[4][39:32] = buffer_data_1[55:48];
        layer4[4][7:0] = buffer_data_0[23:16];
        layer4[4][15:8] = buffer_data_0[31:24];
        layer4[4][23:16] = buffer_data_0[39:32];
        layer4[4][31:24] = buffer_data_0[47:40];
        layer4[4][39:32] = buffer_data_0[55:48];
        layer0[5][7:0] = buffer_data_4[31:24];
        layer0[5][15:8] = buffer_data_4[39:32];
        layer0[5][23:16] = buffer_data_4[47:40];
        layer0[5][31:24] = buffer_data_4[55:48];
        layer0[5][39:32] = buffer_data_4[63:56];
        layer1[5][7:0] = buffer_data_3[31:24];
        layer1[5][15:8] = buffer_data_3[39:32];
        layer1[5][23:16] = buffer_data_3[47:40];
        layer1[5][31:24] = buffer_data_3[55:48];
        layer1[5][39:32] = buffer_data_3[63:56];
        layer2[5][7:0] = buffer_data_2[31:24];
        layer2[5][15:8] = buffer_data_2[39:32];
        layer2[5][23:16] = buffer_data_2[47:40];
        layer2[5][31:24] = buffer_data_2[55:48];
        layer2[5][39:32] = buffer_data_2[63:56];
        layer3[5][7:0] = buffer_data_1[31:24];
        layer3[5][15:8] = buffer_data_1[39:32];
        layer3[5][23:16] = buffer_data_1[47:40];
        layer3[5][31:24] = buffer_data_1[55:48];
        layer3[5][39:32] = buffer_data_1[63:56];
        layer4[5][7:0] = buffer_data_0[31:24];
        layer4[5][15:8] = buffer_data_0[39:32];
        layer4[5][23:16] = buffer_data_0[47:40];
        layer4[5][31:24] = buffer_data_0[55:48];
        layer4[5][39:32] = buffer_data_0[63:56];
        layer0[6][7:0] = buffer_data_4[39:32];
        layer0[6][15:8] = buffer_data_4[47:40];
        layer0[6][23:16] = buffer_data_4[55:48];
        layer0[6][31:24] = buffer_data_4[63:56];
        layer0[6][39:32] = buffer_data_4[71:64];
        layer1[6][7:0] = buffer_data_3[39:32];
        layer1[6][15:8] = buffer_data_3[47:40];
        layer1[6][23:16] = buffer_data_3[55:48];
        layer1[6][31:24] = buffer_data_3[63:56];
        layer1[6][39:32] = buffer_data_3[71:64];
        layer2[6][7:0] = buffer_data_2[39:32];
        layer2[6][15:8] = buffer_data_2[47:40];
        layer2[6][23:16] = buffer_data_2[55:48];
        layer2[6][31:24] = buffer_data_2[63:56];
        layer2[6][39:32] = buffer_data_2[71:64];
        layer3[6][7:0] = buffer_data_1[39:32];
        layer3[6][15:8] = buffer_data_1[47:40];
        layer3[6][23:16] = buffer_data_1[55:48];
        layer3[6][31:24] = buffer_data_1[63:56];
        layer3[6][39:32] = buffer_data_1[71:64];
        layer4[6][7:0] = buffer_data_0[39:32];
        layer4[6][15:8] = buffer_data_0[47:40];
        layer4[6][23:16] = buffer_data_0[55:48];
        layer4[6][31:24] = buffer_data_0[63:56];
        layer4[6][39:32] = buffer_data_0[71:64];
        layer0[7][7:0] = buffer_data_4[47:40];
        layer0[7][15:8] = buffer_data_4[55:48];
        layer0[7][23:16] = buffer_data_4[63:56];
        layer0[7][31:24] = buffer_data_4[71:64];
        layer0[7][39:32] = buffer_data_4[79:72];
        layer1[7][7:0] = buffer_data_3[47:40];
        layer1[7][15:8] = buffer_data_3[55:48];
        layer1[7][23:16] = buffer_data_3[63:56];
        layer1[7][31:24] = buffer_data_3[71:64];
        layer1[7][39:32] = buffer_data_3[79:72];
        layer2[7][7:0] = buffer_data_2[47:40];
        layer2[7][15:8] = buffer_data_2[55:48];
        layer2[7][23:16] = buffer_data_2[63:56];
        layer2[7][31:24] = buffer_data_2[71:64];
        layer2[7][39:32] = buffer_data_2[79:72];
        layer3[7][7:0] = buffer_data_1[47:40];
        layer3[7][15:8] = buffer_data_1[55:48];
        layer3[7][23:16] = buffer_data_1[63:56];
        layer3[7][31:24] = buffer_data_1[71:64];
        layer3[7][39:32] = buffer_data_1[79:72];
        layer4[7][7:0] = buffer_data_0[47:40];
        layer4[7][15:8] = buffer_data_0[55:48];
        layer4[7][23:16] = buffer_data_0[63:56];
        layer4[7][31:24] = buffer_data_0[71:64];
        layer4[7][39:32] = buffer_data_0[79:72];
        layer0[8][7:0] = buffer_data_4[55:48];
        layer0[8][15:8] = buffer_data_4[63:56];
        layer0[8][23:16] = buffer_data_4[71:64];
        layer0[8][31:24] = buffer_data_4[79:72];
        layer0[8][39:32] = buffer_data_4[87:80];
        layer1[8][7:0] = buffer_data_3[55:48];
        layer1[8][15:8] = buffer_data_3[63:56];
        layer1[8][23:16] = buffer_data_3[71:64];
        layer1[8][31:24] = buffer_data_3[79:72];
        layer1[8][39:32] = buffer_data_3[87:80];
        layer2[8][7:0] = buffer_data_2[55:48];
        layer2[8][15:8] = buffer_data_2[63:56];
        layer2[8][23:16] = buffer_data_2[71:64];
        layer2[8][31:24] = buffer_data_2[79:72];
        layer2[8][39:32] = buffer_data_2[87:80];
        layer3[8][7:0] = buffer_data_1[55:48];
        layer3[8][15:8] = buffer_data_1[63:56];
        layer3[8][23:16] = buffer_data_1[71:64];
        layer3[8][31:24] = buffer_data_1[79:72];
        layer3[8][39:32] = buffer_data_1[87:80];
        layer4[8][7:0] = buffer_data_0[55:48];
        layer4[8][15:8] = buffer_data_0[63:56];
        layer4[8][23:16] = buffer_data_0[71:64];
        layer4[8][31:24] = buffer_data_0[79:72];
        layer4[8][39:32] = buffer_data_0[87:80];
        layer0[9][7:0] = buffer_data_4[63:56];
        layer0[9][15:8] = buffer_data_4[71:64];
        layer0[9][23:16] = buffer_data_4[79:72];
        layer0[9][31:24] = buffer_data_4[87:80];
        layer0[9][39:32] = buffer_data_4[95:88];
        layer1[9][7:0] = buffer_data_3[63:56];
        layer1[9][15:8] = buffer_data_3[71:64];
        layer1[9][23:16] = buffer_data_3[79:72];
        layer1[9][31:24] = buffer_data_3[87:80];
        layer1[9][39:32] = buffer_data_3[95:88];
        layer2[9][7:0] = buffer_data_2[63:56];
        layer2[9][15:8] = buffer_data_2[71:64];
        layer2[9][23:16] = buffer_data_2[79:72];
        layer2[9][31:24] = buffer_data_2[87:80];
        layer2[9][39:32] = buffer_data_2[95:88];
        layer3[9][7:0] = buffer_data_1[63:56];
        layer3[9][15:8] = buffer_data_1[71:64];
        layer3[9][23:16] = buffer_data_1[79:72];
        layer3[9][31:24] = buffer_data_1[87:80];
        layer3[9][39:32] = buffer_data_1[95:88];
        layer4[9][7:0] = buffer_data_0[63:56];
        layer4[9][15:8] = buffer_data_0[71:64];
        layer4[9][23:16] = buffer_data_0[79:72];
        layer4[9][31:24] = buffer_data_0[87:80];
        layer4[9][39:32] = buffer_data_0[95:88];
        layer0[10][7:0] = buffer_data_4[71:64];
        layer0[10][15:8] = buffer_data_4[79:72];
        layer0[10][23:16] = buffer_data_4[87:80];
        layer0[10][31:24] = buffer_data_4[95:88];
        layer0[10][39:32] = buffer_data_4[103:96];
        layer1[10][7:0] = buffer_data_3[71:64];
        layer1[10][15:8] = buffer_data_3[79:72];
        layer1[10][23:16] = buffer_data_3[87:80];
        layer1[10][31:24] = buffer_data_3[95:88];
        layer1[10][39:32] = buffer_data_3[103:96];
        layer2[10][7:0] = buffer_data_2[71:64];
        layer2[10][15:8] = buffer_data_2[79:72];
        layer2[10][23:16] = buffer_data_2[87:80];
        layer2[10][31:24] = buffer_data_2[95:88];
        layer2[10][39:32] = buffer_data_2[103:96];
        layer3[10][7:0] = buffer_data_1[71:64];
        layer3[10][15:8] = buffer_data_1[79:72];
        layer3[10][23:16] = buffer_data_1[87:80];
        layer3[10][31:24] = buffer_data_1[95:88];
        layer3[10][39:32] = buffer_data_1[103:96];
        layer4[10][7:0] = buffer_data_0[71:64];
        layer4[10][15:8] = buffer_data_0[79:72];
        layer4[10][23:16] = buffer_data_0[87:80];
        layer4[10][31:24] = buffer_data_0[95:88];
        layer4[10][39:32] = buffer_data_0[103:96];
        layer0[11][7:0] = buffer_data_4[79:72];
        layer0[11][15:8] = buffer_data_4[87:80];
        layer0[11][23:16] = buffer_data_4[95:88];
        layer0[11][31:24] = buffer_data_4[103:96];
        layer0[11][39:32] = buffer_data_4[111:104];
        layer1[11][7:0] = buffer_data_3[79:72];
        layer1[11][15:8] = buffer_data_3[87:80];
        layer1[11][23:16] = buffer_data_3[95:88];
        layer1[11][31:24] = buffer_data_3[103:96];
        layer1[11][39:32] = buffer_data_3[111:104];
        layer2[11][7:0] = buffer_data_2[79:72];
        layer2[11][15:8] = buffer_data_2[87:80];
        layer2[11][23:16] = buffer_data_2[95:88];
        layer2[11][31:24] = buffer_data_2[103:96];
        layer2[11][39:32] = buffer_data_2[111:104];
        layer3[11][7:0] = buffer_data_1[79:72];
        layer3[11][15:8] = buffer_data_1[87:80];
        layer3[11][23:16] = buffer_data_1[95:88];
        layer3[11][31:24] = buffer_data_1[103:96];
        layer3[11][39:32] = buffer_data_1[111:104];
        layer4[11][7:0] = buffer_data_0[79:72];
        layer4[11][15:8] = buffer_data_0[87:80];
        layer4[11][23:16] = buffer_data_0[95:88];
        layer4[11][31:24] = buffer_data_0[103:96];
        layer4[11][39:32] = buffer_data_0[111:104];
        layer0[12][7:0] = buffer_data_4[87:80];
        layer0[12][15:8] = buffer_data_4[95:88];
        layer0[12][23:16] = buffer_data_4[103:96];
        layer0[12][31:24] = buffer_data_4[111:104];
        layer0[12][39:32] = buffer_data_4[119:112];
        layer1[12][7:0] = buffer_data_3[87:80];
        layer1[12][15:8] = buffer_data_3[95:88];
        layer1[12][23:16] = buffer_data_3[103:96];
        layer1[12][31:24] = buffer_data_3[111:104];
        layer1[12][39:32] = buffer_data_3[119:112];
        layer2[12][7:0] = buffer_data_2[87:80];
        layer2[12][15:8] = buffer_data_2[95:88];
        layer2[12][23:16] = buffer_data_2[103:96];
        layer2[12][31:24] = buffer_data_2[111:104];
        layer2[12][39:32] = buffer_data_2[119:112];
        layer3[12][7:0] = buffer_data_1[87:80];
        layer3[12][15:8] = buffer_data_1[95:88];
        layer3[12][23:16] = buffer_data_1[103:96];
        layer3[12][31:24] = buffer_data_1[111:104];
        layer3[12][39:32] = buffer_data_1[119:112];
        layer4[12][7:0] = buffer_data_0[87:80];
        layer4[12][15:8] = buffer_data_0[95:88];
        layer4[12][23:16] = buffer_data_0[103:96];
        layer4[12][31:24] = buffer_data_0[111:104];
        layer4[12][39:32] = buffer_data_0[119:112];
        layer0[13][7:0] = buffer_data_4[95:88];
        layer0[13][15:8] = buffer_data_4[103:96];
        layer0[13][23:16] = buffer_data_4[111:104];
        layer0[13][31:24] = buffer_data_4[119:112];
        layer0[13][39:32] = buffer_data_4[127:120];
        layer1[13][7:0] = buffer_data_3[95:88];
        layer1[13][15:8] = buffer_data_3[103:96];
        layer1[13][23:16] = buffer_data_3[111:104];
        layer1[13][31:24] = buffer_data_3[119:112];
        layer1[13][39:32] = buffer_data_3[127:120];
        layer2[13][7:0] = buffer_data_2[95:88];
        layer2[13][15:8] = buffer_data_2[103:96];
        layer2[13][23:16] = buffer_data_2[111:104];
        layer2[13][31:24] = buffer_data_2[119:112];
        layer2[13][39:32] = buffer_data_2[127:120];
        layer3[13][7:0] = buffer_data_1[95:88];
        layer3[13][15:8] = buffer_data_1[103:96];
        layer3[13][23:16] = buffer_data_1[111:104];
        layer3[13][31:24] = buffer_data_1[119:112];
        layer3[13][39:32] = buffer_data_1[127:120];
        layer4[13][7:0] = buffer_data_0[95:88];
        layer4[13][15:8] = buffer_data_0[103:96];
        layer4[13][23:16] = buffer_data_0[111:104];
        layer4[13][31:24] = buffer_data_0[119:112];
        layer4[13][39:32] = buffer_data_0[127:120];
        layer0[14][7:0] = buffer_data_4[103:96];
        layer0[14][15:8] = buffer_data_4[111:104];
        layer0[14][23:16] = buffer_data_4[119:112];
        layer0[14][31:24] = buffer_data_4[127:120];
        layer0[14][39:32] = buffer_data_4[135:128];
        layer1[14][7:0] = buffer_data_3[103:96];
        layer1[14][15:8] = buffer_data_3[111:104];
        layer1[14][23:16] = buffer_data_3[119:112];
        layer1[14][31:24] = buffer_data_3[127:120];
        layer1[14][39:32] = buffer_data_3[135:128];
        layer2[14][7:0] = buffer_data_2[103:96];
        layer2[14][15:8] = buffer_data_2[111:104];
        layer2[14][23:16] = buffer_data_2[119:112];
        layer2[14][31:24] = buffer_data_2[127:120];
        layer2[14][39:32] = buffer_data_2[135:128];
        layer3[14][7:0] = buffer_data_1[103:96];
        layer3[14][15:8] = buffer_data_1[111:104];
        layer3[14][23:16] = buffer_data_1[119:112];
        layer3[14][31:24] = buffer_data_1[127:120];
        layer3[14][39:32] = buffer_data_1[135:128];
        layer4[14][7:0] = buffer_data_0[103:96];
        layer4[14][15:8] = buffer_data_0[111:104];
        layer4[14][23:16] = buffer_data_0[119:112];
        layer4[14][31:24] = buffer_data_0[127:120];
        layer4[14][39:32] = buffer_data_0[135:128];
        layer0[15][7:0] = buffer_data_4[111:104];
        layer0[15][15:8] = buffer_data_4[119:112];
        layer0[15][23:16] = buffer_data_4[127:120];
        layer0[15][31:24] = buffer_data_4[135:128];
        layer0[15][39:32] = buffer_data_4[143:136];
        layer1[15][7:0] = buffer_data_3[111:104];
        layer1[15][15:8] = buffer_data_3[119:112];
        layer1[15][23:16] = buffer_data_3[127:120];
        layer1[15][31:24] = buffer_data_3[135:128];
        layer1[15][39:32] = buffer_data_3[143:136];
        layer2[15][7:0] = buffer_data_2[111:104];
        layer2[15][15:8] = buffer_data_2[119:112];
        layer2[15][23:16] = buffer_data_2[127:120];
        layer2[15][31:24] = buffer_data_2[135:128];
        layer2[15][39:32] = buffer_data_2[143:136];
        layer3[15][7:0] = buffer_data_1[111:104];
        layer3[15][15:8] = buffer_data_1[119:112];
        layer3[15][23:16] = buffer_data_1[127:120];
        layer3[15][31:24] = buffer_data_1[135:128];
        layer3[15][39:32] = buffer_data_1[143:136];
        layer4[15][7:0] = buffer_data_0[111:104];
        layer4[15][15:8] = buffer_data_0[119:112];
        layer4[15][23:16] = buffer_data_0[127:120];
        layer4[15][31:24] = buffer_data_0[135:128];
        layer4[15][39:32] = buffer_data_0[143:136];
        layer0[16][7:0] = buffer_data_4[119:112];
        layer0[16][15:8] = buffer_data_4[127:120];
        layer0[16][23:16] = buffer_data_4[135:128];
        layer0[16][31:24] = buffer_data_4[143:136];
        layer0[16][39:32] = buffer_data_4[151:144];
        layer1[16][7:0] = buffer_data_3[119:112];
        layer1[16][15:8] = buffer_data_3[127:120];
        layer1[16][23:16] = buffer_data_3[135:128];
        layer1[16][31:24] = buffer_data_3[143:136];
        layer1[16][39:32] = buffer_data_3[151:144];
        layer2[16][7:0] = buffer_data_2[119:112];
        layer2[16][15:8] = buffer_data_2[127:120];
        layer2[16][23:16] = buffer_data_2[135:128];
        layer2[16][31:24] = buffer_data_2[143:136];
        layer2[16][39:32] = buffer_data_2[151:144];
        layer3[16][7:0] = buffer_data_1[119:112];
        layer3[16][15:8] = buffer_data_1[127:120];
        layer3[16][23:16] = buffer_data_1[135:128];
        layer3[16][31:24] = buffer_data_1[143:136];
        layer3[16][39:32] = buffer_data_1[151:144];
        layer4[16][7:0] = buffer_data_0[119:112];
        layer4[16][15:8] = buffer_data_0[127:120];
        layer4[16][23:16] = buffer_data_0[135:128];
        layer4[16][31:24] = buffer_data_0[143:136];
        layer4[16][39:32] = buffer_data_0[151:144];
        layer0[17][7:0] = buffer_data_4[127:120];
        layer0[17][15:8] = buffer_data_4[135:128];
        layer0[17][23:16] = buffer_data_4[143:136];
        layer0[17][31:24] = buffer_data_4[151:144];
        layer0[17][39:32] = buffer_data_4[159:152];
        layer1[17][7:0] = buffer_data_3[127:120];
        layer1[17][15:8] = buffer_data_3[135:128];
        layer1[17][23:16] = buffer_data_3[143:136];
        layer1[17][31:24] = buffer_data_3[151:144];
        layer1[17][39:32] = buffer_data_3[159:152];
        layer2[17][7:0] = buffer_data_2[127:120];
        layer2[17][15:8] = buffer_data_2[135:128];
        layer2[17][23:16] = buffer_data_2[143:136];
        layer2[17][31:24] = buffer_data_2[151:144];
        layer2[17][39:32] = buffer_data_2[159:152];
        layer3[17][7:0] = buffer_data_1[127:120];
        layer3[17][15:8] = buffer_data_1[135:128];
        layer3[17][23:16] = buffer_data_1[143:136];
        layer3[17][31:24] = buffer_data_1[151:144];
        layer3[17][39:32] = buffer_data_1[159:152];
        layer4[17][7:0] = buffer_data_0[127:120];
        layer4[17][15:8] = buffer_data_0[135:128];
        layer4[17][23:16] = buffer_data_0[143:136];
        layer4[17][31:24] = buffer_data_0[151:144];
        layer4[17][39:32] = buffer_data_0[159:152];
        layer0[18][7:0] = buffer_data_4[135:128];
        layer0[18][15:8] = buffer_data_4[143:136];
        layer0[18][23:16] = buffer_data_4[151:144];
        layer0[18][31:24] = buffer_data_4[159:152];
        layer0[18][39:32] = buffer_data_4[167:160];
        layer1[18][7:0] = buffer_data_3[135:128];
        layer1[18][15:8] = buffer_data_3[143:136];
        layer1[18][23:16] = buffer_data_3[151:144];
        layer1[18][31:24] = buffer_data_3[159:152];
        layer1[18][39:32] = buffer_data_3[167:160];
        layer2[18][7:0] = buffer_data_2[135:128];
        layer2[18][15:8] = buffer_data_2[143:136];
        layer2[18][23:16] = buffer_data_2[151:144];
        layer2[18][31:24] = buffer_data_2[159:152];
        layer2[18][39:32] = buffer_data_2[167:160];
        layer3[18][7:0] = buffer_data_1[135:128];
        layer3[18][15:8] = buffer_data_1[143:136];
        layer3[18][23:16] = buffer_data_1[151:144];
        layer3[18][31:24] = buffer_data_1[159:152];
        layer3[18][39:32] = buffer_data_1[167:160];
        layer4[18][7:0] = buffer_data_0[135:128];
        layer4[18][15:8] = buffer_data_0[143:136];
        layer4[18][23:16] = buffer_data_0[151:144];
        layer4[18][31:24] = buffer_data_0[159:152];
        layer4[18][39:32] = buffer_data_0[167:160];
        layer0[19][7:0] = buffer_data_4[143:136];
        layer0[19][15:8] = buffer_data_4[151:144];
        layer0[19][23:16] = buffer_data_4[159:152];
        layer0[19][31:24] = buffer_data_4[167:160];
        layer0[19][39:32] = buffer_data_4[175:168];
        layer1[19][7:0] = buffer_data_3[143:136];
        layer1[19][15:8] = buffer_data_3[151:144];
        layer1[19][23:16] = buffer_data_3[159:152];
        layer1[19][31:24] = buffer_data_3[167:160];
        layer1[19][39:32] = buffer_data_3[175:168];
        layer2[19][7:0] = buffer_data_2[143:136];
        layer2[19][15:8] = buffer_data_2[151:144];
        layer2[19][23:16] = buffer_data_2[159:152];
        layer2[19][31:24] = buffer_data_2[167:160];
        layer2[19][39:32] = buffer_data_2[175:168];
        layer3[19][7:0] = buffer_data_1[143:136];
        layer3[19][15:8] = buffer_data_1[151:144];
        layer3[19][23:16] = buffer_data_1[159:152];
        layer3[19][31:24] = buffer_data_1[167:160];
        layer3[19][39:32] = buffer_data_1[175:168];
        layer4[19][7:0] = buffer_data_0[143:136];
        layer4[19][15:8] = buffer_data_0[151:144];
        layer4[19][23:16] = buffer_data_0[159:152];
        layer4[19][31:24] = buffer_data_0[167:160];
        layer4[19][39:32] = buffer_data_0[175:168];
        layer0[20][7:0] = buffer_data_4[151:144];
        layer0[20][15:8] = buffer_data_4[159:152];
        layer0[20][23:16] = buffer_data_4[167:160];
        layer0[20][31:24] = buffer_data_4[175:168];
        layer0[20][39:32] = buffer_data_4[183:176];
        layer1[20][7:0] = buffer_data_3[151:144];
        layer1[20][15:8] = buffer_data_3[159:152];
        layer1[20][23:16] = buffer_data_3[167:160];
        layer1[20][31:24] = buffer_data_3[175:168];
        layer1[20][39:32] = buffer_data_3[183:176];
        layer2[20][7:0] = buffer_data_2[151:144];
        layer2[20][15:8] = buffer_data_2[159:152];
        layer2[20][23:16] = buffer_data_2[167:160];
        layer2[20][31:24] = buffer_data_2[175:168];
        layer2[20][39:32] = buffer_data_2[183:176];
        layer3[20][7:0] = buffer_data_1[151:144];
        layer3[20][15:8] = buffer_data_1[159:152];
        layer3[20][23:16] = buffer_data_1[167:160];
        layer3[20][31:24] = buffer_data_1[175:168];
        layer3[20][39:32] = buffer_data_1[183:176];
        layer4[20][7:0] = buffer_data_0[151:144];
        layer4[20][15:8] = buffer_data_0[159:152];
        layer4[20][23:16] = buffer_data_0[167:160];
        layer4[20][31:24] = buffer_data_0[175:168];
        layer4[20][39:32] = buffer_data_0[183:176];
        layer0[21][7:0] = buffer_data_4[159:152];
        layer0[21][15:8] = buffer_data_4[167:160];
        layer0[21][23:16] = buffer_data_4[175:168];
        layer0[21][31:24] = buffer_data_4[183:176];
        layer0[21][39:32] = buffer_data_4[191:184];
        layer1[21][7:0] = buffer_data_3[159:152];
        layer1[21][15:8] = buffer_data_3[167:160];
        layer1[21][23:16] = buffer_data_3[175:168];
        layer1[21][31:24] = buffer_data_3[183:176];
        layer1[21][39:32] = buffer_data_3[191:184];
        layer2[21][7:0] = buffer_data_2[159:152];
        layer2[21][15:8] = buffer_data_2[167:160];
        layer2[21][23:16] = buffer_data_2[175:168];
        layer2[21][31:24] = buffer_data_2[183:176];
        layer2[21][39:32] = buffer_data_2[191:184];
        layer3[21][7:0] = buffer_data_1[159:152];
        layer3[21][15:8] = buffer_data_1[167:160];
        layer3[21][23:16] = buffer_data_1[175:168];
        layer3[21][31:24] = buffer_data_1[183:176];
        layer3[21][39:32] = buffer_data_1[191:184];
        layer4[21][7:0] = buffer_data_0[159:152];
        layer4[21][15:8] = buffer_data_0[167:160];
        layer4[21][23:16] = buffer_data_0[175:168];
        layer4[21][31:24] = buffer_data_0[183:176];
        layer4[21][39:32] = buffer_data_0[191:184];
        layer0[22][7:0] = buffer_data_4[167:160];
        layer0[22][15:8] = buffer_data_4[175:168];
        layer0[22][23:16] = buffer_data_4[183:176];
        layer0[22][31:24] = buffer_data_4[191:184];
        layer0[22][39:32] = buffer_data_4[199:192];
        layer1[22][7:0] = buffer_data_3[167:160];
        layer1[22][15:8] = buffer_data_3[175:168];
        layer1[22][23:16] = buffer_data_3[183:176];
        layer1[22][31:24] = buffer_data_3[191:184];
        layer1[22][39:32] = buffer_data_3[199:192];
        layer2[22][7:0] = buffer_data_2[167:160];
        layer2[22][15:8] = buffer_data_2[175:168];
        layer2[22][23:16] = buffer_data_2[183:176];
        layer2[22][31:24] = buffer_data_2[191:184];
        layer2[22][39:32] = buffer_data_2[199:192];
        layer3[22][7:0] = buffer_data_1[167:160];
        layer3[22][15:8] = buffer_data_1[175:168];
        layer3[22][23:16] = buffer_data_1[183:176];
        layer3[22][31:24] = buffer_data_1[191:184];
        layer3[22][39:32] = buffer_data_1[199:192];
        layer4[22][7:0] = buffer_data_0[167:160];
        layer4[22][15:8] = buffer_data_0[175:168];
        layer4[22][23:16] = buffer_data_0[183:176];
        layer4[22][31:24] = buffer_data_0[191:184];
        layer4[22][39:32] = buffer_data_0[199:192];
        layer0[23][7:0] = buffer_data_4[175:168];
        layer0[23][15:8] = buffer_data_4[183:176];
        layer0[23][23:16] = buffer_data_4[191:184];
        layer0[23][31:24] = buffer_data_4[199:192];
        layer0[23][39:32] = buffer_data_4[207:200];
        layer1[23][7:0] = buffer_data_3[175:168];
        layer1[23][15:8] = buffer_data_3[183:176];
        layer1[23][23:16] = buffer_data_3[191:184];
        layer1[23][31:24] = buffer_data_3[199:192];
        layer1[23][39:32] = buffer_data_3[207:200];
        layer2[23][7:0] = buffer_data_2[175:168];
        layer2[23][15:8] = buffer_data_2[183:176];
        layer2[23][23:16] = buffer_data_2[191:184];
        layer2[23][31:24] = buffer_data_2[199:192];
        layer2[23][39:32] = buffer_data_2[207:200];
        layer3[23][7:0] = buffer_data_1[175:168];
        layer3[23][15:8] = buffer_data_1[183:176];
        layer3[23][23:16] = buffer_data_1[191:184];
        layer3[23][31:24] = buffer_data_1[199:192];
        layer3[23][39:32] = buffer_data_1[207:200];
        layer4[23][7:0] = buffer_data_0[175:168];
        layer4[23][15:8] = buffer_data_0[183:176];
        layer4[23][23:16] = buffer_data_0[191:184];
        layer4[23][31:24] = buffer_data_0[199:192];
        layer4[23][39:32] = buffer_data_0[207:200];
        layer0[24][7:0] = buffer_data_4[183:176];
        layer0[24][15:8] = buffer_data_4[191:184];
        layer0[24][23:16] = buffer_data_4[199:192];
        layer0[24][31:24] = buffer_data_4[207:200];
        layer0[24][39:32] = buffer_data_4[215:208];
        layer1[24][7:0] = buffer_data_3[183:176];
        layer1[24][15:8] = buffer_data_3[191:184];
        layer1[24][23:16] = buffer_data_3[199:192];
        layer1[24][31:24] = buffer_data_3[207:200];
        layer1[24][39:32] = buffer_data_3[215:208];
        layer2[24][7:0] = buffer_data_2[183:176];
        layer2[24][15:8] = buffer_data_2[191:184];
        layer2[24][23:16] = buffer_data_2[199:192];
        layer2[24][31:24] = buffer_data_2[207:200];
        layer2[24][39:32] = buffer_data_2[215:208];
        layer3[24][7:0] = buffer_data_1[183:176];
        layer3[24][15:8] = buffer_data_1[191:184];
        layer3[24][23:16] = buffer_data_1[199:192];
        layer3[24][31:24] = buffer_data_1[207:200];
        layer3[24][39:32] = buffer_data_1[215:208];
        layer4[24][7:0] = buffer_data_0[183:176];
        layer4[24][15:8] = buffer_data_0[191:184];
        layer4[24][23:16] = buffer_data_0[199:192];
        layer4[24][31:24] = buffer_data_0[207:200];
        layer4[24][39:32] = buffer_data_0[215:208];
        layer0[25][7:0] = buffer_data_4[191:184];
        layer0[25][15:8] = buffer_data_4[199:192];
        layer0[25][23:16] = buffer_data_4[207:200];
        layer0[25][31:24] = buffer_data_4[215:208];
        layer0[25][39:32] = buffer_data_4[223:216];
        layer1[25][7:0] = buffer_data_3[191:184];
        layer1[25][15:8] = buffer_data_3[199:192];
        layer1[25][23:16] = buffer_data_3[207:200];
        layer1[25][31:24] = buffer_data_3[215:208];
        layer1[25][39:32] = buffer_data_3[223:216];
        layer2[25][7:0] = buffer_data_2[191:184];
        layer2[25][15:8] = buffer_data_2[199:192];
        layer2[25][23:16] = buffer_data_2[207:200];
        layer2[25][31:24] = buffer_data_2[215:208];
        layer2[25][39:32] = buffer_data_2[223:216];
        layer3[25][7:0] = buffer_data_1[191:184];
        layer3[25][15:8] = buffer_data_1[199:192];
        layer3[25][23:16] = buffer_data_1[207:200];
        layer3[25][31:24] = buffer_data_1[215:208];
        layer3[25][39:32] = buffer_data_1[223:216];
        layer4[25][7:0] = buffer_data_0[191:184];
        layer4[25][15:8] = buffer_data_0[199:192];
        layer4[25][23:16] = buffer_data_0[207:200];
        layer4[25][31:24] = buffer_data_0[215:208];
        layer4[25][39:32] = buffer_data_0[223:216];
        layer0[26][7:0] = buffer_data_4[199:192];
        layer0[26][15:8] = buffer_data_4[207:200];
        layer0[26][23:16] = buffer_data_4[215:208];
        layer0[26][31:24] = buffer_data_4[223:216];
        layer0[26][39:32] = buffer_data_4[231:224];
        layer1[26][7:0] = buffer_data_3[199:192];
        layer1[26][15:8] = buffer_data_3[207:200];
        layer1[26][23:16] = buffer_data_3[215:208];
        layer1[26][31:24] = buffer_data_3[223:216];
        layer1[26][39:32] = buffer_data_3[231:224];
        layer2[26][7:0] = buffer_data_2[199:192];
        layer2[26][15:8] = buffer_data_2[207:200];
        layer2[26][23:16] = buffer_data_2[215:208];
        layer2[26][31:24] = buffer_data_2[223:216];
        layer2[26][39:32] = buffer_data_2[231:224];
        layer3[26][7:0] = buffer_data_1[199:192];
        layer3[26][15:8] = buffer_data_1[207:200];
        layer3[26][23:16] = buffer_data_1[215:208];
        layer3[26][31:24] = buffer_data_1[223:216];
        layer3[26][39:32] = buffer_data_1[231:224];
        layer4[26][7:0] = buffer_data_0[199:192];
        layer4[26][15:8] = buffer_data_0[207:200];
        layer4[26][23:16] = buffer_data_0[215:208];
        layer4[26][31:24] = buffer_data_0[223:216];
        layer4[26][39:32] = buffer_data_0[231:224];
        layer0[27][7:0] = buffer_data_4[207:200];
        layer0[27][15:8] = buffer_data_4[215:208];
        layer0[27][23:16] = buffer_data_4[223:216];
        layer0[27][31:24] = buffer_data_4[231:224];
        layer0[27][39:32] = buffer_data_4[239:232];
        layer1[27][7:0] = buffer_data_3[207:200];
        layer1[27][15:8] = buffer_data_3[215:208];
        layer1[27][23:16] = buffer_data_3[223:216];
        layer1[27][31:24] = buffer_data_3[231:224];
        layer1[27][39:32] = buffer_data_3[239:232];
        layer2[27][7:0] = buffer_data_2[207:200];
        layer2[27][15:8] = buffer_data_2[215:208];
        layer2[27][23:16] = buffer_data_2[223:216];
        layer2[27][31:24] = buffer_data_2[231:224];
        layer2[27][39:32] = buffer_data_2[239:232];
        layer3[27][7:0] = buffer_data_1[207:200];
        layer3[27][15:8] = buffer_data_1[215:208];
        layer3[27][23:16] = buffer_data_1[223:216];
        layer3[27][31:24] = buffer_data_1[231:224];
        layer3[27][39:32] = buffer_data_1[239:232];
        layer4[27][7:0] = buffer_data_0[207:200];
        layer4[27][15:8] = buffer_data_0[215:208];
        layer4[27][23:16] = buffer_data_0[223:216];
        layer4[27][31:24] = buffer_data_0[231:224];
        layer4[27][39:32] = buffer_data_0[239:232];
        layer0[28][7:0] = buffer_data_4[215:208];
        layer0[28][15:8] = buffer_data_4[223:216];
        layer0[28][23:16] = buffer_data_4[231:224];
        layer0[28][31:24] = buffer_data_4[239:232];
        layer0[28][39:32] = buffer_data_4[247:240];
        layer1[28][7:0] = buffer_data_3[215:208];
        layer1[28][15:8] = buffer_data_3[223:216];
        layer1[28][23:16] = buffer_data_3[231:224];
        layer1[28][31:24] = buffer_data_3[239:232];
        layer1[28][39:32] = buffer_data_3[247:240];
        layer2[28][7:0] = buffer_data_2[215:208];
        layer2[28][15:8] = buffer_data_2[223:216];
        layer2[28][23:16] = buffer_data_2[231:224];
        layer2[28][31:24] = buffer_data_2[239:232];
        layer2[28][39:32] = buffer_data_2[247:240];
        layer3[28][7:0] = buffer_data_1[215:208];
        layer3[28][15:8] = buffer_data_1[223:216];
        layer3[28][23:16] = buffer_data_1[231:224];
        layer3[28][31:24] = buffer_data_1[239:232];
        layer3[28][39:32] = buffer_data_1[247:240];
        layer4[28][7:0] = buffer_data_0[215:208];
        layer4[28][15:8] = buffer_data_0[223:216];
        layer4[28][23:16] = buffer_data_0[231:224];
        layer4[28][31:24] = buffer_data_0[239:232];
        layer4[28][39:32] = buffer_data_0[247:240];
        layer0[29][7:0] = buffer_data_4[223:216];
        layer0[29][15:8] = buffer_data_4[231:224];
        layer0[29][23:16] = buffer_data_4[239:232];
        layer0[29][31:24] = buffer_data_4[247:240];
        layer0[29][39:32] = buffer_data_4[255:248];
        layer1[29][7:0] = buffer_data_3[223:216];
        layer1[29][15:8] = buffer_data_3[231:224];
        layer1[29][23:16] = buffer_data_3[239:232];
        layer1[29][31:24] = buffer_data_3[247:240];
        layer1[29][39:32] = buffer_data_3[255:248];
        layer2[29][7:0] = buffer_data_2[223:216];
        layer2[29][15:8] = buffer_data_2[231:224];
        layer2[29][23:16] = buffer_data_2[239:232];
        layer2[29][31:24] = buffer_data_2[247:240];
        layer2[29][39:32] = buffer_data_2[255:248];
        layer3[29][7:0] = buffer_data_1[223:216];
        layer3[29][15:8] = buffer_data_1[231:224];
        layer3[29][23:16] = buffer_data_1[239:232];
        layer3[29][31:24] = buffer_data_1[247:240];
        layer3[29][39:32] = buffer_data_1[255:248];
        layer4[29][7:0] = buffer_data_0[223:216];
        layer4[29][15:8] = buffer_data_0[231:224];
        layer4[29][23:16] = buffer_data_0[239:232];
        layer4[29][31:24] = buffer_data_0[247:240];
        layer4[29][39:32] = buffer_data_0[255:248];
        layer0[30][7:0] = buffer_data_4[231:224];
        layer0[30][15:8] = buffer_data_4[239:232];
        layer0[30][23:16] = buffer_data_4[247:240];
        layer0[30][31:24] = buffer_data_4[255:248];
        layer0[30][39:32] = buffer_data_4[263:256];
        layer1[30][7:0] = buffer_data_3[231:224];
        layer1[30][15:8] = buffer_data_3[239:232];
        layer1[30][23:16] = buffer_data_3[247:240];
        layer1[30][31:24] = buffer_data_3[255:248];
        layer1[30][39:32] = buffer_data_3[263:256];
        layer2[30][7:0] = buffer_data_2[231:224];
        layer2[30][15:8] = buffer_data_2[239:232];
        layer2[30][23:16] = buffer_data_2[247:240];
        layer2[30][31:24] = buffer_data_2[255:248];
        layer2[30][39:32] = buffer_data_2[263:256];
        layer3[30][7:0] = buffer_data_1[231:224];
        layer3[30][15:8] = buffer_data_1[239:232];
        layer3[30][23:16] = buffer_data_1[247:240];
        layer3[30][31:24] = buffer_data_1[255:248];
        layer3[30][39:32] = buffer_data_1[263:256];
        layer4[30][7:0] = buffer_data_0[231:224];
        layer4[30][15:8] = buffer_data_0[239:232];
        layer4[30][23:16] = buffer_data_0[247:240];
        layer4[30][31:24] = buffer_data_0[255:248];
        layer4[30][39:32] = buffer_data_0[263:256];
        layer0[31][7:0] = buffer_data_4[239:232];
        layer0[31][15:8] = buffer_data_4[247:240];
        layer0[31][23:16] = buffer_data_4[255:248];
        layer0[31][31:24] = buffer_data_4[263:256];
        layer0[31][39:32] = buffer_data_4[271:264];
        layer1[31][7:0] = buffer_data_3[239:232];
        layer1[31][15:8] = buffer_data_3[247:240];
        layer1[31][23:16] = buffer_data_3[255:248];
        layer1[31][31:24] = buffer_data_3[263:256];
        layer1[31][39:32] = buffer_data_3[271:264];
        layer2[31][7:0] = buffer_data_2[239:232];
        layer2[31][15:8] = buffer_data_2[247:240];
        layer2[31][23:16] = buffer_data_2[255:248];
        layer2[31][31:24] = buffer_data_2[263:256];
        layer2[31][39:32] = buffer_data_2[271:264];
        layer3[31][7:0] = buffer_data_1[239:232];
        layer3[31][15:8] = buffer_data_1[247:240];
        layer3[31][23:16] = buffer_data_1[255:248];
        layer3[31][31:24] = buffer_data_1[263:256];
        layer3[31][39:32] = buffer_data_1[271:264];
        layer4[31][7:0] = buffer_data_0[239:232];
        layer4[31][15:8] = buffer_data_0[247:240];
        layer4[31][23:16] = buffer_data_0[255:248];
        layer4[31][31:24] = buffer_data_0[263:256];
        layer4[31][39:32] = buffer_data_0[271:264];
        layer0[32][7:0] = buffer_data_4[247:240];
        layer0[32][15:8] = buffer_data_4[255:248];
        layer0[32][23:16] = buffer_data_4[263:256];
        layer0[32][31:24] = buffer_data_4[271:264];
        layer0[32][39:32] = buffer_data_4[279:272];
        layer1[32][7:0] = buffer_data_3[247:240];
        layer1[32][15:8] = buffer_data_3[255:248];
        layer1[32][23:16] = buffer_data_3[263:256];
        layer1[32][31:24] = buffer_data_3[271:264];
        layer1[32][39:32] = buffer_data_3[279:272];
        layer2[32][7:0] = buffer_data_2[247:240];
        layer2[32][15:8] = buffer_data_2[255:248];
        layer2[32][23:16] = buffer_data_2[263:256];
        layer2[32][31:24] = buffer_data_2[271:264];
        layer2[32][39:32] = buffer_data_2[279:272];
        layer3[32][7:0] = buffer_data_1[247:240];
        layer3[32][15:8] = buffer_data_1[255:248];
        layer3[32][23:16] = buffer_data_1[263:256];
        layer3[32][31:24] = buffer_data_1[271:264];
        layer3[32][39:32] = buffer_data_1[279:272];
        layer4[32][7:0] = buffer_data_0[247:240];
        layer4[32][15:8] = buffer_data_0[255:248];
        layer4[32][23:16] = buffer_data_0[263:256];
        layer4[32][31:24] = buffer_data_0[271:264];
        layer4[32][39:32] = buffer_data_0[279:272];
        layer0[33][7:0] = buffer_data_4[255:248];
        layer0[33][15:8] = buffer_data_4[263:256];
        layer0[33][23:16] = buffer_data_4[271:264];
        layer0[33][31:24] = buffer_data_4[279:272];
        layer0[33][39:32] = buffer_data_4[287:280];
        layer1[33][7:0] = buffer_data_3[255:248];
        layer1[33][15:8] = buffer_data_3[263:256];
        layer1[33][23:16] = buffer_data_3[271:264];
        layer1[33][31:24] = buffer_data_3[279:272];
        layer1[33][39:32] = buffer_data_3[287:280];
        layer2[33][7:0] = buffer_data_2[255:248];
        layer2[33][15:8] = buffer_data_2[263:256];
        layer2[33][23:16] = buffer_data_2[271:264];
        layer2[33][31:24] = buffer_data_2[279:272];
        layer2[33][39:32] = buffer_data_2[287:280];
        layer3[33][7:0] = buffer_data_1[255:248];
        layer3[33][15:8] = buffer_data_1[263:256];
        layer3[33][23:16] = buffer_data_1[271:264];
        layer3[33][31:24] = buffer_data_1[279:272];
        layer3[33][39:32] = buffer_data_1[287:280];
        layer4[33][7:0] = buffer_data_0[255:248];
        layer4[33][15:8] = buffer_data_0[263:256];
        layer4[33][23:16] = buffer_data_0[271:264];
        layer4[33][31:24] = buffer_data_0[279:272];
        layer4[33][39:32] = buffer_data_0[287:280];
        layer0[34][7:0] = buffer_data_4[263:256];
        layer0[34][15:8] = buffer_data_4[271:264];
        layer0[34][23:16] = buffer_data_4[279:272];
        layer0[34][31:24] = buffer_data_4[287:280];
        layer0[34][39:32] = buffer_data_4[295:288];
        layer1[34][7:0] = buffer_data_3[263:256];
        layer1[34][15:8] = buffer_data_3[271:264];
        layer1[34][23:16] = buffer_data_3[279:272];
        layer1[34][31:24] = buffer_data_3[287:280];
        layer1[34][39:32] = buffer_data_3[295:288];
        layer2[34][7:0] = buffer_data_2[263:256];
        layer2[34][15:8] = buffer_data_2[271:264];
        layer2[34][23:16] = buffer_data_2[279:272];
        layer2[34][31:24] = buffer_data_2[287:280];
        layer2[34][39:32] = buffer_data_2[295:288];
        layer3[34][7:0] = buffer_data_1[263:256];
        layer3[34][15:8] = buffer_data_1[271:264];
        layer3[34][23:16] = buffer_data_1[279:272];
        layer3[34][31:24] = buffer_data_1[287:280];
        layer3[34][39:32] = buffer_data_1[295:288];
        layer4[34][7:0] = buffer_data_0[263:256];
        layer4[34][15:8] = buffer_data_0[271:264];
        layer4[34][23:16] = buffer_data_0[279:272];
        layer4[34][31:24] = buffer_data_0[287:280];
        layer4[34][39:32] = buffer_data_0[295:288];
        layer0[35][7:0] = buffer_data_4[271:264];
        layer0[35][15:8] = buffer_data_4[279:272];
        layer0[35][23:16] = buffer_data_4[287:280];
        layer0[35][31:24] = buffer_data_4[295:288];
        layer0[35][39:32] = buffer_data_4[303:296];
        layer1[35][7:0] = buffer_data_3[271:264];
        layer1[35][15:8] = buffer_data_3[279:272];
        layer1[35][23:16] = buffer_data_3[287:280];
        layer1[35][31:24] = buffer_data_3[295:288];
        layer1[35][39:32] = buffer_data_3[303:296];
        layer2[35][7:0] = buffer_data_2[271:264];
        layer2[35][15:8] = buffer_data_2[279:272];
        layer2[35][23:16] = buffer_data_2[287:280];
        layer2[35][31:24] = buffer_data_2[295:288];
        layer2[35][39:32] = buffer_data_2[303:296];
        layer3[35][7:0] = buffer_data_1[271:264];
        layer3[35][15:8] = buffer_data_1[279:272];
        layer3[35][23:16] = buffer_data_1[287:280];
        layer3[35][31:24] = buffer_data_1[295:288];
        layer3[35][39:32] = buffer_data_1[303:296];
        layer4[35][7:0] = buffer_data_0[271:264];
        layer4[35][15:8] = buffer_data_0[279:272];
        layer4[35][23:16] = buffer_data_0[287:280];
        layer4[35][31:24] = buffer_data_0[295:288];
        layer4[35][39:32] = buffer_data_0[303:296];
        layer0[36][7:0] = buffer_data_4[279:272];
        layer0[36][15:8] = buffer_data_4[287:280];
        layer0[36][23:16] = buffer_data_4[295:288];
        layer0[36][31:24] = buffer_data_4[303:296];
        layer0[36][39:32] = buffer_data_4[311:304];
        layer1[36][7:0] = buffer_data_3[279:272];
        layer1[36][15:8] = buffer_data_3[287:280];
        layer1[36][23:16] = buffer_data_3[295:288];
        layer1[36][31:24] = buffer_data_3[303:296];
        layer1[36][39:32] = buffer_data_3[311:304];
        layer2[36][7:0] = buffer_data_2[279:272];
        layer2[36][15:8] = buffer_data_2[287:280];
        layer2[36][23:16] = buffer_data_2[295:288];
        layer2[36][31:24] = buffer_data_2[303:296];
        layer2[36][39:32] = buffer_data_2[311:304];
        layer3[36][7:0] = buffer_data_1[279:272];
        layer3[36][15:8] = buffer_data_1[287:280];
        layer3[36][23:16] = buffer_data_1[295:288];
        layer3[36][31:24] = buffer_data_1[303:296];
        layer3[36][39:32] = buffer_data_1[311:304];
        layer4[36][7:0] = buffer_data_0[279:272];
        layer4[36][15:8] = buffer_data_0[287:280];
        layer4[36][23:16] = buffer_data_0[295:288];
        layer4[36][31:24] = buffer_data_0[303:296];
        layer4[36][39:32] = buffer_data_0[311:304];
        layer0[37][7:0] = buffer_data_4[287:280];
        layer0[37][15:8] = buffer_data_4[295:288];
        layer0[37][23:16] = buffer_data_4[303:296];
        layer0[37][31:24] = buffer_data_4[311:304];
        layer0[37][39:32] = buffer_data_4[319:312];
        layer1[37][7:0] = buffer_data_3[287:280];
        layer1[37][15:8] = buffer_data_3[295:288];
        layer1[37][23:16] = buffer_data_3[303:296];
        layer1[37][31:24] = buffer_data_3[311:304];
        layer1[37][39:32] = buffer_data_3[319:312];
        layer2[37][7:0] = buffer_data_2[287:280];
        layer2[37][15:8] = buffer_data_2[295:288];
        layer2[37][23:16] = buffer_data_2[303:296];
        layer2[37][31:24] = buffer_data_2[311:304];
        layer2[37][39:32] = buffer_data_2[319:312];
        layer3[37][7:0] = buffer_data_1[287:280];
        layer3[37][15:8] = buffer_data_1[295:288];
        layer3[37][23:16] = buffer_data_1[303:296];
        layer3[37][31:24] = buffer_data_1[311:304];
        layer3[37][39:32] = buffer_data_1[319:312];
        layer4[37][7:0] = buffer_data_0[287:280];
        layer4[37][15:8] = buffer_data_0[295:288];
        layer4[37][23:16] = buffer_data_0[303:296];
        layer4[37][31:24] = buffer_data_0[311:304];
        layer4[37][39:32] = buffer_data_0[319:312];
        layer0[38][7:0] = buffer_data_4[295:288];
        layer0[38][15:8] = buffer_data_4[303:296];
        layer0[38][23:16] = buffer_data_4[311:304];
        layer0[38][31:24] = buffer_data_4[319:312];
        layer0[38][39:32] = buffer_data_4[327:320];
        layer1[38][7:0] = buffer_data_3[295:288];
        layer1[38][15:8] = buffer_data_3[303:296];
        layer1[38][23:16] = buffer_data_3[311:304];
        layer1[38][31:24] = buffer_data_3[319:312];
        layer1[38][39:32] = buffer_data_3[327:320];
        layer2[38][7:0] = buffer_data_2[295:288];
        layer2[38][15:8] = buffer_data_2[303:296];
        layer2[38][23:16] = buffer_data_2[311:304];
        layer2[38][31:24] = buffer_data_2[319:312];
        layer2[38][39:32] = buffer_data_2[327:320];
        layer3[38][7:0] = buffer_data_1[295:288];
        layer3[38][15:8] = buffer_data_1[303:296];
        layer3[38][23:16] = buffer_data_1[311:304];
        layer3[38][31:24] = buffer_data_1[319:312];
        layer3[38][39:32] = buffer_data_1[327:320];
        layer4[38][7:0] = buffer_data_0[295:288];
        layer4[38][15:8] = buffer_data_0[303:296];
        layer4[38][23:16] = buffer_data_0[311:304];
        layer4[38][31:24] = buffer_data_0[319:312];
        layer4[38][39:32] = buffer_data_0[327:320];
        layer0[39][7:0] = buffer_data_4[303:296];
        layer0[39][15:8] = buffer_data_4[311:304];
        layer0[39][23:16] = buffer_data_4[319:312];
        layer0[39][31:24] = buffer_data_4[327:320];
        layer0[39][39:32] = buffer_data_4[335:328];
        layer1[39][7:0] = buffer_data_3[303:296];
        layer1[39][15:8] = buffer_data_3[311:304];
        layer1[39][23:16] = buffer_data_3[319:312];
        layer1[39][31:24] = buffer_data_3[327:320];
        layer1[39][39:32] = buffer_data_3[335:328];
        layer2[39][7:0] = buffer_data_2[303:296];
        layer2[39][15:8] = buffer_data_2[311:304];
        layer2[39][23:16] = buffer_data_2[319:312];
        layer2[39][31:24] = buffer_data_2[327:320];
        layer2[39][39:32] = buffer_data_2[335:328];
        layer3[39][7:0] = buffer_data_1[303:296];
        layer3[39][15:8] = buffer_data_1[311:304];
        layer3[39][23:16] = buffer_data_1[319:312];
        layer3[39][31:24] = buffer_data_1[327:320];
        layer3[39][39:32] = buffer_data_1[335:328];
        layer4[39][7:0] = buffer_data_0[303:296];
        layer4[39][15:8] = buffer_data_0[311:304];
        layer4[39][23:16] = buffer_data_0[319:312];
        layer4[39][31:24] = buffer_data_0[327:320];
        layer4[39][39:32] = buffer_data_0[335:328];
        layer0[40][7:0] = buffer_data_4[311:304];
        layer0[40][15:8] = buffer_data_4[319:312];
        layer0[40][23:16] = buffer_data_4[327:320];
        layer0[40][31:24] = buffer_data_4[335:328];
        layer0[40][39:32] = buffer_data_4[343:336];
        layer1[40][7:0] = buffer_data_3[311:304];
        layer1[40][15:8] = buffer_data_3[319:312];
        layer1[40][23:16] = buffer_data_3[327:320];
        layer1[40][31:24] = buffer_data_3[335:328];
        layer1[40][39:32] = buffer_data_3[343:336];
        layer2[40][7:0] = buffer_data_2[311:304];
        layer2[40][15:8] = buffer_data_2[319:312];
        layer2[40][23:16] = buffer_data_2[327:320];
        layer2[40][31:24] = buffer_data_2[335:328];
        layer2[40][39:32] = buffer_data_2[343:336];
        layer3[40][7:0] = buffer_data_1[311:304];
        layer3[40][15:8] = buffer_data_1[319:312];
        layer3[40][23:16] = buffer_data_1[327:320];
        layer3[40][31:24] = buffer_data_1[335:328];
        layer3[40][39:32] = buffer_data_1[343:336];
        layer4[40][7:0] = buffer_data_0[311:304];
        layer4[40][15:8] = buffer_data_0[319:312];
        layer4[40][23:16] = buffer_data_0[327:320];
        layer4[40][31:24] = buffer_data_0[335:328];
        layer4[40][39:32] = buffer_data_0[343:336];
        layer0[41][7:0] = buffer_data_4[319:312];
        layer0[41][15:8] = buffer_data_4[327:320];
        layer0[41][23:16] = buffer_data_4[335:328];
        layer0[41][31:24] = buffer_data_4[343:336];
        layer0[41][39:32] = buffer_data_4[351:344];
        layer1[41][7:0] = buffer_data_3[319:312];
        layer1[41][15:8] = buffer_data_3[327:320];
        layer1[41][23:16] = buffer_data_3[335:328];
        layer1[41][31:24] = buffer_data_3[343:336];
        layer1[41][39:32] = buffer_data_3[351:344];
        layer2[41][7:0] = buffer_data_2[319:312];
        layer2[41][15:8] = buffer_data_2[327:320];
        layer2[41][23:16] = buffer_data_2[335:328];
        layer2[41][31:24] = buffer_data_2[343:336];
        layer2[41][39:32] = buffer_data_2[351:344];
        layer3[41][7:0] = buffer_data_1[319:312];
        layer3[41][15:8] = buffer_data_1[327:320];
        layer3[41][23:16] = buffer_data_1[335:328];
        layer3[41][31:24] = buffer_data_1[343:336];
        layer3[41][39:32] = buffer_data_1[351:344];
        layer4[41][7:0] = buffer_data_0[319:312];
        layer4[41][15:8] = buffer_data_0[327:320];
        layer4[41][23:16] = buffer_data_0[335:328];
        layer4[41][31:24] = buffer_data_0[343:336];
        layer4[41][39:32] = buffer_data_0[351:344];
        layer0[42][7:0] = buffer_data_4[327:320];
        layer0[42][15:8] = buffer_data_4[335:328];
        layer0[42][23:16] = buffer_data_4[343:336];
        layer0[42][31:24] = buffer_data_4[351:344];
        layer0[42][39:32] = buffer_data_4[359:352];
        layer1[42][7:0] = buffer_data_3[327:320];
        layer1[42][15:8] = buffer_data_3[335:328];
        layer1[42][23:16] = buffer_data_3[343:336];
        layer1[42][31:24] = buffer_data_3[351:344];
        layer1[42][39:32] = buffer_data_3[359:352];
        layer2[42][7:0] = buffer_data_2[327:320];
        layer2[42][15:8] = buffer_data_2[335:328];
        layer2[42][23:16] = buffer_data_2[343:336];
        layer2[42][31:24] = buffer_data_2[351:344];
        layer2[42][39:32] = buffer_data_2[359:352];
        layer3[42][7:0] = buffer_data_1[327:320];
        layer3[42][15:8] = buffer_data_1[335:328];
        layer3[42][23:16] = buffer_data_1[343:336];
        layer3[42][31:24] = buffer_data_1[351:344];
        layer3[42][39:32] = buffer_data_1[359:352];
        layer4[42][7:0] = buffer_data_0[327:320];
        layer4[42][15:8] = buffer_data_0[335:328];
        layer4[42][23:16] = buffer_data_0[343:336];
        layer4[42][31:24] = buffer_data_0[351:344];
        layer4[42][39:32] = buffer_data_0[359:352];
        layer0[43][7:0] = buffer_data_4[335:328];
        layer0[43][15:8] = buffer_data_4[343:336];
        layer0[43][23:16] = buffer_data_4[351:344];
        layer0[43][31:24] = buffer_data_4[359:352];
        layer0[43][39:32] = buffer_data_4[367:360];
        layer1[43][7:0] = buffer_data_3[335:328];
        layer1[43][15:8] = buffer_data_3[343:336];
        layer1[43][23:16] = buffer_data_3[351:344];
        layer1[43][31:24] = buffer_data_3[359:352];
        layer1[43][39:32] = buffer_data_3[367:360];
        layer2[43][7:0] = buffer_data_2[335:328];
        layer2[43][15:8] = buffer_data_2[343:336];
        layer2[43][23:16] = buffer_data_2[351:344];
        layer2[43][31:24] = buffer_data_2[359:352];
        layer2[43][39:32] = buffer_data_2[367:360];
        layer3[43][7:0] = buffer_data_1[335:328];
        layer3[43][15:8] = buffer_data_1[343:336];
        layer3[43][23:16] = buffer_data_1[351:344];
        layer3[43][31:24] = buffer_data_1[359:352];
        layer3[43][39:32] = buffer_data_1[367:360];
        layer4[43][7:0] = buffer_data_0[335:328];
        layer4[43][15:8] = buffer_data_0[343:336];
        layer4[43][23:16] = buffer_data_0[351:344];
        layer4[43][31:24] = buffer_data_0[359:352];
        layer4[43][39:32] = buffer_data_0[367:360];
        layer0[44][7:0] = buffer_data_4[343:336];
        layer0[44][15:8] = buffer_data_4[351:344];
        layer0[44][23:16] = buffer_data_4[359:352];
        layer0[44][31:24] = buffer_data_4[367:360];
        layer0[44][39:32] = buffer_data_4[375:368];
        layer1[44][7:0] = buffer_data_3[343:336];
        layer1[44][15:8] = buffer_data_3[351:344];
        layer1[44][23:16] = buffer_data_3[359:352];
        layer1[44][31:24] = buffer_data_3[367:360];
        layer1[44][39:32] = buffer_data_3[375:368];
        layer2[44][7:0] = buffer_data_2[343:336];
        layer2[44][15:8] = buffer_data_2[351:344];
        layer2[44][23:16] = buffer_data_2[359:352];
        layer2[44][31:24] = buffer_data_2[367:360];
        layer2[44][39:32] = buffer_data_2[375:368];
        layer3[44][7:0] = buffer_data_1[343:336];
        layer3[44][15:8] = buffer_data_1[351:344];
        layer3[44][23:16] = buffer_data_1[359:352];
        layer3[44][31:24] = buffer_data_1[367:360];
        layer3[44][39:32] = buffer_data_1[375:368];
        layer4[44][7:0] = buffer_data_0[343:336];
        layer4[44][15:8] = buffer_data_0[351:344];
        layer4[44][23:16] = buffer_data_0[359:352];
        layer4[44][31:24] = buffer_data_0[367:360];
        layer4[44][39:32] = buffer_data_0[375:368];
        layer0[45][7:0] = buffer_data_4[351:344];
        layer0[45][15:8] = buffer_data_4[359:352];
        layer0[45][23:16] = buffer_data_4[367:360];
        layer0[45][31:24] = buffer_data_4[375:368];
        layer0[45][39:32] = buffer_data_4[383:376];
        layer1[45][7:0] = buffer_data_3[351:344];
        layer1[45][15:8] = buffer_data_3[359:352];
        layer1[45][23:16] = buffer_data_3[367:360];
        layer1[45][31:24] = buffer_data_3[375:368];
        layer1[45][39:32] = buffer_data_3[383:376];
        layer2[45][7:0] = buffer_data_2[351:344];
        layer2[45][15:8] = buffer_data_2[359:352];
        layer2[45][23:16] = buffer_data_2[367:360];
        layer2[45][31:24] = buffer_data_2[375:368];
        layer2[45][39:32] = buffer_data_2[383:376];
        layer3[45][7:0] = buffer_data_1[351:344];
        layer3[45][15:8] = buffer_data_1[359:352];
        layer3[45][23:16] = buffer_data_1[367:360];
        layer3[45][31:24] = buffer_data_1[375:368];
        layer3[45][39:32] = buffer_data_1[383:376];
        layer4[45][7:0] = buffer_data_0[351:344];
        layer4[45][15:8] = buffer_data_0[359:352];
        layer4[45][23:16] = buffer_data_0[367:360];
        layer4[45][31:24] = buffer_data_0[375:368];
        layer4[45][39:32] = buffer_data_0[383:376];
        layer0[46][7:0] = buffer_data_4[359:352];
        layer0[46][15:8] = buffer_data_4[367:360];
        layer0[46][23:16] = buffer_data_4[375:368];
        layer0[46][31:24] = buffer_data_4[383:376];
        layer0[46][39:32] = buffer_data_4[391:384];
        layer1[46][7:0] = buffer_data_3[359:352];
        layer1[46][15:8] = buffer_data_3[367:360];
        layer1[46][23:16] = buffer_data_3[375:368];
        layer1[46][31:24] = buffer_data_3[383:376];
        layer1[46][39:32] = buffer_data_3[391:384];
        layer2[46][7:0] = buffer_data_2[359:352];
        layer2[46][15:8] = buffer_data_2[367:360];
        layer2[46][23:16] = buffer_data_2[375:368];
        layer2[46][31:24] = buffer_data_2[383:376];
        layer2[46][39:32] = buffer_data_2[391:384];
        layer3[46][7:0] = buffer_data_1[359:352];
        layer3[46][15:8] = buffer_data_1[367:360];
        layer3[46][23:16] = buffer_data_1[375:368];
        layer3[46][31:24] = buffer_data_1[383:376];
        layer3[46][39:32] = buffer_data_1[391:384];
        layer4[46][7:0] = buffer_data_0[359:352];
        layer4[46][15:8] = buffer_data_0[367:360];
        layer4[46][23:16] = buffer_data_0[375:368];
        layer4[46][31:24] = buffer_data_0[383:376];
        layer4[46][39:32] = buffer_data_0[391:384];
        layer0[47][7:0] = buffer_data_4[367:360];
        layer0[47][15:8] = buffer_data_4[375:368];
        layer0[47][23:16] = buffer_data_4[383:376];
        layer0[47][31:24] = buffer_data_4[391:384];
        layer0[47][39:32] = buffer_data_4[399:392];
        layer1[47][7:0] = buffer_data_3[367:360];
        layer1[47][15:8] = buffer_data_3[375:368];
        layer1[47][23:16] = buffer_data_3[383:376];
        layer1[47][31:24] = buffer_data_3[391:384];
        layer1[47][39:32] = buffer_data_3[399:392];
        layer2[47][7:0] = buffer_data_2[367:360];
        layer2[47][15:8] = buffer_data_2[375:368];
        layer2[47][23:16] = buffer_data_2[383:376];
        layer2[47][31:24] = buffer_data_2[391:384];
        layer2[47][39:32] = buffer_data_2[399:392];
        layer3[47][7:0] = buffer_data_1[367:360];
        layer3[47][15:8] = buffer_data_1[375:368];
        layer3[47][23:16] = buffer_data_1[383:376];
        layer3[47][31:24] = buffer_data_1[391:384];
        layer3[47][39:32] = buffer_data_1[399:392];
        layer4[47][7:0] = buffer_data_0[367:360];
        layer4[47][15:8] = buffer_data_0[375:368];
        layer4[47][23:16] = buffer_data_0[383:376];
        layer4[47][31:24] = buffer_data_0[391:384];
        layer4[47][39:32] = buffer_data_0[399:392];
        layer0[48][7:0] = buffer_data_4[375:368];
        layer0[48][15:8] = buffer_data_4[383:376];
        layer0[48][23:16] = buffer_data_4[391:384];
        layer0[48][31:24] = buffer_data_4[399:392];
        layer0[48][39:32] = buffer_data_4[407:400];
        layer1[48][7:0] = buffer_data_3[375:368];
        layer1[48][15:8] = buffer_data_3[383:376];
        layer1[48][23:16] = buffer_data_3[391:384];
        layer1[48][31:24] = buffer_data_3[399:392];
        layer1[48][39:32] = buffer_data_3[407:400];
        layer2[48][7:0] = buffer_data_2[375:368];
        layer2[48][15:8] = buffer_data_2[383:376];
        layer2[48][23:16] = buffer_data_2[391:384];
        layer2[48][31:24] = buffer_data_2[399:392];
        layer2[48][39:32] = buffer_data_2[407:400];
        layer3[48][7:0] = buffer_data_1[375:368];
        layer3[48][15:8] = buffer_data_1[383:376];
        layer3[48][23:16] = buffer_data_1[391:384];
        layer3[48][31:24] = buffer_data_1[399:392];
        layer3[48][39:32] = buffer_data_1[407:400];
        layer4[48][7:0] = buffer_data_0[375:368];
        layer4[48][15:8] = buffer_data_0[383:376];
        layer4[48][23:16] = buffer_data_0[391:384];
        layer4[48][31:24] = buffer_data_0[399:392];
        layer4[48][39:32] = buffer_data_0[407:400];
        layer0[49][7:0] = buffer_data_4[383:376];
        layer0[49][15:8] = buffer_data_4[391:384];
        layer0[49][23:16] = buffer_data_4[399:392];
        layer0[49][31:24] = buffer_data_4[407:400];
        layer0[49][39:32] = buffer_data_4[415:408];
        layer1[49][7:0] = buffer_data_3[383:376];
        layer1[49][15:8] = buffer_data_3[391:384];
        layer1[49][23:16] = buffer_data_3[399:392];
        layer1[49][31:24] = buffer_data_3[407:400];
        layer1[49][39:32] = buffer_data_3[415:408];
        layer2[49][7:0] = buffer_data_2[383:376];
        layer2[49][15:8] = buffer_data_2[391:384];
        layer2[49][23:16] = buffer_data_2[399:392];
        layer2[49][31:24] = buffer_data_2[407:400];
        layer2[49][39:32] = buffer_data_2[415:408];
        layer3[49][7:0] = buffer_data_1[383:376];
        layer3[49][15:8] = buffer_data_1[391:384];
        layer3[49][23:16] = buffer_data_1[399:392];
        layer3[49][31:24] = buffer_data_1[407:400];
        layer3[49][39:32] = buffer_data_1[415:408];
        layer4[49][7:0] = buffer_data_0[383:376];
        layer4[49][15:8] = buffer_data_0[391:384];
        layer4[49][23:16] = buffer_data_0[399:392];
        layer4[49][31:24] = buffer_data_0[407:400];
        layer4[49][39:32] = buffer_data_0[415:408];
        layer0[50][7:0] = buffer_data_4[391:384];
        layer0[50][15:8] = buffer_data_4[399:392];
        layer0[50][23:16] = buffer_data_4[407:400];
        layer0[50][31:24] = buffer_data_4[415:408];
        layer0[50][39:32] = buffer_data_4[423:416];
        layer1[50][7:0] = buffer_data_3[391:384];
        layer1[50][15:8] = buffer_data_3[399:392];
        layer1[50][23:16] = buffer_data_3[407:400];
        layer1[50][31:24] = buffer_data_3[415:408];
        layer1[50][39:32] = buffer_data_3[423:416];
        layer2[50][7:0] = buffer_data_2[391:384];
        layer2[50][15:8] = buffer_data_2[399:392];
        layer2[50][23:16] = buffer_data_2[407:400];
        layer2[50][31:24] = buffer_data_2[415:408];
        layer2[50][39:32] = buffer_data_2[423:416];
        layer3[50][7:0] = buffer_data_1[391:384];
        layer3[50][15:8] = buffer_data_1[399:392];
        layer3[50][23:16] = buffer_data_1[407:400];
        layer3[50][31:24] = buffer_data_1[415:408];
        layer3[50][39:32] = buffer_data_1[423:416];
        layer4[50][7:0] = buffer_data_0[391:384];
        layer4[50][15:8] = buffer_data_0[399:392];
        layer4[50][23:16] = buffer_data_0[407:400];
        layer4[50][31:24] = buffer_data_0[415:408];
        layer4[50][39:32] = buffer_data_0[423:416];
        layer0[51][7:0] = buffer_data_4[399:392];
        layer0[51][15:8] = buffer_data_4[407:400];
        layer0[51][23:16] = buffer_data_4[415:408];
        layer0[51][31:24] = buffer_data_4[423:416];
        layer0[51][39:32] = buffer_data_4[431:424];
        layer1[51][7:0] = buffer_data_3[399:392];
        layer1[51][15:8] = buffer_data_3[407:400];
        layer1[51][23:16] = buffer_data_3[415:408];
        layer1[51][31:24] = buffer_data_3[423:416];
        layer1[51][39:32] = buffer_data_3[431:424];
        layer2[51][7:0] = buffer_data_2[399:392];
        layer2[51][15:8] = buffer_data_2[407:400];
        layer2[51][23:16] = buffer_data_2[415:408];
        layer2[51][31:24] = buffer_data_2[423:416];
        layer2[51][39:32] = buffer_data_2[431:424];
        layer3[51][7:0] = buffer_data_1[399:392];
        layer3[51][15:8] = buffer_data_1[407:400];
        layer3[51][23:16] = buffer_data_1[415:408];
        layer3[51][31:24] = buffer_data_1[423:416];
        layer3[51][39:32] = buffer_data_1[431:424];
        layer4[51][7:0] = buffer_data_0[399:392];
        layer4[51][15:8] = buffer_data_0[407:400];
        layer4[51][23:16] = buffer_data_0[415:408];
        layer4[51][31:24] = buffer_data_0[423:416];
        layer4[51][39:32] = buffer_data_0[431:424];
        layer0[52][7:0] = buffer_data_4[407:400];
        layer0[52][15:8] = buffer_data_4[415:408];
        layer0[52][23:16] = buffer_data_4[423:416];
        layer0[52][31:24] = buffer_data_4[431:424];
        layer0[52][39:32] = buffer_data_4[439:432];
        layer1[52][7:0] = buffer_data_3[407:400];
        layer1[52][15:8] = buffer_data_3[415:408];
        layer1[52][23:16] = buffer_data_3[423:416];
        layer1[52][31:24] = buffer_data_3[431:424];
        layer1[52][39:32] = buffer_data_3[439:432];
        layer2[52][7:0] = buffer_data_2[407:400];
        layer2[52][15:8] = buffer_data_2[415:408];
        layer2[52][23:16] = buffer_data_2[423:416];
        layer2[52][31:24] = buffer_data_2[431:424];
        layer2[52][39:32] = buffer_data_2[439:432];
        layer3[52][7:0] = buffer_data_1[407:400];
        layer3[52][15:8] = buffer_data_1[415:408];
        layer3[52][23:16] = buffer_data_1[423:416];
        layer3[52][31:24] = buffer_data_1[431:424];
        layer3[52][39:32] = buffer_data_1[439:432];
        layer4[52][7:0] = buffer_data_0[407:400];
        layer4[52][15:8] = buffer_data_0[415:408];
        layer4[52][23:16] = buffer_data_0[423:416];
        layer4[52][31:24] = buffer_data_0[431:424];
        layer4[52][39:32] = buffer_data_0[439:432];
        layer0[53][7:0] = buffer_data_4[415:408];
        layer0[53][15:8] = buffer_data_4[423:416];
        layer0[53][23:16] = buffer_data_4[431:424];
        layer0[53][31:24] = buffer_data_4[439:432];
        layer0[53][39:32] = buffer_data_4[447:440];
        layer1[53][7:0] = buffer_data_3[415:408];
        layer1[53][15:8] = buffer_data_3[423:416];
        layer1[53][23:16] = buffer_data_3[431:424];
        layer1[53][31:24] = buffer_data_3[439:432];
        layer1[53][39:32] = buffer_data_3[447:440];
        layer2[53][7:0] = buffer_data_2[415:408];
        layer2[53][15:8] = buffer_data_2[423:416];
        layer2[53][23:16] = buffer_data_2[431:424];
        layer2[53][31:24] = buffer_data_2[439:432];
        layer2[53][39:32] = buffer_data_2[447:440];
        layer3[53][7:0] = buffer_data_1[415:408];
        layer3[53][15:8] = buffer_data_1[423:416];
        layer3[53][23:16] = buffer_data_1[431:424];
        layer3[53][31:24] = buffer_data_1[439:432];
        layer3[53][39:32] = buffer_data_1[447:440];
        layer4[53][7:0] = buffer_data_0[415:408];
        layer4[53][15:8] = buffer_data_0[423:416];
        layer4[53][23:16] = buffer_data_0[431:424];
        layer4[53][31:24] = buffer_data_0[439:432];
        layer4[53][39:32] = buffer_data_0[447:440];
        layer0[54][7:0] = buffer_data_4[423:416];
        layer0[54][15:8] = buffer_data_4[431:424];
        layer0[54][23:16] = buffer_data_4[439:432];
        layer0[54][31:24] = buffer_data_4[447:440];
        layer0[54][39:32] = buffer_data_4[455:448];
        layer1[54][7:0] = buffer_data_3[423:416];
        layer1[54][15:8] = buffer_data_3[431:424];
        layer1[54][23:16] = buffer_data_3[439:432];
        layer1[54][31:24] = buffer_data_3[447:440];
        layer1[54][39:32] = buffer_data_3[455:448];
        layer2[54][7:0] = buffer_data_2[423:416];
        layer2[54][15:8] = buffer_data_2[431:424];
        layer2[54][23:16] = buffer_data_2[439:432];
        layer2[54][31:24] = buffer_data_2[447:440];
        layer2[54][39:32] = buffer_data_2[455:448];
        layer3[54][7:0] = buffer_data_1[423:416];
        layer3[54][15:8] = buffer_data_1[431:424];
        layer3[54][23:16] = buffer_data_1[439:432];
        layer3[54][31:24] = buffer_data_1[447:440];
        layer3[54][39:32] = buffer_data_1[455:448];
        layer4[54][7:0] = buffer_data_0[423:416];
        layer4[54][15:8] = buffer_data_0[431:424];
        layer4[54][23:16] = buffer_data_0[439:432];
        layer4[54][31:24] = buffer_data_0[447:440];
        layer4[54][39:32] = buffer_data_0[455:448];
        layer0[55][7:0] = buffer_data_4[431:424];
        layer0[55][15:8] = buffer_data_4[439:432];
        layer0[55][23:16] = buffer_data_4[447:440];
        layer0[55][31:24] = buffer_data_4[455:448];
        layer0[55][39:32] = buffer_data_4[463:456];
        layer1[55][7:0] = buffer_data_3[431:424];
        layer1[55][15:8] = buffer_data_3[439:432];
        layer1[55][23:16] = buffer_data_3[447:440];
        layer1[55][31:24] = buffer_data_3[455:448];
        layer1[55][39:32] = buffer_data_3[463:456];
        layer2[55][7:0] = buffer_data_2[431:424];
        layer2[55][15:8] = buffer_data_2[439:432];
        layer2[55][23:16] = buffer_data_2[447:440];
        layer2[55][31:24] = buffer_data_2[455:448];
        layer2[55][39:32] = buffer_data_2[463:456];
        layer3[55][7:0] = buffer_data_1[431:424];
        layer3[55][15:8] = buffer_data_1[439:432];
        layer3[55][23:16] = buffer_data_1[447:440];
        layer3[55][31:24] = buffer_data_1[455:448];
        layer3[55][39:32] = buffer_data_1[463:456];
        layer4[55][7:0] = buffer_data_0[431:424];
        layer4[55][15:8] = buffer_data_0[439:432];
        layer4[55][23:16] = buffer_data_0[447:440];
        layer4[55][31:24] = buffer_data_0[455:448];
        layer4[55][39:32] = buffer_data_0[463:456];
        layer0[56][7:0] = buffer_data_4[439:432];
        layer0[56][15:8] = buffer_data_4[447:440];
        layer0[56][23:16] = buffer_data_4[455:448];
        layer0[56][31:24] = buffer_data_4[463:456];
        layer0[56][39:32] = buffer_data_4[471:464];
        layer1[56][7:0] = buffer_data_3[439:432];
        layer1[56][15:8] = buffer_data_3[447:440];
        layer1[56][23:16] = buffer_data_3[455:448];
        layer1[56][31:24] = buffer_data_3[463:456];
        layer1[56][39:32] = buffer_data_3[471:464];
        layer2[56][7:0] = buffer_data_2[439:432];
        layer2[56][15:8] = buffer_data_2[447:440];
        layer2[56][23:16] = buffer_data_2[455:448];
        layer2[56][31:24] = buffer_data_2[463:456];
        layer2[56][39:32] = buffer_data_2[471:464];
        layer3[56][7:0] = buffer_data_1[439:432];
        layer3[56][15:8] = buffer_data_1[447:440];
        layer3[56][23:16] = buffer_data_1[455:448];
        layer3[56][31:24] = buffer_data_1[463:456];
        layer3[56][39:32] = buffer_data_1[471:464];
        layer4[56][7:0] = buffer_data_0[439:432];
        layer4[56][15:8] = buffer_data_0[447:440];
        layer4[56][23:16] = buffer_data_0[455:448];
        layer4[56][31:24] = buffer_data_0[463:456];
        layer4[56][39:32] = buffer_data_0[471:464];
        layer0[57][7:0] = buffer_data_4[447:440];
        layer0[57][15:8] = buffer_data_4[455:448];
        layer0[57][23:16] = buffer_data_4[463:456];
        layer0[57][31:24] = buffer_data_4[471:464];
        layer0[57][39:32] = buffer_data_4[479:472];
        layer1[57][7:0] = buffer_data_3[447:440];
        layer1[57][15:8] = buffer_data_3[455:448];
        layer1[57][23:16] = buffer_data_3[463:456];
        layer1[57][31:24] = buffer_data_3[471:464];
        layer1[57][39:32] = buffer_data_3[479:472];
        layer2[57][7:0] = buffer_data_2[447:440];
        layer2[57][15:8] = buffer_data_2[455:448];
        layer2[57][23:16] = buffer_data_2[463:456];
        layer2[57][31:24] = buffer_data_2[471:464];
        layer2[57][39:32] = buffer_data_2[479:472];
        layer3[57][7:0] = buffer_data_1[447:440];
        layer3[57][15:8] = buffer_data_1[455:448];
        layer3[57][23:16] = buffer_data_1[463:456];
        layer3[57][31:24] = buffer_data_1[471:464];
        layer3[57][39:32] = buffer_data_1[479:472];
        layer4[57][7:0] = buffer_data_0[447:440];
        layer4[57][15:8] = buffer_data_0[455:448];
        layer4[57][23:16] = buffer_data_0[463:456];
        layer4[57][31:24] = buffer_data_0[471:464];
        layer4[57][39:32] = buffer_data_0[479:472];
        layer0[58][7:0] = buffer_data_4[455:448];
        layer0[58][15:8] = buffer_data_4[463:456];
        layer0[58][23:16] = buffer_data_4[471:464];
        layer0[58][31:24] = buffer_data_4[479:472];
        layer0[58][39:32] = buffer_data_4[487:480];
        layer1[58][7:0] = buffer_data_3[455:448];
        layer1[58][15:8] = buffer_data_3[463:456];
        layer1[58][23:16] = buffer_data_3[471:464];
        layer1[58][31:24] = buffer_data_3[479:472];
        layer1[58][39:32] = buffer_data_3[487:480];
        layer2[58][7:0] = buffer_data_2[455:448];
        layer2[58][15:8] = buffer_data_2[463:456];
        layer2[58][23:16] = buffer_data_2[471:464];
        layer2[58][31:24] = buffer_data_2[479:472];
        layer2[58][39:32] = buffer_data_2[487:480];
        layer3[58][7:0] = buffer_data_1[455:448];
        layer3[58][15:8] = buffer_data_1[463:456];
        layer3[58][23:16] = buffer_data_1[471:464];
        layer3[58][31:24] = buffer_data_1[479:472];
        layer3[58][39:32] = buffer_data_1[487:480];
        layer4[58][7:0] = buffer_data_0[455:448];
        layer4[58][15:8] = buffer_data_0[463:456];
        layer4[58][23:16] = buffer_data_0[471:464];
        layer4[58][31:24] = buffer_data_0[479:472];
        layer4[58][39:32] = buffer_data_0[487:480];
        layer0[59][7:0] = buffer_data_4[463:456];
        layer0[59][15:8] = buffer_data_4[471:464];
        layer0[59][23:16] = buffer_data_4[479:472];
        layer0[59][31:24] = buffer_data_4[487:480];
        layer0[59][39:32] = buffer_data_4[495:488];
        layer1[59][7:0] = buffer_data_3[463:456];
        layer1[59][15:8] = buffer_data_3[471:464];
        layer1[59][23:16] = buffer_data_3[479:472];
        layer1[59][31:24] = buffer_data_3[487:480];
        layer1[59][39:32] = buffer_data_3[495:488];
        layer2[59][7:0] = buffer_data_2[463:456];
        layer2[59][15:8] = buffer_data_2[471:464];
        layer2[59][23:16] = buffer_data_2[479:472];
        layer2[59][31:24] = buffer_data_2[487:480];
        layer2[59][39:32] = buffer_data_2[495:488];
        layer3[59][7:0] = buffer_data_1[463:456];
        layer3[59][15:8] = buffer_data_1[471:464];
        layer3[59][23:16] = buffer_data_1[479:472];
        layer3[59][31:24] = buffer_data_1[487:480];
        layer3[59][39:32] = buffer_data_1[495:488];
        layer4[59][7:0] = buffer_data_0[463:456];
        layer4[59][15:8] = buffer_data_0[471:464];
        layer4[59][23:16] = buffer_data_0[479:472];
        layer4[59][31:24] = buffer_data_0[487:480];
        layer4[59][39:32] = buffer_data_0[495:488];
        layer0[60][7:0] = buffer_data_4[471:464];
        layer0[60][15:8] = buffer_data_4[479:472];
        layer0[60][23:16] = buffer_data_4[487:480];
        layer0[60][31:24] = buffer_data_4[495:488];
        layer0[60][39:32] = buffer_data_4[503:496];
        layer1[60][7:0] = buffer_data_3[471:464];
        layer1[60][15:8] = buffer_data_3[479:472];
        layer1[60][23:16] = buffer_data_3[487:480];
        layer1[60][31:24] = buffer_data_3[495:488];
        layer1[60][39:32] = buffer_data_3[503:496];
        layer2[60][7:0] = buffer_data_2[471:464];
        layer2[60][15:8] = buffer_data_2[479:472];
        layer2[60][23:16] = buffer_data_2[487:480];
        layer2[60][31:24] = buffer_data_2[495:488];
        layer2[60][39:32] = buffer_data_2[503:496];
        layer3[60][7:0] = buffer_data_1[471:464];
        layer3[60][15:8] = buffer_data_1[479:472];
        layer3[60][23:16] = buffer_data_1[487:480];
        layer3[60][31:24] = buffer_data_1[495:488];
        layer3[60][39:32] = buffer_data_1[503:496];
        layer4[60][7:0] = buffer_data_0[471:464];
        layer4[60][15:8] = buffer_data_0[479:472];
        layer4[60][23:16] = buffer_data_0[487:480];
        layer4[60][31:24] = buffer_data_0[495:488];
        layer4[60][39:32] = buffer_data_0[503:496];
        layer0[61][7:0] = buffer_data_4[479:472];
        layer0[61][15:8] = buffer_data_4[487:480];
        layer0[61][23:16] = buffer_data_4[495:488];
        layer0[61][31:24] = buffer_data_4[503:496];
        layer0[61][39:32] = buffer_data_4[511:504];
        layer1[61][7:0] = buffer_data_3[479:472];
        layer1[61][15:8] = buffer_data_3[487:480];
        layer1[61][23:16] = buffer_data_3[495:488];
        layer1[61][31:24] = buffer_data_3[503:496];
        layer1[61][39:32] = buffer_data_3[511:504];
        layer2[61][7:0] = buffer_data_2[479:472];
        layer2[61][15:8] = buffer_data_2[487:480];
        layer2[61][23:16] = buffer_data_2[495:488];
        layer2[61][31:24] = buffer_data_2[503:496];
        layer2[61][39:32] = buffer_data_2[511:504];
        layer3[61][7:0] = buffer_data_1[479:472];
        layer3[61][15:8] = buffer_data_1[487:480];
        layer3[61][23:16] = buffer_data_1[495:488];
        layer3[61][31:24] = buffer_data_1[503:496];
        layer3[61][39:32] = buffer_data_1[511:504];
        layer4[61][7:0] = buffer_data_0[479:472];
        layer4[61][15:8] = buffer_data_0[487:480];
        layer4[61][23:16] = buffer_data_0[495:488];
        layer4[61][31:24] = buffer_data_0[503:496];
        layer4[61][39:32] = buffer_data_0[511:504];
        layer0[62][7:0] = buffer_data_4[487:480];
        layer0[62][15:8] = buffer_data_4[495:488];
        layer0[62][23:16] = buffer_data_4[503:496];
        layer0[62][31:24] = buffer_data_4[511:504];
        layer0[62][39:32] = buffer_data_4[519:512];
        layer1[62][7:0] = buffer_data_3[487:480];
        layer1[62][15:8] = buffer_data_3[495:488];
        layer1[62][23:16] = buffer_data_3[503:496];
        layer1[62][31:24] = buffer_data_3[511:504];
        layer1[62][39:32] = buffer_data_3[519:512];
        layer2[62][7:0] = buffer_data_2[487:480];
        layer2[62][15:8] = buffer_data_2[495:488];
        layer2[62][23:16] = buffer_data_2[503:496];
        layer2[62][31:24] = buffer_data_2[511:504];
        layer2[62][39:32] = buffer_data_2[519:512];
        layer3[62][7:0] = buffer_data_1[487:480];
        layer3[62][15:8] = buffer_data_1[495:488];
        layer3[62][23:16] = buffer_data_1[503:496];
        layer3[62][31:24] = buffer_data_1[511:504];
        layer3[62][39:32] = buffer_data_1[519:512];
        layer4[62][7:0] = buffer_data_0[487:480];
        layer4[62][15:8] = buffer_data_0[495:488];
        layer4[62][23:16] = buffer_data_0[503:496];
        layer4[62][31:24] = buffer_data_0[511:504];
        layer4[62][39:32] = buffer_data_0[519:512];
        layer0[63][7:0] = buffer_data_4[495:488];
        layer0[63][15:8] = buffer_data_4[503:496];
        layer0[63][23:16] = buffer_data_4[511:504];
        layer0[63][31:24] = buffer_data_4[519:512];
        layer0[63][39:32] = buffer_data_4[527:520];
        layer1[63][7:0] = buffer_data_3[495:488];
        layer1[63][15:8] = buffer_data_3[503:496];
        layer1[63][23:16] = buffer_data_3[511:504];
        layer1[63][31:24] = buffer_data_3[519:512];
        layer1[63][39:32] = buffer_data_3[527:520];
        layer2[63][7:0] = buffer_data_2[495:488];
        layer2[63][15:8] = buffer_data_2[503:496];
        layer2[63][23:16] = buffer_data_2[511:504];
        layer2[63][31:24] = buffer_data_2[519:512];
        layer2[63][39:32] = buffer_data_2[527:520];
        layer3[63][7:0] = buffer_data_1[495:488];
        layer3[63][15:8] = buffer_data_1[503:496];
        layer3[63][23:16] = buffer_data_1[511:504];
        layer3[63][31:24] = buffer_data_1[519:512];
        layer3[63][39:32] = buffer_data_1[527:520];
        layer4[63][7:0] = buffer_data_0[495:488];
        layer4[63][15:8] = buffer_data_0[503:496];
        layer4[63][23:16] = buffer_data_0[511:504];
        layer4[63][31:24] = buffer_data_0[519:512];
        layer4[63][39:32] = buffer_data_0[527:520];
    end
    ST_GAUSSIAN_1: begin
        layer0[0][7:0] = buffer_data_4[503:496];
        layer0[0][15:8] = buffer_data_4[511:504];
        layer0[0][23:16] = buffer_data_4[519:512];
        layer0[0][31:24] = buffer_data_4[527:520];
        layer0[0][39:32] = buffer_data_4[535:528];
        layer1[0][7:0] = buffer_data_3[503:496];
        layer1[0][15:8] = buffer_data_3[511:504];
        layer1[0][23:16] = buffer_data_3[519:512];
        layer1[0][31:24] = buffer_data_3[527:520];
        layer1[0][39:32] = buffer_data_3[535:528];
        layer2[0][7:0] = buffer_data_2[503:496];
        layer2[0][15:8] = buffer_data_2[511:504];
        layer2[0][23:16] = buffer_data_2[519:512];
        layer2[0][31:24] = buffer_data_2[527:520];
        layer2[0][39:32] = buffer_data_2[535:528];
        layer3[0][7:0] = buffer_data_1[503:496];
        layer3[0][15:8] = buffer_data_1[511:504];
        layer3[0][23:16] = buffer_data_1[519:512];
        layer3[0][31:24] = buffer_data_1[527:520];
        layer3[0][39:32] = buffer_data_1[535:528];
        layer4[0][7:0] = buffer_data_0[503:496];
        layer4[0][15:8] = buffer_data_0[511:504];
        layer4[0][23:16] = buffer_data_0[519:512];
        layer4[0][31:24] = buffer_data_0[527:520];
        layer4[0][39:32] = buffer_data_0[535:528];
        layer0[1][7:0] = buffer_data_4[511:504];
        layer0[1][15:8] = buffer_data_4[519:512];
        layer0[1][23:16] = buffer_data_4[527:520];
        layer0[1][31:24] = buffer_data_4[535:528];
        layer0[1][39:32] = buffer_data_4[543:536];
        layer1[1][7:0] = buffer_data_3[511:504];
        layer1[1][15:8] = buffer_data_3[519:512];
        layer1[1][23:16] = buffer_data_3[527:520];
        layer1[1][31:24] = buffer_data_3[535:528];
        layer1[1][39:32] = buffer_data_3[543:536];
        layer2[1][7:0] = buffer_data_2[511:504];
        layer2[1][15:8] = buffer_data_2[519:512];
        layer2[1][23:16] = buffer_data_2[527:520];
        layer2[1][31:24] = buffer_data_2[535:528];
        layer2[1][39:32] = buffer_data_2[543:536];
        layer3[1][7:0] = buffer_data_1[511:504];
        layer3[1][15:8] = buffer_data_1[519:512];
        layer3[1][23:16] = buffer_data_1[527:520];
        layer3[1][31:24] = buffer_data_1[535:528];
        layer3[1][39:32] = buffer_data_1[543:536];
        layer4[1][7:0] = buffer_data_0[511:504];
        layer4[1][15:8] = buffer_data_0[519:512];
        layer4[1][23:16] = buffer_data_0[527:520];
        layer4[1][31:24] = buffer_data_0[535:528];
        layer4[1][39:32] = buffer_data_0[543:536];
        layer0[2][7:0] = buffer_data_4[519:512];
        layer0[2][15:8] = buffer_data_4[527:520];
        layer0[2][23:16] = buffer_data_4[535:528];
        layer0[2][31:24] = buffer_data_4[543:536];
        layer0[2][39:32] = buffer_data_4[551:544];
        layer1[2][7:0] = buffer_data_3[519:512];
        layer1[2][15:8] = buffer_data_3[527:520];
        layer1[2][23:16] = buffer_data_3[535:528];
        layer1[2][31:24] = buffer_data_3[543:536];
        layer1[2][39:32] = buffer_data_3[551:544];
        layer2[2][7:0] = buffer_data_2[519:512];
        layer2[2][15:8] = buffer_data_2[527:520];
        layer2[2][23:16] = buffer_data_2[535:528];
        layer2[2][31:24] = buffer_data_2[543:536];
        layer2[2][39:32] = buffer_data_2[551:544];
        layer3[2][7:0] = buffer_data_1[519:512];
        layer3[2][15:8] = buffer_data_1[527:520];
        layer3[2][23:16] = buffer_data_1[535:528];
        layer3[2][31:24] = buffer_data_1[543:536];
        layer3[2][39:32] = buffer_data_1[551:544];
        layer4[2][7:0] = buffer_data_0[519:512];
        layer4[2][15:8] = buffer_data_0[527:520];
        layer4[2][23:16] = buffer_data_0[535:528];
        layer4[2][31:24] = buffer_data_0[543:536];
        layer4[2][39:32] = buffer_data_0[551:544];
        layer0[3][7:0] = buffer_data_4[527:520];
        layer0[3][15:8] = buffer_data_4[535:528];
        layer0[3][23:16] = buffer_data_4[543:536];
        layer0[3][31:24] = buffer_data_4[551:544];
        layer0[3][39:32] = buffer_data_4[559:552];
        layer1[3][7:0] = buffer_data_3[527:520];
        layer1[3][15:8] = buffer_data_3[535:528];
        layer1[3][23:16] = buffer_data_3[543:536];
        layer1[3][31:24] = buffer_data_3[551:544];
        layer1[3][39:32] = buffer_data_3[559:552];
        layer2[3][7:0] = buffer_data_2[527:520];
        layer2[3][15:8] = buffer_data_2[535:528];
        layer2[3][23:16] = buffer_data_2[543:536];
        layer2[3][31:24] = buffer_data_2[551:544];
        layer2[3][39:32] = buffer_data_2[559:552];
        layer3[3][7:0] = buffer_data_1[527:520];
        layer3[3][15:8] = buffer_data_1[535:528];
        layer3[3][23:16] = buffer_data_1[543:536];
        layer3[3][31:24] = buffer_data_1[551:544];
        layer3[3][39:32] = buffer_data_1[559:552];
        layer4[3][7:0] = buffer_data_0[527:520];
        layer4[3][15:8] = buffer_data_0[535:528];
        layer4[3][23:16] = buffer_data_0[543:536];
        layer4[3][31:24] = buffer_data_0[551:544];
        layer4[3][39:32] = buffer_data_0[559:552];
        layer0[4][7:0] = buffer_data_4[535:528];
        layer0[4][15:8] = buffer_data_4[543:536];
        layer0[4][23:16] = buffer_data_4[551:544];
        layer0[4][31:24] = buffer_data_4[559:552];
        layer0[4][39:32] = buffer_data_4[567:560];
        layer1[4][7:0] = buffer_data_3[535:528];
        layer1[4][15:8] = buffer_data_3[543:536];
        layer1[4][23:16] = buffer_data_3[551:544];
        layer1[4][31:24] = buffer_data_3[559:552];
        layer1[4][39:32] = buffer_data_3[567:560];
        layer2[4][7:0] = buffer_data_2[535:528];
        layer2[4][15:8] = buffer_data_2[543:536];
        layer2[4][23:16] = buffer_data_2[551:544];
        layer2[4][31:24] = buffer_data_2[559:552];
        layer2[4][39:32] = buffer_data_2[567:560];
        layer3[4][7:0] = buffer_data_1[535:528];
        layer3[4][15:8] = buffer_data_1[543:536];
        layer3[4][23:16] = buffer_data_1[551:544];
        layer3[4][31:24] = buffer_data_1[559:552];
        layer3[4][39:32] = buffer_data_1[567:560];
        layer4[4][7:0] = buffer_data_0[535:528];
        layer4[4][15:8] = buffer_data_0[543:536];
        layer4[4][23:16] = buffer_data_0[551:544];
        layer4[4][31:24] = buffer_data_0[559:552];
        layer4[4][39:32] = buffer_data_0[567:560];
        layer0[5][7:0] = buffer_data_4[543:536];
        layer0[5][15:8] = buffer_data_4[551:544];
        layer0[5][23:16] = buffer_data_4[559:552];
        layer0[5][31:24] = buffer_data_4[567:560];
        layer0[5][39:32] = buffer_data_4[575:568];
        layer1[5][7:0] = buffer_data_3[543:536];
        layer1[5][15:8] = buffer_data_3[551:544];
        layer1[5][23:16] = buffer_data_3[559:552];
        layer1[5][31:24] = buffer_data_3[567:560];
        layer1[5][39:32] = buffer_data_3[575:568];
        layer2[5][7:0] = buffer_data_2[543:536];
        layer2[5][15:8] = buffer_data_2[551:544];
        layer2[5][23:16] = buffer_data_2[559:552];
        layer2[5][31:24] = buffer_data_2[567:560];
        layer2[5][39:32] = buffer_data_2[575:568];
        layer3[5][7:0] = buffer_data_1[543:536];
        layer3[5][15:8] = buffer_data_1[551:544];
        layer3[5][23:16] = buffer_data_1[559:552];
        layer3[5][31:24] = buffer_data_1[567:560];
        layer3[5][39:32] = buffer_data_1[575:568];
        layer4[5][7:0] = buffer_data_0[543:536];
        layer4[5][15:8] = buffer_data_0[551:544];
        layer4[5][23:16] = buffer_data_0[559:552];
        layer4[5][31:24] = buffer_data_0[567:560];
        layer4[5][39:32] = buffer_data_0[575:568];
        layer0[6][7:0] = buffer_data_4[551:544];
        layer0[6][15:8] = buffer_data_4[559:552];
        layer0[6][23:16] = buffer_data_4[567:560];
        layer0[6][31:24] = buffer_data_4[575:568];
        layer0[6][39:32] = buffer_data_4[583:576];
        layer1[6][7:0] = buffer_data_3[551:544];
        layer1[6][15:8] = buffer_data_3[559:552];
        layer1[6][23:16] = buffer_data_3[567:560];
        layer1[6][31:24] = buffer_data_3[575:568];
        layer1[6][39:32] = buffer_data_3[583:576];
        layer2[6][7:0] = buffer_data_2[551:544];
        layer2[6][15:8] = buffer_data_2[559:552];
        layer2[6][23:16] = buffer_data_2[567:560];
        layer2[6][31:24] = buffer_data_2[575:568];
        layer2[6][39:32] = buffer_data_2[583:576];
        layer3[6][7:0] = buffer_data_1[551:544];
        layer3[6][15:8] = buffer_data_1[559:552];
        layer3[6][23:16] = buffer_data_1[567:560];
        layer3[6][31:24] = buffer_data_1[575:568];
        layer3[6][39:32] = buffer_data_1[583:576];
        layer4[6][7:0] = buffer_data_0[551:544];
        layer4[6][15:8] = buffer_data_0[559:552];
        layer4[6][23:16] = buffer_data_0[567:560];
        layer4[6][31:24] = buffer_data_0[575:568];
        layer4[6][39:32] = buffer_data_0[583:576];
        layer0[7][7:0] = buffer_data_4[559:552];
        layer0[7][15:8] = buffer_data_4[567:560];
        layer0[7][23:16] = buffer_data_4[575:568];
        layer0[7][31:24] = buffer_data_4[583:576];
        layer0[7][39:32] = buffer_data_4[591:584];
        layer1[7][7:0] = buffer_data_3[559:552];
        layer1[7][15:8] = buffer_data_3[567:560];
        layer1[7][23:16] = buffer_data_3[575:568];
        layer1[7][31:24] = buffer_data_3[583:576];
        layer1[7][39:32] = buffer_data_3[591:584];
        layer2[7][7:0] = buffer_data_2[559:552];
        layer2[7][15:8] = buffer_data_2[567:560];
        layer2[7][23:16] = buffer_data_2[575:568];
        layer2[7][31:24] = buffer_data_2[583:576];
        layer2[7][39:32] = buffer_data_2[591:584];
        layer3[7][7:0] = buffer_data_1[559:552];
        layer3[7][15:8] = buffer_data_1[567:560];
        layer3[7][23:16] = buffer_data_1[575:568];
        layer3[7][31:24] = buffer_data_1[583:576];
        layer3[7][39:32] = buffer_data_1[591:584];
        layer4[7][7:0] = buffer_data_0[559:552];
        layer4[7][15:8] = buffer_data_0[567:560];
        layer4[7][23:16] = buffer_data_0[575:568];
        layer4[7][31:24] = buffer_data_0[583:576];
        layer4[7][39:32] = buffer_data_0[591:584];
        layer0[8][7:0] = buffer_data_4[567:560];
        layer0[8][15:8] = buffer_data_4[575:568];
        layer0[8][23:16] = buffer_data_4[583:576];
        layer0[8][31:24] = buffer_data_4[591:584];
        layer0[8][39:32] = buffer_data_4[599:592];
        layer1[8][7:0] = buffer_data_3[567:560];
        layer1[8][15:8] = buffer_data_3[575:568];
        layer1[8][23:16] = buffer_data_3[583:576];
        layer1[8][31:24] = buffer_data_3[591:584];
        layer1[8][39:32] = buffer_data_3[599:592];
        layer2[8][7:0] = buffer_data_2[567:560];
        layer2[8][15:8] = buffer_data_2[575:568];
        layer2[8][23:16] = buffer_data_2[583:576];
        layer2[8][31:24] = buffer_data_2[591:584];
        layer2[8][39:32] = buffer_data_2[599:592];
        layer3[8][7:0] = buffer_data_1[567:560];
        layer3[8][15:8] = buffer_data_1[575:568];
        layer3[8][23:16] = buffer_data_1[583:576];
        layer3[8][31:24] = buffer_data_1[591:584];
        layer3[8][39:32] = buffer_data_1[599:592];
        layer4[8][7:0] = buffer_data_0[567:560];
        layer4[8][15:8] = buffer_data_0[575:568];
        layer4[8][23:16] = buffer_data_0[583:576];
        layer4[8][31:24] = buffer_data_0[591:584];
        layer4[8][39:32] = buffer_data_0[599:592];
        layer0[9][7:0] = buffer_data_4[575:568];
        layer0[9][15:8] = buffer_data_4[583:576];
        layer0[9][23:16] = buffer_data_4[591:584];
        layer0[9][31:24] = buffer_data_4[599:592];
        layer0[9][39:32] = buffer_data_4[607:600];
        layer1[9][7:0] = buffer_data_3[575:568];
        layer1[9][15:8] = buffer_data_3[583:576];
        layer1[9][23:16] = buffer_data_3[591:584];
        layer1[9][31:24] = buffer_data_3[599:592];
        layer1[9][39:32] = buffer_data_3[607:600];
        layer2[9][7:0] = buffer_data_2[575:568];
        layer2[9][15:8] = buffer_data_2[583:576];
        layer2[9][23:16] = buffer_data_2[591:584];
        layer2[9][31:24] = buffer_data_2[599:592];
        layer2[9][39:32] = buffer_data_2[607:600];
        layer3[9][7:0] = buffer_data_1[575:568];
        layer3[9][15:8] = buffer_data_1[583:576];
        layer3[9][23:16] = buffer_data_1[591:584];
        layer3[9][31:24] = buffer_data_1[599:592];
        layer3[9][39:32] = buffer_data_1[607:600];
        layer4[9][7:0] = buffer_data_0[575:568];
        layer4[9][15:8] = buffer_data_0[583:576];
        layer4[9][23:16] = buffer_data_0[591:584];
        layer4[9][31:24] = buffer_data_0[599:592];
        layer4[9][39:32] = buffer_data_0[607:600];
        layer0[10][7:0] = buffer_data_4[583:576];
        layer0[10][15:8] = buffer_data_4[591:584];
        layer0[10][23:16] = buffer_data_4[599:592];
        layer0[10][31:24] = buffer_data_4[607:600];
        layer0[10][39:32] = buffer_data_4[615:608];
        layer1[10][7:0] = buffer_data_3[583:576];
        layer1[10][15:8] = buffer_data_3[591:584];
        layer1[10][23:16] = buffer_data_3[599:592];
        layer1[10][31:24] = buffer_data_3[607:600];
        layer1[10][39:32] = buffer_data_3[615:608];
        layer2[10][7:0] = buffer_data_2[583:576];
        layer2[10][15:8] = buffer_data_2[591:584];
        layer2[10][23:16] = buffer_data_2[599:592];
        layer2[10][31:24] = buffer_data_2[607:600];
        layer2[10][39:32] = buffer_data_2[615:608];
        layer3[10][7:0] = buffer_data_1[583:576];
        layer3[10][15:8] = buffer_data_1[591:584];
        layer3[10][23:16] = buffer_data_1[599:592];
        layer3[10][31:24] = buffer_data_1[607:600];
        layer3[10][39:32] = buffer_data_1[615:608];
        layer4[10][7:0] = buffer_data_0[583:576];
        layer4[10][15:8] = buffer_data_0[591:584];
        layer4[10][23:16] = buffer_data_0[599:592];
        layer4[10][31:24] = buffer_data_0[607:600];
        layer4[10][39:32] = buffer_data_0[615:608];
        layer0[11][7:0] = buffer_data_4[591:584];
        layer0[11][15:8] = buffer_data_4[599:592];
        layer0[11][23:16] = buffer_data_4[607:600];
        layer0[11][31:24] = buffer_data_4[615:608];
        layer0[11][39:32] = buffer_data_4[623:616];
        layer1[11][7:0] = buffer_data_3[591:584];
        layer1[11][15:8] = buffer_data_3[599:592];
        layer1[11][23:16] = buffer_data_3[607:600];
        layer1[11][31:24] = buffer_data_3[615:608];
        layer1[11][39:32] = buffer_data_3[623:616];
        layer2[11][7:0] = buffer_data_2[591:584];
        layer2[11][15:8] = buffer_data_2[599:592];
        layer2[11][23:16] = buffer_data_2[607:600];
        layer2[11][31:24] = buffer_data_2[615:608];
        layer2[11][39:32] = buffer_data_2[623:616];
        layer3[11][7:0] = buffer_data_1[591:584];
        layer3[11][15:8] = buffer_data_1[599:592];
        layer3[11][23:16] = buffer_data_1[607:600];
        layer3[11][31:24] = buffer_data_1[615:608];
        layer3[11][39:32] = buffer_data_1[623:616];
        layer4[11][7:0] = buffer_data_0[591:584];
        layer4[11][15:8] = buffer_data_0[599:592];
        layer4[11][23:16] = buffer_data_0[607:600];
        layer4[11][31:24] = buffer_data_0[615:608];
        layer4[11][39:32] = buffer_data_0[623:616];
        layer0[12][7:0] = buffer_data_4[599:592];
        layer0[12][15:8] = buffer_data_4[607:600];
        layer0[12][23:16] = buffer_data_4[615:608];
        layer0[12][31:24] = buffer_data_4[623:616];
        layer0[12][39:32] = buffer_data_4[631:624];
        layer1[12][7:0] = buffer_data_3[599:592];
        layer1[12][15:8] = buffer_data_3[607:600];
        layer1[12][23:16] = buffer_data_3[615:608];
        layer1[12][31:24] = buffer_data_3[623:616];
        layer1[12][39:32] = buffer_data_3[631:624];
        layer2[12][7:0] = buffer_data_2[599:592];
        layer2[12][15:8] = buffer_data_2[607:600];
        layer2[12][23:16] = buffer_data_2[615:608];
        layer2[12][31:24] = buffer_data_2[623:616];
        layer2[12][39:32] = buffer_data_2[631:624];
        layer3[12][7:0] = buffer_data_1[599:592];
        layer3[12][15:8] = buffer_data_1[607:600];
        layer3[12][23:16] = buffer_data_1[615:608];
        layer3[12][31:24] = buffer_data_1[623:616];
        layer3[12][39:32] = buffer_data_1[631:624];
        layer4[12][7:0] = buffer_data_0[599:592];
        layer4[12][15:8] = buffer_data_0[607:600];
        layer4[12][23:16] = buffer_data_0[615:608];
        layer4[12][31:24] = buffer_data_0[623:616];
        layer4[12][39:32] = buffer_data_0[631:624];
        layer0[13][7:0] = buffer_data_4[607:600];
        layer0[13][15:8] = buffer_data_4[615:608];
        layer0[13][23:16] = buffer_data_4[623:616];
        layer0[13][31:24] = buffer_data_4[631:624];
        layer0[13][39:32] = buffer_data_4[639:632];
        layer1[13][7:0] = buffer_data_3[607:600];
        layer1[13][15:8] = buffer_data_3[615:608];
        layer1[13][23:16] = buffer_data_3[623:616];
        layer1[13][31:24] = buffer_data_3[631:624];
        layer1[13][39:32] = buffer_data_3[639:632];
        layer2[13][7:0] = buffer_data_2[607:600];
        layer2[13][15:8] = buffer_data_2[615:608];
        layer2[13][23:16] = buffer_data_2[623:616];
        layer2[13][31:24] = buffer_data_2[631:624];
        layer2[13][39:32] = buffer_data_2[639:632];
        layer3[13][7:0] = buffer_data_1[607:600];
        layer3[13][15:8] = buffer_data_1[615:608];
        layer3[13][23:16] = buffer_data_1[623:616];
        layer3[13][31:24] = buffer_data_1[631:624];
        layer3[13][39:32] = buffer_data_1[639:632];
        layer4[13][7:0] = buffer_data_0[607:600];
        layer4[13][15:8] = buffer_data_0[615:608];
        layer4[13][23:16] = buffer_data_0[623:616];
        layer4[13][31:24] = buffer_data_0[631:624];
        layer4[13][39:32] = buffer_data_0[639:632];
        layer0[14][7:0] = buffer_data_4[615:608];
        layer0[14][15:8] = buffer_data_4[623:616];
        layer0[14][23:16] = buffer_data_4[631:624];
        layer0[14][31:24] = buffer_data_4[639:632];
        layer0[14][39:32] = buffer_data_4[647:640];
        layer1[14][7:0] = buffer_data_3[615:608];
        layer1[14][15:8] = buffer_data_3[623:616];
        layer1[14][23:16] = buffer_data_3[631:624];
        layer1[14][31:24] = buffer_data_3[639:632];
        layer1[14][39:32] = buffer_data_3[647:640];
        layer2[14][7:0] = buffer_data_2[615:608];
        layer2[14][15:8] = buffer_data_2[623:616];
        layer2[14][23:16] = buffer_data_2[631:624];
        layer2[14][31:24] = buffer_data_2[639:632];
        layer2[14][39:32] = buffer_data_2[647:640];
        layer3[14][7:0] = buffer_data_1[615:608];
        layer3[14][15:8] = buffer_data_1[623:616];
        layer3[14][23:16] = buffer_data_1[631:624];
        layer3[14][31:24] = buffer_data_1[639:632];
        layer3[14][39:32] = buffer_data_1[647:640];
        layer4[14][7:0] = buffer_data_0[615:608];
        layer4[14][15:8] = buffer_data_0[623:616];
        layer4[14][23:16] = buffer_data_0[631:624];
        layer4[14][31:24] = buffer_data_0[639:632];
        layer4[14][39:32] = buffer_data_0[647:640];
        layer0[15][7:0] = buffer_data_4[623:616];
        layer0[15][15:8] = buffer_data_4[631:624];
        layer0[15][23:16] = buffer_data_4[639:632];
        layer0[15][31:24] = buffer_data_4[647:640];
        layer0[15][39:32] = buffer_data_4[655:648];
        layer1[15][7:0] = buffer_data_3[623:616];
        layer1[15][15:8] = buffer_data_3[631:624];
        layer1[15][23:16] = buffer_data_3[639:632];
        layer1[15][31:24] = buffer_data_3[647:640];
        layer1[15][39:32] = buffer_data_3[655:648];
        layer2[15][7:0] = buffer_data_2[623:616];
        layer2[15][15:8] = buffer_data_2[631:624];
        layer2[15][23:16] = buffer_data_2[639:632];
        layer2[15][31:24] = buffer_data_2[647:640];
        layer2[15][39:32] = buffer_data_2[655:648];
        layer3[15][7:0] = buffer_data_1[623:616];
        layer3[15][15:8] = buffer_data_1[631:624];
        layer3[15][23:16] = buffer_data_1[639:632];
        layer3[15][31:24] = buffer_data_1[647:640];
        layer3[15][39:32] = buffer_data_1[655:648];
        layer4[15][7:0] = buffer_data_0[623:616];
        layer4[15][15:8] = buffer_data_0[631:624];
        layer4[15][23:16] = buffer_data_0[639:632];
        layer4[15][31:24] = buffer_data_0[647:640];
        layer4[15][39:32] = buffer_data_0[655:648];
        layer0[16][7:0] = buffer_data_4[631:624];
        layer0[16][15:8] = buffer_data_4[639:632];
        layer0[16][23:16] = buffer_data_4[647:640];
        layer0[16][31:24] = buffer_data_4[655:648];
        layer0[16][39:32] = buffer_data_4[663:656];
        layer1[16][7:0] = buffer_data_3[631:624];
        layer1[16][15:8] = buffer_data_3[639:632];
        layer1[16][23:16] = buffer_data_3[647:640];
        layer1[16][31:24] = buffer_data_3[655:648];
        layer1[16][39:32] = buffer_data_3[663:656];
        layer2[16][7:0] = buffer_data_2[631:624];
        layer2[16][15:8] = buffer_data_2[639:632];
        layer2[16][23:16] = buffer_data_2[647:640];
        layer2[16][31:24] = buffer_data_2[655:648];
        layer2[16][39:32] = buffer_data_2[663:656];
        layer3[16][7:0] = buffer_data_1[631:624];
        layer3[16][15:8] = buffer_data_1[639:632];
        layer3[16][23:16] = buffer_data_1[647:640];
        layer3[16][31:24] = buffer_data_1[655:648];
        layer3[16][39:32] = buffer_data_1[663:656];
        layer4[16][7:0] = buffer_data_0[631:624];
        layer4[16][15:8] = buffer_data_0[639:632];
        layer4[16][23:16] = buffer_data_0[647:640];
        layer4[16][31:24] = buffer_data_0[655:648];
        layer4[16][39:32] = buffer_data_0[663:656];
        layer0[17][7:0] = buffer_data_4[639:632];
        layer0[17][15:8] = buffer_data_4[647:640];
        layer0[17][23:16] = buffer_data_4[655:648];
        layer0[17][31:24] = buffer_data_4[663:656];
        layer0[17][39:32] = buffer_data_4[671:664];
        layer1[17][7:0] = buffer_data_3[639:632];
        layer1[17][15:8] = buffer_data_3[647:640];
        layer1[17][23:16] = buffer_data_3[655:648];
        layer1[17][31:24] = buffer_data_3[663:656];
        layer1[17][39:32] = buffer_data_3[671:664];
        layer2[17][7:0] = buffer_data_2[639:632];
        layer2[17][15:8] = buffer_data_2[647:640];
        layer2[17][23:16] = buffer_data_2[655:648];
        layer2[17][31:24] = buffer_data_2[663:656];
        layer2[17][39:32] = buffer_data_2[671:664];
        layer3[17][7:0] = buffer_data_1[639:632];
        layer3[17][15:8] = buffer_data_1[647:640];
        layer3[17][23:16] = buffer_data_1[655:648];
        layer3[17][31:24] = buffer_data_1[663:656];
        layer3[17][39:32] = buffer_data_1[671:664];
        layer4[17][7:0] = buffer_data_0[639:632];
        layer4[17][15:8] = buffer_data_0[647:640];
        layer4[17][23:16] = buffer_data_0[655:648];
        layer4[17][31:24] = buffer_data_0[663:656];
        layer4[17][39:32] = buffer_data_0[671:664];
        layer0[18][7:0] = buffer_data_4[647:640];
        layer0[18][15:8] = buffer_data_4[655:648];
        layer0[18][23:16] = buffer_data_4[663:656];
        layer0[18][31:24] = buffer_data_4[671:664];
        layer0[18][39:32] = buffer_data_4[679:672];
        layer1[18][7:0] = buffer_data_3[647:640];
        layer1[18][15:8] = buffer_data_3[655:648];
        layer1[18][23:16] = buffer_data_3[663:656];
        layer1[18][31:24] = buffer_data_3[671:664];
        layer1[18][39:32] = buffer_data_3[679:672];
        layer2[18][7:0] = buffer_data_2[647:640];
        layer2[18][15:8] = buffer_data_2[655:648];
        layer2[18][23:16] = buffer_data_2[663:656];
        layer2[18][31:24] = buffer_data_2[671:664];
        layer2[18][39:32] = buffer_data_2[679:672];
        layer3[18][7:0] = buffer_data_1[647:640];
        layer3[18][15:8] = buffer_data_1[655:648];
        layer3[18][23:16] = buffer_data_1[663:656];
        layer3[18][31:24] = buffer_data_1[671:664];
        layer3[18][39:32] = buffer_data_1[679:672];
        layer4[18][7:0] = buffer_data_0[647:640];
        layer4[18][15:8] = buffer_data_0[655:648];
        layer4[18][23:16] = buffer_data_0[663:656];
        layer4[18][31:24] = buffer_data_0[671:664];
        layer4[18][39:32] = buffer_data_0[679:672];
        layer0[19][7:0] = buffer_data_4[655:648];
        layer0[19][15:8] = buffer_data_4[663:656];
        layer0[19][23:16] = buffer_data_4[671:664];
        layer0[19][31:24] = buffer_data_4[679:672];
        layer0[19][39:32] = buffer_data_4[687:680];
        layer1[19][7:0] = buffer_data_3[655:648];
        layer1[19][15:8] = buffer_data_3[663:656];
        layer1[19][23:16] = buffer_data_3[671:664];
        layer1[19][31:24] = buffer_data_3[679:672];
        layer1[19][39:32] = buffer_data_3[687:680];
        layer2[19][7:0] = buffer_data_2[655:648];
        layer2[19][15:8] = buffer_data_2[663:656];
        layer2[19][23:16] = buffer_data_2[671:664];
        layer2[19][31:24] = buffer_data_2[679:672];
        layer2[19][39:32] = buffer_data_2[687:680];
        layer3[19][7:0] = buffer_data_1[655:648];
        layer3[19][15:8] = buffer_data_1[663:656];
        layer3[19][23:16] = buffer_data_1[671:664];
        layer3[19][31:24] = buffer_data_1[679:672];
        layer3[19][39:32] = buffer_data_1[687:680];
        layer4[19][7:0] = buffer_data_0[655:648];
        layer4[19][15:8] = buffer_data_0[663:656];
        layer4[19][23:16] = buffer_data_0[671:664];
        layer4[19][31:24] = buffer_data_0[679:672];
        layer4[19][39:32] = buffer_data_0[687:680];
        layer0[20][7:0] = buffer_data_4[663:656];
        layer0[20][15:8] = buffer_data_4[671:664];
        layer0[20][23:16] = buffer_data_4[679:672];
        layer0[20][31:24] = buffer_data_4[687:680];
        layer0[20][39:32] = buffer_data_4[695:688];
        layer1[20][7:0] = buffer_data_3[663:656];
        layer1[20][15:8] = buffer_data_3[671:664];
        layer1[20][23:16] = buffer_data_3[679:672];
        layer1[20][31:24] = buffer_data_3[687:680];
        layer1[20][39:32] = buffer_data_3[695:688];
        layer2[20][7:0] = buffer_data_2[663:656];
        layer2[20][15:8] = buffer_data_2[671:664];
        layer2[20][23:16] = buffer_data_2[679:672];
        layer2[20][31:24] = buffer_data_2[687:680];
        layer2[20][39:32] = buffer_data_2[695:688];
        layer3[20][7:0] = buffer_data_1[663:656];
        layer3[20][15:8] = buffer_data_1[671:664];
        layer3[20][23:16] = buffer_data_1[679:672];
        layer3[20][31:24] = buffer_data_1[687:680];
        layer3[20][39:32] = buffer_data_1[695:688];
        layer4[20][7:0] = buffer_data_0[663:656];
        layer4[20][15:8] = buffer_data_0[671:664];
        layer4[20][23:16] = buffer_data_0[679:672];
        layer4[20][31:24] = buffer_data_0[687:680];
        layer4[20][39:32] = buffer_data_0[695:688];
        layer0[21][7:0] = buffer_data_4[671:664];
        layer0[21][15:8] = buffer_data_4[679:672];
        layer0[21][23:16] = buffer_data_4[687:680];
        layer0[21][31:24] = buffer_data_4[695:688];
        layer0[21][39:32] = buffer_data_4[703:696];
        layer1[21][7:0] = buffer_data_3[671:664];
        layer1[21][15:8] = buffer_data_3[679:672];
        layer1[21][23:16] = buffer_data_3[687:680];
        layer1[21][31:24] = buffer_data_3[695:688];
        layer1[21][39:32] = buffer_data_3[703:696];
        layer2[21][7:0] = buffer_data_2[671:664];
        layer2[21][15:8] = buffer_data_2[679:672];
        layer2[21][23:16] = buffer_data_2[687:680];
        layer2[21][31:24] = buffer_data_2[695:688];
        layer2[21][39:32] = buffer_data_2[703:696];
        layer3[21][7:0] = buffer_data_1[671:664];
        layer3[21][15:8] = buffer_data_1[679:672];
        layer3[21][23:16] = buffer_data_1[687:680];
        layer3[21][31:24] = buffer_data_1[695:688];
        layer3[21][39:32] = buffer_data_1[703:696];
        layer4[21][7:0] = buffer_data_0[671:664];
        layer4[21][15:8] = buffer_data_0[679:672];
        layer4[21][23:16] = buffer_data_0[687:680];
        layer4[21][31:24] = buffer_data_0[695:688];
        layer4[21][39:32] = buffer_data_0[703:696];
        layer0[22][7:0] = buffer_data_4[679:672];
        layer0[22][15:8] = buffer_data_4[687:680];
        layer0[22][23:16] = buffer_data_4[695:688];
        layer0[22][31:24] = buffer_data_4[703:696];
        layer0[22][39:32] = buffer_data_4[711:704];
        layer1[22][7:0] = buffer_data_3[679:672];
        layer1[22][15:8] = buffer_data_3[687:680];
        layer1[22][23:16] = buffer_data_3[695:688];
        layer1[22][31:24] = buffer_data_3[703:696];
        layer1[22][39:32] = buffer_data_3[711:704];
        layer2[22][7:0] = buffer_data_2[679:672];
        layer2[22][15:8] = buffer_data_2[687:680];
        layer2[22][23:16] = buffer_data_2[695:688];
        layer2[22][31:24] = buffer_data_2[703:696];
        layer2[22][39:32] = buffer_data_2[711:704];
        layer3[22][7:0] = buffer_data_1[679:672];
        layer3[22][15:8] = buffer_data_1[687:680];
        layer3[22][23:16] = buffer_data_1[695:688];
        layer3[22][31:24] = buffer_data_1[703:696];
        layer3[22][39:32] = buffer_data_1[711:704];
        layer4[22][7:0] = buffer_data_0[679:672];
        layer4[22][15:8] = buffer_data_0[687:680];
        layer4[22][23:16] = buffer_data_0[695:688];
        layer4[22][31:24] = buffer_data_0[703:696];
        layer4[22][39:32] = buffer_data_0[711:704];
        layer0[23][7:0] = buffer_data_4[687:680];
        layer0[23][15:8] = buffer_data_4[695:688];
        layer0[23][23:16] = buffer_data_4[703:696];
        layer0[23][31:24] = buffer_data_4[711:704];
        layer0[23][39:32] = buffer_data_4[719:712];
        layer1[23][7:0] = buffer_data_3[687:680];
        layer1[23][15:8] = buffer_data_3[695:688];
        layer1[23][23:16] = buffer_data_3[703:696];
        layer1[23][31:24] = buffer_data_3[711:704];
        layer1[23][39:32] = buffer_data_3[719:712];
        layer2[23][7:0] = buffer_data_2[687:680];
        layer2[23][15:8] = buffer_data_2[695:688];
        layer2[23][23:16] = buffer_data_2[703:696];
        layer2[23][31:24] = buffer_data_2[711:704];
        layer2[23][39:32] = buffer_data_2[719:712];
        layer3[23][7:0] = buffer_data_1[687:680];
        layer3[23][15:8] = buffer_data_1[695:688];
        layer3[23][23:16] = buffer_data_1[703:696];
        layer3[23][31:24] = buffer_data_1[711:704];
        layer3[23][39:32] = buffer_data_1[719:712];
        layer4[23][7:0] = buffer_data_0[687:680];
        layer4[23][15:8] = buffer_data_0[695:688];
        layer4[23][23:16] = buffer_data_0[703:696];
        layer4[23][31:24] = buffer_data_0[711:704];
        layer4[23][39:32] = buffer_data_0[719:712];
        layer0[24][7:0] = buffer_data_4[695:688];
        layer0[24][15:8] = buffer_data_4[703:696];
        layer0[24][23:16] = buffer_data_4[711:704];
        layer0[24][31:24] = buffer_data_4[719:712];
        layer0[24][39:32] = buffer_data_4[727:720];
        layer1[24][7:0] = buffer_data_3[695:688];
        layer1[24][15:8] = buffer_data_3[703:696];
        layer1[24][23:16] = buffer_data_3[711:704];
        layer1[24][31:24] = buffer_data_3[719:712];
        layer1[24][39:32] = buffer_data_3[727:720];
        layer2[24][7:0] = buffer_data_2[695:688];
        layer2[24][15:8] = buffer_data_2[703:696];
        layer2[24][23:16] = buffer_data_2[711:704];
        layer2[24][31:24] = buffer_data_2[719:712];
        layer2[24][39:32] = buffer_data_2[727:720];
        layer3[24][7:0] = buffer_data_1[695:688];
        layer3[24][15:8] = buffer_data_1[703:696];
        layer3[24][23:16] = buffer_data_1[711:704];
        layer3[24][31:24] = buffer_data_1[719:712];
        layer3[24][39:32] = buffer_data_1[727:720];
        layer4[24][7:0] = buffer_data_0[695:688];
        layer4[24][15:8] = buffer_data_0[703:696];
        layer4[24][23:16] = buffer_data_0[711:704];
        layer4[24][31:24] = buffer_data_0[719:712];
        layer4[24][39:32] = buffer_data_0[727:720];
        layer0[25][7:0] = buffer_data_4[703:696];
        layer0[25][15:8] = buffer_data_4[711:704];
        layer0[25][23:16] = buffer_data_4[719:712];
        layer0[25][31:24] = buffer_data_4[727:720];
        layer0[25][39:32] = buffer_data_4[735:728];
        layer1[25][7:0] = buffer_data_3[703:696];
        layer1[25][15:8] = buffer_data_3[711:704];
        layer1[25][23:16] = buffer_data_3[719:712];
        layer1[25][31:24] = buffer_data_3[727:720];
        layer1[25][39:32] = buffer_data_3[735:728];
        layer2[25][7:0] = buffer_data_2[703:696];
        layer2[25][15:8] = buffer_data_2[711:704];
        layer2[25][23:16] = buffer_data_2[719:712];
        layer2[25][31:24] = buffer_data_2[727:720];
        layer2[25][39:32] = buffer_data_2[735:728];
        layer3[25][7:0] = buffer_data_1[703:696];
        layer3[25][15:8] = buffer_data_1[711:704];
        layer3[25][23:16] = buffer_data_1[719:712];
        layer3[25][31:24] = buffer_data_1[727:720];
        layer3[25][39:32] = buffer_data_1[735:728];
        layer4[25][7:0] = buffer_data_0[703:696];
        layer4[25][15:8] = buffer_data_0[711:704];
        layer4[25][23:16] = buffer_data_0[719:712];
        layer4[25][31:24] = buffer_data_0[727:720];
        layer4[25][39:32] = buffer_data_0[735:728];
        layer0[26][7:0] = buffer_data_4[711:704];
        layer0[26][15:8] = buffer_data_4[719:712];
        layer0[26][23:16] = buffer_data_4[727:720];
        layer0[26][31:24] = buffer_data_4[735:728];
        layer0[26][39:32] = buffer_data_4[743:736];
        layer1[26][7:0] = buffer_data_3[711:704];
        layer1[26][15:8] = buffer_data_3[719:712];
        layer1[26][23:16] = buffer_data_3[727:720];
        layer1[26][31:24] = buffer_data_3[735:728];
        layer1[26][39:32] = buffer_data_3[743:736];
        layer2[26][7:0] = buffer_data_2[711:704];
        layer2[26][15:8] = buffer_data_2[719:712];
        layer2[26][23:16] = buffer_data_2[727:720];
        layer2[26][31:24] = buffer_data_2[735:728];
        layer2[26][39:32] = buffer_data_2[743:736];
        layer3[26][7:0] = buffer_data_1[711:704];
        layer3[26][15:8] = buffer_data_1[719:712];
        layer3[26][23:16] = buffer_data_1[727:720];
        layer3[26][31:24] = buffer_data_1[735:728];
        layer3[26][39:32] = buffer_data_1[743:736];
        layer4[26][7:0] = buffer_data_0[711:704];
        layer4[26][15:8] = buffer_data_0[719:712];
        layer4[26][23:16] = buffer_data_0[727:720];
        layer4[26][31:24] = buffer_data_0[735:728];
        layer4[26][39:32] = buffer_data_0[743:736];
        layer0[27][7:0] = buffer_data_4[719:712];
        layer0[27][15:8] = buffer_data_4[727:720];
        layer0[27][23:16] = buffer_data_4[735:728];
        layer0[27][31:24] = buffer_data_4[743:736];
        layer0[27][39:32] = buffer_data_4[751:744];
        layer1[27][7:0] = buffer_data_3[719:712];
        layer1[27][15:8] = buffer_data_3[727:720];
        layer1[27][23:16] = buffer_data_3[735:728];
        layer1[27][31:24] = buffer_data_3[743:736];
        layer1[27][39:32] = buffer_data_3[751:744];
        layer2[27][7:0] = buffer_data_2[719:712];
        layer2[27][15:8] = buffer_data_2[727:720];
        layer2[27][23:16] = buffer_data_2[735:728];
        layer2[27][31:24] = buffer_data_2[743:736];
        layer2[27][39:32] = buffer_data_2[751:744];
        layer3[27][7:0] = buffer_data_1[719:712];
        layer3[27][15:8] = buffer_data_1[727:720];
        layer3[27][23:16] = buffer_data_1[735:728];
        layer3[27][31:24] = buffer_data_1[743:736];
        layer3[27][39:32] = buffer_data_1[751:744];
        layer4[27][7:0] = buffer_data_0[719:712];
        layer4[27][15:8] = buffer_data_0[727:720];
        layer4[27][23:16] = buffer_data_0[735:728];
        layer4[27][31:24] = buffer_data_0[743:736];
        layer4[27][39:32] = buffer_data_0[751:744];
        layer0[28][7:0] = buffer_data_4[727:720];
        layer0[28][15:8] = buffer_data_4[735:728];
        layer0[28][23:16] = buffer_data_4[743:736];
        layer0[28][31:24] = buffer_data_4[751:744];
        layer0[28][39:32] = buffer_data_4[759:752];
        layer1[28][7:0] = buffer_data_3[727:720];
        layer1[28][15:8] = buffer_data_3[735:728];
        layer1[28][23:16] = buffer_data_3[743:736];
        layer1[28][31:24] = buffer_data_3[751:744];
        layer1[28][39:32] = buffer_data_3[759:752];
        layer2[28][7:0] = buffer_data_2[727:720];
        layer2[28][15:8] = buffer_data_2[735:728];
        layer2[28][23:16] = buffer_data_2[743:736];
        layer2[28][31:24] = buffer_data_2[751:744];
        layer2[28][39:32] = buffer_data_2[759:752];
        layer3[28][7:0] = buffer_data_1[727:720];
        layer3[28][15:8] = buffer_data_1[735:728];
        layer3[28][23:16] = buffer_data_1[743:736];
        layer3[28][31:24] = buffer_data_1[751:744];
        layer3[28][39:32] = buffer_data_1[759:752];
        layer4[28][7:0] = buffer_data_0[727:720];
        layer4[28][15:8] = buffer_data_0[735:728];
        layer4[28][23:16] = buffer_data_0[743:736];
        layer4[28][31:24] = buffer_data_0[751:744];
        layer4[28][39:32] = buffer_data_0[759:752];
        layer0[29][7:0] = buffer_data_4[735:728];
        layer0[29][15:8] = buffer_data_4[743:736];
        layer0[29][23:16] = buffer_data_4[751:744];
        layer0[29][31:24] = buffer_data_4[759:752];
        layer0[29][39:32] = buffer_data_4[767:760];
        layer1[29][7:0] = buffer_data_3[735:728];
        layer1[29][15:8] = buffer_data_3[743:736];
        layer1[29][23:16] = buffer_data_3[751:744];
        layer1[29][31:24] = buffer_data_3[759:752];
        layer1[29][39:32] = buffer_data_3[767:760];
        layer2[29][7:0] = buffer_data_2[735:728];
        layer2[29][15:8] = buffer_data_2[743:736];
        layer2[29][23:16] = buffer_data_2[751:744];
        layer2[29][31:24] = buffer_data_2[759:752];
        layer2[29][39:32] = buffer_data_2[767:760];
        layer3[29][7:0] = buffer_data_1[735:728];
        layer3[29][15:8] = buffer_data_1[743:736];
        layer3[29][23:16] = buffer_data_1[751:744];
        layer3[29][31:24] = buffer_data_1[759:752];
        layer3[29][39:32] = buffer_data_1[767:760];
        layer4[29][7:0] = buffer_data_0[735:728];
        layer4[29][15:8] = buffer_data_0[743:736];
        layer4[29][23:16] = buffer_data_0[751:744];
        layer4[29][31:24] = buffer_data_0[759:752];
        layer4[29][39:32] = buffer_data_0[767:760];
        layer0[30][7:0] = buffer_data_4[743:736];
        layer0[30][15:8] = buffer_data_4[751:744];
        layer0[30][23:16] = buffer_data_4[759:752];
        layer0[30][31:24] = buffer_data_4[767:760];
        layer0[30][39:32] = buffer_data_4[775:768];
        layer1[30][7:0] = buffer_data_3[743:736];
        layer1[30][15:8] = buffer_data_3[751:744];
        layer1[30][23:16] = buffer_data_3[759:752];
        layer1[30][31:24] = buffer_data_3[767:760];
        layer1[30][39:32] = buffer_data_3[775:768];
        layer2[30][7:0] = buffer_data_2[743:736];
        layer2[30][15:8] = buffer_data_2[751:744];
        layer2[30][23:16] = buffer_data_2[759:752];
        layer2[30][31:24] = buffer_data_2[767:760];
        layer2[30][39:32] = buffer_data_2[775:768];
        layer3[30][7:0] = buffer_data_1[743:736];
        layer3[30][15:8] = buffer_data_1[751:744];
        layer3[30][23:16] = buffer_data_1[759:752];
        layer3[30][31:24] = buffer_data_1[767:760];
        layer3[30][39:32] = buffer_data_1[775:768];
        layer4[30][7:0] = buffer_data_0[743:736];
        layer4[30][15:8] = buffer_data_0[751:744];
        layer4[30][23:16] = buffer_data_0[759:752];
        layer4[30][31:24] = buffer_data_0[767:760];
        layer4[30][39:32] = buffer_data_0[775:768];
        layer0[31][7:0] = buffer_data_4[751:744];
        layer0[31][15:8] = buffer_data_4[759:752];
        layer0[31][23:16] = buffer_data_4[767:760];
        layer0[31][31:24] = buffer_data_4[775:768];
        layer0[31][39:32] = buffer_data_4[783:776];
        layer1[31][7:0] = buffer_data_3[751:744];
        layer1[31][15:8] = buffer_data_3[759:752];
        layer1[31][23:16] = buffer_data_3[767:760];
        layer1[31][31:24] = buffer_data_3[775:768];
        layer1[31][39:32] = buffer_data_3[783:776];
        layer2[31][7:0] = buffer_data_2[751:744];
        layer2[31][15:8] = buffer_data_2[759:752];
        layer2[31][23:16] = buffer_data_2[767:760];
        layer2[31][31:24] = buffer_data_2[775:768];
        layer2[31][39:32] = buffer_data_2[783:776];
        layer3[31][7:0] = buffer_data_1[751:744];
        layer3[31][15:8] = buffer_data_1[759:752];
        layer3[31][23:16] = buffer_data_1[767:760];
        layer3[31][31:24] = buffer_data_1[775:768];
        layer3[31][39:32] = buffer_data_1[783:776];
        layer4[31][7:0] = buffer_data_0[751:744];
        layer4[31][15:8] = buffer_data_0[759:752];
        layer4[31][23:16] = buffer_data_0[767:760];
        layer4[31][31:24] = buffer_data_0[775:768];
        layer4[31][39:32] = buffer_data_0[783:776];
        layer0[32][7:0] = buffer_data_4[759:752];
        layer0[32][15:8] = buffer_data_4[767:760];
        layer0[32][23:16] = buffer_data_4[775:768];
        layer0[32][31:24] = buffer_data_4[783:776];
        layer0[32][39:32] = buffer_data_4[791:784];
        layer1[32][7:0] = buffer_data_3[759:752];
        layer1[32][15:8] = buffer_data_3[767:760];
        layer1[32][23:16] = buffer_data_3[775:768];
        layer1[32][31:24] = buffer_data_3[783:776];
        layer1[32][39:32] = buffer_data_3[791:784];
        layer2[32][7:0] = buffer_data_2[759:752];
        layer2[32][15:8] = buffer_data_2[767:760];
        layer2[32][23:16] = buffer_data_2[775:768];
        layer2[32][31:24] = buffer_data_2[783:776];
        layer2[32][39:32] = buffer_data_2[791:784];
        layer3[32][7:0] = buffer_data_1[759:752];
        layer3[32][15:8] = buffer_data_1[767:760];
        layer3[32][23:16] = buffer_data_1[775:768];
        layer3[32][31:24] = buffer_data_1[783:776];
        layer3[32][39:32] = buffer_data_1[791:784];
        layer4[32][7:0] = buffer_data_0[759:752];
        layer4[32][15:8] = buffer_data_0[767:760];
        layer4[32][23:16] = buffer_data_0[775:768];
        layer4[32][31:24] = buffer_data_0[783:776];
        layer4[32][39:32] = buffer_data_0[791:784];
        layer0[33][7:0] = buffer_data_4[767:760];
        layer0[33][15:8] = buffer_data_4[775:768];
        layer0[33][23:16] = buffer_data_4[783:776];
        layer0[33][31:24] = buffer_data_4[791:784];
        layer0[33][39:32] = buffer_data_4[799:792];
        layer1[33][7:0] = buffer_data_3[767:760];
        layer1[33][15:8] = buffer_data_3[775:768];
        layer1[33][23:16] = buffer_data_3[783:776];
        layer1[33][31:24] = buffer_data_3[791:784];
        layer1[33][39:32] = buffer_data_3[799:792];
        layer2[33][7:0] = buffer_data_2[767:760];
        layer2[33][15:8] = buffer_data_2[775:768];
        layer2[33][23:16] = buffer_data_2[783:776];
        layer2[33][31:24] = buffer_data_2[791:784];
        layer2[33][39:32] = buffer_data_2[799:792];
        layer3[33][7:0] = buffer_data_1[767:760];
        layer3[33][15:8] = buffer_data_1[775:768];
        layer3[33][23:16] = buffer_data_1[783:776];
        layer3[33][31:24] = buffer_data_1[791:784];
        layer3[33][39:32] = buffer_data_1[799:792];
        layer4[33][7:0] = buffer_data_0[767:760];
        layer4[33][15:8] = buffer_data_0[775:768];
        layer4[33][23:16] = buffer_data_0[783:776];
        layer4[33][31:24] = buffer_data_0[791:784];
        layer4[33][39:32] = buffer_data_0[799:792];
        layer0[34][7:0] = buffer_data_4[775:768];
        layer0[34][15:8] = buffer_data_4[783:776];
        layer0[34][23:16] = buffer_data_4[791:784];
        layer0[34][31:24] = buffer_data_4[799:792];
        layer0[34][39:32] = buffer_data_4[807:800];
        layer1[34][7:0] = buffer_data_3[775:768];
        layer1[34][15:8] = buffer_data_3[783:776];
        layer1[34][23:16] = buffer_data_3[791:784];
        layer1[34][31:24] = buffer_data_3[799:792];
        layer1[34][39:32] = buffer_data_3[807:800];
        layer2[34][7:0] = buffer_data_2[775:768];
        layer2[34][15:8] = buffer_data_2[783:776];
        layer2[34][23:16] = buffer_data_2[791:784];
        layer2[34][31:24] = buffer_data_2[799:792];
        layer2[34][39:32] = buffer_data_2[807:800];
        layer3[34][7:0] = buffer_data_1[775:768];
        layer3[34][15:8] = buffer_data_1[783:776];
        layer3[34][23:16] = buffer_data_1[791:784];
        layer3[34][31:24] = buffer_data_1[799:792];
        layer3[34][39:32] = buffer_data_1[807:800];
        layer4[34][7:0] = buffer_data_0[775:768];
        layer4[34][15:8] = buffer_data_0[783:776];
        layer4[34][23:16] = buffer_data_0[791:784];
        layer4[34][31:24] = buffer_data_0[799:792];
        layer4[34][39:32] = buffer_data_0[807:800];
        layer0[35][7:0] = buffer_data_4[783:776];
        layer0[35][15:8] = buffer_data_4[791:784];
        layer0[35][23:16] = buffer_data_4[799:792];
        layer0[35][31:24] = buffer_data_4[807:800];
        layer0[35][39:32] = buffer_data_4[815:808];
        layer1[35][7:0] = buffer_data_3[783:776];
        layer1[35][15:8] = buffer_data_3[791:784];
        layer1[35][23:16] = buffer_data_3[799:792];
        layer1[35][31:24] = buffer_data_3[807:800];
        layer1[35][39:32] = buffer_data_3[815:808];
        layer2[35][7:0] = buffer_data_2[783:776];
        layer2[35][15:8] = buffer_data_2[791:784];
        layer2[35][23:16] = buffer_data_2[799:792];
        layer2[35][31:24] = buffer_data_2[807:800];
        layer2[35][39:32] = buffer_data_2[815:808];
        layer3[35][7:0] = buffer_data_1[783:776];
        layer3[35][15:8] = buffer_data_1[791:784];
        layer3[35][23:16] = buffer_data_1[799:792];
        layer3[35][31:24] = buffer_data_1[807:800];
        layer3[35][39:32] = buffer_data_1[815:808];
        layer4[35][7:0] = buffer_data_0[783:776];
        layer4[35][15:8] = buffer_data_0[791:784];
        layer4[35][23:16] = buffer_data_0[799:792];
        layer4[35][31:24] = buffer_data_0[807:800];
        layer4[35][39:32] = buffer_data_0[815:808];
        layer0[36][7:0] = buffer_data_4[791:784];
        layer0[36][15:8] = buffer_data_4[799:792];
        layer0[36][23:16] = buffer_data_4[807:800];
        layer0[36][31:24] = buffer_data_4[815:808];
        layer0[36][39:32] = buffer_data_4[823:816];
        layer1[36][7:0] = buffer_data_3[791:784];
        layer1[36][15:8] = buffer_data_3[799:792];
        layer1[36][23:16] = buffer_data_3[807:800];
        layer1[36][31:24] = buffer_data_3[815:808];
        layer1[36][39:32] = buffer_data_3[823:816];
        layer2[36][7:0] = buffer_data_2[791:784];
        layer2[36][15:8] = buffer_data_2[799:792];
        layer2[36][23:16] = buffer_data_2[807:800];
        layer2[36][31:24] = buffer_data_2[815:808];
        layer2[36][39:32] = buffer_data_2[823:816];
        layer3[36][7:0] = buffer_data_1[791:784];
        layer3[36][15:8] = buffer_data_1[799:792];
        layer3[36][23:16] = buffer_data_1[807:800];
        layer3[36][31:24] = buffer_data_1[815:808];
        layer3[36][39:32] = buffer_data_1[823:816];
        layer4[36][7:0] = buffer_data_0[791:784];
        layer4[36][15:8] = buffer_data_0[799:792];
        layer4[36][23:16] = buffer_data_0[807:800];
        layer4[36][31:24] = buffer_data_0[815:808];
        layer4[36][39:32] = buffer_data_0[823:816];
        layer0[37][7:0] = buffer_data_4[799:792];
        layer0[37][15:8] = buffer_data_4[807:800];
        layer0[37][23:16] = buffer_data_4[815:808];
        layer0[37][31:24] = buffer_data_4[823:816];
        layer0[37][39:32] = buffer_data_4[831:824];
        layer1[37][7:0] = buffer_data_3[799:792];
        layer1[37][15:8] = buffer_data_3[807:800];
        layer1[37][23:16] = buffer_data_3[815:808];
        layer1[37][31:24] = buffer_data_3[823:816];
        layer1[37][39:32] = buffer_data_3[831:824];
        layer2[37][7:0] = buffer_data_2[799:792];
        layer2[37][15:8] = buffer_data_2[807:800];
        layer2[37][23:16] = buffer_data_2[815:808];
        layer2[37][31:24] = buffer_data_2[823:816];
        layer2[37][39:32] = buffer_data_2[831:824];
        layer3[37][7:0] = buffer_data_1[799:792];
        layer3[37][15:8] = buffer_data_1[807:800];
        layer3[37][23:16] = buffer_data_1[815:808];
        layer3[37][31:24] = buffer_data_1[823:816];
        layer3[37][39:32] = buffer_data_1[831:824];
        layer4[37][7:0] = buffer_data_0[799:792];
        layer4[37][15:8] = buffer_data_0[807:800];
        layer4[37][23:16] = buffer_data_0[815:808];
        layer4[37][31:24] = buffer_data_0[823:816];
        layer4[37][39:32] = buffer_data_0[831:824];
        layer0[38][7:0] = buffer_data_4[807:800];
        layer0[38][15:8] = buffer_data_4[815:808];
        layer0[38][23:16] = buffer_data_4[823:816];
        layer0[38][31:24] = buffer_data_4[831:824];
        layer0[38][39:32] = buffer_data_4[839:832];
        layer1[38][7:0] = buffer_data_3[807:800];
        layer1[38][15:8] = buffer_data_3[815:808];
        layer1[38][23:16] = buffer_data_3[823:816];
        layer1[38][31:24] = buffer_data_3[831:824];
        layer1[38][39:32] = buffer_data_3[839:832];
        layer2[38][7:0] = buffer_data_2[807:800];
        layer2[38][15:8] = buffer_data_2[815:808];
        layer2[38][23:16] = buffer_data_2[823:816];
        layer2[38][31:24] = buffer_data_2[831:824];
        layer2[38][39:32] = buffer_data_2[839:832];
        layer3[38][7:0] = buffer_data_1[807:800];
        layer3[38][15:8] = buffer_data_1[815:808];
        layer3[38][23:16] = buffer_data_1[823:816];
        layer3[38][31:24] = buffer_data_1[831:824];
        layer3[38][39:32] = buffer_data_1[839:832];
        layer4[38][7:0] = buffer_data_0[807:800];
        layer4[38][15:8] = buffer_data_0[815:808];
        layer4[38][23:16] = buffer_data_0[823:816];
        layer4[38][31:24] = buffer_data_0[831:824];
        layer4[38][39:32] = buffer_data_0[839:832];
        layer0[39][7:0] = buffer_data_4[815:808];
        layer0[39][15:8] = buffer_data_4[823:816];
        layer0[39][23:16] = buffer_data_4[831:824];
        layer0[39][31:24] = buffer_data_4[839:832];
        layer0[39][39:32] = buffer_data_4[847:840];
        layer1[39][7:0] = buffer_data_3[815:808];
        layer1[39][15:8] = buffer_data_3[823:816];
        layer1[39][23:16] = buffer_data_3[831:824];
        layer1[39][31:24] = buffer_data_3[839:832];
        layer1[39][39:32] = buffer_data_3[847:840];
        layer2[39][7:0] = buffer_data_2[815:808];
        layer2[39][15:8] = buffer_data_2[823:816];
        layer2[39][23:16] = buffer_data_2[831:824];
        layer2[39][31:24] = buffer_data_2[839:832];
        layer2[39][39:32] = buffer_data_2[847:840];
        layer3[39][7:0] = buffer_data_1[815:808];
        layer3[39][15:8] = buffer_data_1[823:816];
        layer3[39][23:16] = buffer_data_1[831:824];
        layer3[39][31:24] = buffer_data_1[839:832];
        layer3[39][39:32] = buffer_data_1[847:840];
        layer4[39][7:0] = buffer_data_0[815:808];
        layer4[39][15:8] = buffer_data_0[823:816];
        layer4[39][23:16] = buffer_data_0[831:824];
        layer4[39][31:24] = buffer_data_0[839:832];
        layer4[39][39:32] = buffer_data_0[847:840];
        layer0[40][7:0] = buffer_data_4[823:816];
        layer0[40][15:8] = buffer_data_4[831:824];
        layer0[40][23:16] = buffer_data_4[839:832];
        layer0[40][31:24] = buffer_data_4[847:840];
        layer0[40][39:32] = buffer_data_4[855:848];
        layer1[40][7:0] = buffer_data_3[823:816];
        layer1[40][15:8] = buffer_data_3[831:824];
        layer1[40][23:16] = buffer_data_3[839:832];
        layer1[40][31:24] = buffer_data_3[847:840];
        layer1[40][39:32] = buffer_data_3[855:848];
        layer2[40][7:0] = buffer_data_2[823:816];
        layer2[40][15:8] = buffer_data_2[831:824];
        layer2[40][23:16] = buffer_data_2[839:832];
        layer2[40][31:24] = buffer_data_2[847:840];
        layer2[40][39:32] = buffer_data_2[855:848];
        layer3[40][7:0] = buffer_data_1[823:816];
        layer3[40][15:8] = buffer_data_1[831:824];
        layer3[40][23:16] = buffer_data_1[839:832];
        layer3[40][31:24] = buffer_data_1[847:840];
        layer3[40][39:32] = buffer_data_1[855:848];
        layer4[40][7:0] = buffer_data_0[823:816];
        layer4[40][15:8] = buffer_data_0[831:824];
        layer4[40][23:16] = buffer_data_0[839:832];
        layer4[40][31:24] = buffer_data_0[847:840];
        layer4[40][39:32] = buffer_data_0[855:848];
        layer0[41][7:0] = buffer_data_4[831:824];
        layer0[41][15:8] = buffer_data_4[839:832];
        layer0[41][23:16] = buffer_data_4[847:840];
        layer0[41][31:24] = buffer_data_4[855:848];
        layer0[41][39:32] = buffer_data_4[863:856];
        layer1[41][7:0] = buffer_data_3[831:824];
        layer1[41][15:8] = buffer_data_3[839:832];
        layer1[41][23:16] = buffer_data_3[847:840];
        layer1[41][31:24] = buffer_data_3[855:848];
        layer1[41][39:32] = buffer_data_3[863:856];
        layer2[41][7:0] = buffer_data_2[831:824];
        layer2[41][15:8] = buffer_data_2[839:832];
        layer2[41][23:16] = buffer_data_2[847:840];
        layer2[41][31:24] = buffer_data_2[855:848];
        layer2[41][39:32] = buffer_data_2[863:856];
        layer3[41][7:0] = buffer_data_1[831:824];
        layer3[41][15:8] = buffer_data_1[839:832];
        layer3[41][23:16] = buffer_data_1[847:840];
        layer3[41][31:24] = buffer_data_1[855:848];
        layer3[41][39:32] = buffer_data_1[863:856];
        layer4[41][7:0] = buffer_data_0[831:824];
        layer4[41][15:8] = buffer_data_0[839:832];
        layer4[41][23:16] = buffer_data_0[847:840];
        layer4[41][31:24] = buffer_data_0[855:848];
        layer4[41][39:32] = buffer_data_0[863:856];
        layer0[42][7:0] = buffer_data_4[839:832];
        layer0[42][15:8] = buffer_data_4[847:840];
        layer0[42][23:16] = buffer_data_4[855:848];
        layer0[42][31:24] = buffer_data_4[863:856];
        layer0[42][39:32] = buffer_data_4[871:864];
        layer1[42][7:0] = buffer_data_3[839:832];
        layer1[42][15:8] = buffer_data_3[847:840];
        layer1[42][23:16] = buffer_data_3[855:848];
        layer1[42][31:24] = buffer_data_3[863:856];
        layer1[42][39:32] = buffer_data_3[871:864];
        layer2[42][7:0] = buffer_data_2[839:832];
        layer2[42][15:8] = buffer_data_2[847:840];
        layer2[42][23:16] = buffer_data_2[855:848];
        layer2[42][31:24] = buffer_data_2[863:856];
        layer2[42][39:32] = buffer_data_2[871:864];
        layer3[42][7:0] = buffer_data_1[839:832];
        layer3[42][15:8] = buffer_data_1[847:840];
        layer3[42][23:16] = buffer_data_1[855:848];
        layer3[42][31:24] = buffer_data_1[863:856];
        layer3[42][39:32] = buffer_data_1[871:864];
        layer4[42][7:0] = buffer_data_0[839:832];
        layer4[42][15:8] = buffer_data_0[847:840];
        layer4[42][23:16] = buffer_data_0[855:848];
        layer4[42][31:24] = buffer_data_0[863:856];
        layer4[42][39:32] = buffer_data_0[871:864];
        layer0[43][7:0] = buffer_data_4[847:840];
        layer0[43][15:8] = buffer_data_4[855:848];
        layer0[43][23:16] = buffer_data_4[863:856];
        layer0[43][31:24] = buffer_data_4[871:864];
        layer0[43][39:32] = buffer_data_4[879:872];
        layer1[43][7:0] = buffer_data_3[847:840];
        layer1[43][15:8] = buffer_data_3[855:848];
        layer1[43][23:16] = buffer_data_3[863:856];
        layer1[43][31:24] = buffer_data_3[871:864];
        layer1[43][39:32] = buffer_data_3[879:872];
        layer2[43][7:0] = buffer_data_2[847:840];
        layer2[43][15:8] = buffer_data_2[855:848];
        layer2[43][23:16] = buffer_data_2[863:856];
        layer2[43][31:24] = buffer_data_2[871:864];
        layer2[43][39:32] = buffer_data_2[879:872];
        layer3[43][7:0] = buffer_data_1[847:840];
        layer3[43][15:8] = buffer_data_1[855:848];
        layer3[43][23:16] = buffer_data_1[863:856];
        layer3[43][31:24] = buffer_data_1[871:864];
        layer3[43][39:32] = buffer_data_1[879:872];
        layer4[43][7:0] = buffer_data_0[847:840];
        layer4[43][15:8] = buffer_data_0[855:848];
        layer4[43][23:16] = buffer_data_0[863:856];
        layer4[43][31:24] = buffer_data_0[871:864];
        layer4[43][39:32] = buffer_data_0[879:872];
        layer0[44][7:0] = buffer_data_4[855:848];
        layer0[44][15:8] = buffer_data_4[863:856];
        layer0[44][23:16] = buffer_data_4[871:864];
        layer0[44][31:24] = buffer_data_4[879:872];
        layer0[44][39:32] = buffer_data_4[887:880];
        layer1[44][7:0] = buffer_data_3[855:848];
        layer1[44][15:8] = buffer_data_3[863:856];
        layer1[44][23:16] = buffer_data_3[871:864];
        layer1[44][31:24] = buffer_data_3[879:872];
        layer1[44][39:32] = buffer_data_3[887:880];
        layer2[44][7:0] = buffer_data_2[855:848];
        layer2[44][15:8] = buffer_data_2[863:856];
        layer2[44][23:16] = buffer_data_2[871:864];
        layer2[44][31:24] = buffer_data_2[879:872];
        layer2[44][39:32] = buffer_data_2[887:880];
        layer3[44][7:0] = buffer_data_1[855:848];
        layer3[44][15:8] = buffer_data_1[863:856];
        layer3[44][23:16] = buffer_data_1[871:864];
        layer3[44][31:24] = buffer_data_1[879:872];
        layer3[44][39:32] = buffer_data_1[887:880];
        layer4[44][7:0] = buffer_data_0[855:848];
        layer4[44][15:8] = buffer_data_0[863:856];
        layer4[44][23:16] = buffer_data_0[871:864];
        layer4[44][31:24] = buffer_data_0[879:872];
        layer4[44][39:32] = buffer_data_0[887:880];
        layer0[45][7:0] = buffer_data_4[863:856];
        layer0[45][15:8] = buffer_data_4[871:864];
        layer0[45][23:16] = buffer_data_4[879:872];
        layer0[45][31:24] = buffer_data_4[887:880];
        layer0[45][39:32] = buffer_data_4[895:888];
        layer1[45][7:0] = buffer_data_3[863:856];
        layer1[45][15:8] = buffer_data_3[871:864];
        layer1[45][23:16] = buffer_data_3[879:872];
        layer1[45][31:24] = buffer_data_3[887:880];
        layer1[45][39:32] = buffer_data_3[895:888];
        layer2[45][7:0] = buffer_data_2[863:856];
        layer2[45][15:8] = buffer_data_2[871:864];
        layer2[45][23:16] = buffer_data_2[879:872];
        layer2[45][31:24] = buffer_data_2[887:880];
        layer2[45][39:32] = buffer_data_2[895:888];
        layer3[45][7:0] = buffer_data_1[863:856];
        layer3[45][15:8] = buffer_data_1[871:864];
        layer3[45][23:16] = buffer_data_1[879:872];
        layer3[45][31:24] = buffer_data_1[887:880];
        layer3[45][39:32] = buffer_data_1[895:888];
        layer4[45][7:0] = buffer_data_0[863:856];
        layer4[45][15:8] = buffer_data_0[871:864];
        layer4[45][23:16] = buffer_data_0[879:872];
        layer4[45][31:24] = buffer_data_0[887:880];
        layer4[45][39:32] = buffer_data_0[895:888];
        layer0[46][7:0] = buffer_data_4[871:864];
        layer0[46][15:8] = buffer_data_4[879:872];
        layer0[46][23:16] = buffer_data_4[887:880];
        layer0[46][31:24] = buffer_data_4[895:888];
        layer0[46][39:32] = buffer_data_4[903:896];
        layer1[46][7:0] = buffer_data_3[871:864];
        layer1[46][15:8] = buffer_data_3[879:872];
        layer1[46][23:16] = buffer_data_3[887:880];
        layer1[46][31:24] = buffer_data_3[895:888];
        layer1[46][39:32] = buffer_data_3[903:896];
        layer2[46][7:0] = buffer_data_2[871:864];
        layer2[46][15:8] = buffer_data_2[879:872];
        layer2[46][23:16] = buffer_data_2[887:880];
        layer2[46][31:24] = buffer_data_2[895:888];
        layer2[46][39:32] = buffer_data_2[903:896];
        layer3[46][7:0] = buffer_data_1[871:864];
        layer3[46][15:8] = buffer_data_1[879:872];
        layer3[46][23:16] = buffer_data_1[887:880];
        layer3[46][31:24] = buffer_data_1[895:888];
        layer3[46][39:32] = buffer_data_1[903:896];
        layer4[46][7:0] = buffer_data_0[871:864];
        layer4[46][15:8] = buffer_data_0[879:872];
        layer4[46][23:16] = buffer_data_0[887:880];
        layer4[46][31:24] = buffer_data_0[895:888];
        layer4[46][39:32] = buffer_data_0[903:896];
        layer0[47][7:0] = buffer_data_4[879:872];
        layer0[47][15:8] = buffer_data_4[887:880];
        layer0[47][23:16] = buffer_data_4[895:888];
        layer0[47][31:24] = buffer_data_4[903:896];
        layer0[47][39:32] = buffer_data_4[911:904];
        layer1[47][7:0] = buffer_data_3[879:872];
        layer1[47][15:8] = buffer_data_3[887:880];
        layer1[47][23:16] = buffer_data_3[895:888];
        layer1[47][31:24] = buffer_data_3[903:896];
        layer1[47][39:32] = buffer_data_3[911:904];
        layer2[47][7:0] = buffer_data_2[879:872];
        layer2[47][15:8] = buffer_data_2[887:880];
        layer2[47][23:16] = buffer_data_2[895:888];
        layer2[47][31:24] = buffer_data_2[903:896];
        layer2[47][39:32] = buffer_data_2[911:904];
        layer3[47][7:0] = buffer_data_1[879:872];
        layer3[47][15:8] = buffer_data_1[887:880];
        layer3[47][23:16] = buffer_data_1[895:888];
        layer3[47][31:24] = buffer_data_1[903:896];
        layer3[47][39:32] = buffer_data_1[911:904];
        layer4[47][7:0] = buffer_data_0[879:872];
        layer4[47][15:8] = buffer_data_0[887:880];
        layer4[47][23:16] = buffer_data_0[895:888];
        layer4[47][31:24] = buffer_data_0[903:896];
        layer4[47][39:32] = buffer_data_0[911:904];
        layer0[48][7:0] = buffer_data_4[887:880];
        layer0[48][15:8] = buffer_data_4[895:888];
        layer0[48][23:16] = buffer_data_4[903:896];
        layer0[48][31:24] = buffer_data_4[911:904];
        layer0[48][39:32] = buffer_data_4[919:912];
        layer1[48][7:0] = buffer_data_3[887:880];
        layer1[48][15:8] = buffer_data_3[895:888];
        layer1[48][23:16] = buffer_data_3[903:896];
        layer1[48][31:24] = buffer_data_3[911:904];
        layer1[48][39:32] = buffer_data_3[919:912];
        layer2[48][7:0] = buffer_data_2[887:880];
        layer2[48][15:8] = buffer_data_2[895:888];
        layer2[48][23:16] = buffer_data_2[903:896];
        layer2[48][31:24] = buffer_data_2[911:904];
        layer2[48][39:32] = buffer_data_2[919:912];
        layer3[48][7:0] = buffer_data_1[887:880];
        layer3[48][15:8] = buffer_data_1[895:888];
        layer3[48][23:16] = buffer_data_1[903:896];
        layer3[48][31:24] = buffer_data_1[911:904];
        layer3[48][39:32] = buffer_data_1[919:912];
        layer4[48][7:0] = buffer_data_0[887:880];
        layer4[48][15:8] = buffer_data_0[895:888];
        layer4[48][23:16] = buffer_data_0[903:896];
        layer4[48][31:24] = buffer_data_0[911:904];
        layer4[48][39:32] = buffer_data_0[919:912];
        layer0[49][7:0] = buffer_data_4[895:888];
        layer0[49][15:8] = buffer_data_4[903:896];
        layer0[49][23:16] = buffer_data_4[911:904];
        layer0[49][31:24] = buffer_data_4[919:912];
        layer0[49][39:32] = buffer_data_4[927:920];
        layer1[49][7:0] = buffer_data_3[895:888];
        layer1[49][15:8] = buffer_data_3[903:896];
        layer1[49][23:16] = buffer_data_3[911:904];
        layer1[49][31:24] = buffer_data_3[919:912];
        layer1[49][39:32] = buffer_data_3[927:920];
        layer2[49][7:0] = buffer_data_2[895:888];
        layer2[49][15:8] = buffer_data_2[903:896];
        layer2[49][23:16] = buffer_data_2[911:904];
        layer2[49][31:24] = buffer_data_2[919:912];
        layer2[49][39:32] = buffer_data_2[927:920];
        layer3[49][7:0] = buffer_data_1[895:888];
        layer3[49][15:8] = buffer_data_1[903:896];
        layer3[49][23:16] = buffer_data_1[911:904];
        layer3[49][31:24] = buffer_data_1[919:912];
        layer3[49][39:32] = buffer_data_1[927:920];
        layer4[49][7:0] = buffer_data_0[895:888];
        layer4[49][15:8] = buffer_data_0[903:896];
        layer4[49][23:16] = buffer_data_0[911:904];
        layer4[49][31:24] = buffer_data_0[919:912];
        layer4[49][39:32] = buffer_data_0[927:920];
        layer0[50][7:0] = buffer_data_4[903:896];
        layer0[50][15:8] = buffer_data_4[911:904];
        layer0[50][23:16] = buffer_data_4[919:912];
        layer0[50][31:24] = buffer_data_4[927:920];
        layer0[50][39:32] = buffer_data_4[935:928];
        layer1[50][7:0] = buffer_data_3[903:896];
        layer1[50][15:8] = buffer_data_3[911:904];
        layer1[50][23:16] = buffer_data_3[919:912];
        layer1[50][31:24] = buffer_data_3[927:920];
        layer1[50][39:32] = buffer_data_3[935:928];
        layer2[50][7:0] = buffer_data_2[903:896];
        layer2[50][15:8] = buffer_data_2[911:904];
        layer2[50][23:16] = buffer_data_2[919:912];
        layer2[50][31:24] = buffer_data_2[927:920];
        layer2[50][39:32] = buffer_data_2[935:928];
        layer3[50][7:0] = buffer_data_1[903:896];
        layer3[50][15:8] = buffer_data_1[911:904];
        layer3[50][23:16] = buffer_data_1[919:912];
        layer3[50][31:24] = buffer_data_1[927:920];
        layer3[50][39:32] = buffer_data_1[935:928];
        layer4[50][7:0] = buffer_data_0[903:896];
        layer4[50][15:8] = buffer_data_0[911:904];
        layer4[50][23:16] = buffer_data_0[919:912];
        layer4[50][31:24] = buffer_data_0[927:920];
        layer4[50][39:32] = buffer_data_0[935:928];
        layer0[51][7:0] = buffer_data_4[911:904];
        layer0[51][15:8] = buffer_data_4[919:912];
        layer0[51][23:16] = buffer_data_4[927:920];
        layer0[51][31:24] = buffer_data_4[935:928];
        layer0[51][39:32] = buffer_data_4[943:936];
        layer1[51][7:0] = buffer_data_3[911:904];
        layer1[51][15:8] = buffer_data_3[919:912];
        layer1[51][23:16] = buffer_data_3[927:920];
        layer1[51][31:24] = buffer_data_3[935:928];
        layer1[51][39:32] = buffer_data_3[943:936];
        layer2[51][7:0] = buffer_data_2[911:904];
        layer2[51][15:8] = buffer_data_2[919:912];
        layer2[51][23:16] = buffer_data_2[927:920];
        layer2[51][31:24] = buffer_data_2[935:928];
        layer2[51][39:32] = buffer_data_2[943:936];
        layer3[51][7:0] = buffer_data_1[911:904];
        layer3[51][15:8] = buffer_data_1[919:912];
        layer3[51][23:16] = buffer_data_1[927:920];
        layer3[51][31:24] = buffer_data_1[935:928];
        layer3[51][39:32] = buffer_data_1[943:936];
        layer4[51][7:0] = buffer_data_0[911:904];
        layer4[51][15:8] = buffer_data_0[919:912];
        layer4[51][23:16] = buffer_data_0[927:920];
        layer4[51][31:24] = buffer_data_0[935:928];
        layer4[51][39:32] = buffer_data_0[943:936];
        layer0[52][7:0] = buffer_data_4[919:912];
        layer0[52][15:8] = buffer_data_4[927:920];
        layer0[52][23:16] = buffer_data_4[935:928];
        layer0[52][31:24] = buffer_data_4[943:936];
        layer0[52][39:32] = buffer_data_4[951:944];
        layer1[52][7:0] = buffer_data_3[919:912];
        layer1[52][15:8] = buffer_data_3[927:920];
        layer1[52][23:16] = buffer_data_3[935:928];
        layer1[52][31:24] = buffer_data_3[943:936];
        layer1[52][39:32] = buffer_data_3[951:944];
        layer2[52][7:0] = buffer_data_2[919:912];
        layer2[52][15:8] = buffer_data_2[927:920];
        layer2[52][23:16] = buffer_data_2[935:928];
        layer2[52][31:24] = buffer_data_2[943:936];
        layer2[52][39:32] = buffer_data_2[951:944];
        layer3[52][7:0] = buffer_data_1[919:912];
        layer3[52][15:8] = buffer_data_1[927:920];
        layer3[52][23:16] = buffer_data_1[935:928];
        layer3[52][31:24] = buffer_data_1[943:936];
        layer3[52][39:32] = buffer_data_1[951:944];
        layer4[52][7:0] = buffer_data_0[919:912];
        layer4[52][15:8] = buffer_data_0[927:920];
        layer4[52][23:16] = buffer_data_0[935:928];
        layer4[52][31:24] = buffer_data_0[943:936];
        layer4[52][39:32] = buffer_data_0[951:944];
        layer0[53][7:0] = buffer_data_4[927:920];
        layer0[53][15:8] = buffer_data_4[935:928];
        layer0[53][23:16] = buffer_data_4[943:936];
        layer0[53][31:24] = buffer_data_4[951:944];
        layer0[53][39:32] = buffer_data_4[959:952];
        layer1[53][7:0] = buffer_data_3[927:920];
        layer1[53][15:8] = buffer_data_3[935:928];
        layer1[53][23:16] = buffer_data_3[943:936];
        layer1[53][31:24] = buffer_data_3[951:944];
        layer1[53][39:32] = buffer_data_3[959:952];
        layer2[53][7:0] = buffer_data_2[927:920];
        layer2[53][15:8] = buffer_data_2[935:928];
        layer2[53][23:16] = buffer_data_2[943:936];
        layer2[53][31:24] = buffer_data_2[951:944];
        layer2[53][39:32] = buffer_data_2[959:952];
        layer3[53][7:0] = buffer_data_1[927:920];
        layer3[53][15:8] = buffer_data_1[935:928];
        layer3[53][23:16] = buffer_data_1[943:936];
        layer3[53][31:24] = buffer_data_1[951:944];
        layer3[53][39:32] = buffer_data_1[959:952];
        layer4[53][7:0] = buffer_data_0[927:920];
        layer4[53][15:8] = buffer_data_0[935:928];
        layer4[53][23:16] = buffer_data_0[943:936];
        layer4[53][31:24] = buffer_data_0[951:944];
        layer4[53][39:32] = buffer_data_0[959:952];
        layer0[54][7:0] = buffer_data_4[935:928];
        layer0[54][15:8] = buffer_data_4[943:936];
        layer0[54][23:16] = buffer_data_4[951:944];
        layer0[54][31:24] = buffer_data_4[959:952];
        layer0[54][39:32] = buffer_data_4[967:960];
        layer1[54][7:0] = buffer_data_3[935:928];
        layer1[54][15:8] = buffer_data_3[943:936];
        layer1[54][23:16] = buffer_data_3[951:944];
        layer1[54][31:24] = buffer_data_3[959:952];
        layer1[54][39:32] = buffer_data_3[967:960];
        layer2[54][7:0] = buffer_data_2[935:928];
        layer2[54][15:8] = buffer_data_2[943:936];
        layer2[54][23:16] = buffer_data_2[951:944];
        layer2[54][31:24] = buffer_data_2[959:952];
        layer2[54][39:32] = buffer_data_2[967:960];
        layer3[54][7:0] = buffer_data_1[935:928];
        layer3[54][15:8] = buffer_data_1[943:936];
        layer3[54][23:16] = buffer_data_1[951:944];
        layer3[54][31:24] = buffer_data_1[959:952];
        layer3[54][39:32] = buffer_data_1[967:960];
        layer4[54][7:0] = buffer_data_0[935:928];
        layer4[54][15:8] = buffer_data_0[943:936];
        layer4[54][23:16] = buffer_data_0[951:944];
        layer4[54][31:24] = buffer_data_0[959:952];
        layer4[54][39:32] = buffer_data_0[967:960];
        layer0[55][7:0] = buffer_data_4[943:936];
        layer0[55][15:8] = buffer_data_4[951:944];
        layer0[55][23:16] = buffer_data_4[959:952];
        layer0[55][31:24] = buffer_data_4[967:960];
        layer0[55][39:32] = buffer_data_4[975:968];
        layer1[55][7:0] = buffer_data_3[943:936];
        layer1[55][15:8] = buffer_data_3[951:944];
        layer1[55][23:16] = buffer_data_3[959:952];
        layer1[55][31:24] = buffer_data_3[967:960];
        layer1[55][39:32] = buffer_data_3[975:968];
        layer2[55][7:0] = buffer_data_2[943:936];
        layer2[55][15:8] = buffer_data_2[951:944];
        layer2[55][23:16] = buffer_data_2[959:952];
        layer2[55][31:24] = buffer_data_2[967:960];
        layer2[55][39:32] = buffer_data_2[975:968];
        layer3[55][7:0] = buffer_data_1[943:936];
        layer3[55][15:8] = buffer_data_1[951:944];
        layer3[55][23:16] = buffer_data_1[959:952];
        layer3[55][31:24] = buffer_data_1[967:960];
        layer3[55][39:32] = buffer_data_1[975:968];
        layer4[55][7:0] = buffer_data_0[943:936];
        layer4[55][15:8] = buffer_data_0[951:944];
        layer4[55][23:16] = buffer_data_0[959:952];
        layer4[55][31:24] = buffer_data_0[967:960];
        layer4[55][39:32] = buffer_data_0[975:968];
        layer0[56][7:0] = buffer_data_4[951:944];
        layer0[56][15:8] = buffer_data_4[959:952];
        layer0[56][23:16] = buffer_data_4[967:960];
        layer0[56][31:24] = buffer_data_4[975:968];
        layer0[56][39:32] = buffer_data_4[983:976];
        layer1[56][7:0] = buffer_data_3[951:944];
        layer1[56][15:8] = buffer_data_3[959:952];
        layer1[56][23:16] = buffer_data_3[967:960];
        layer1[56][31:24] = buffer_data_3[975:968];
        layer1[56][39:32] = buffer_data_3[983:976];
        layer2[56][7:0] = buffer_data_2[951:944];
        layer2[56][15:8] = buffer_data_2[959:952];
        layer2[56][23:16] = buffer_data_2[967:960];
        layer2[56][31:24] = buffer_data_2[975:968];
        layer2[56][39:32] = buffer_data_2[983:976];
        layer3[56][7:0] = buffer_data_1[951:944];
        layer3[56][15:8] = buffer_data_1[959:952];
        layer3[56][23:16] = buffer_data_1[967:960];
        layer3[56][31:24] = buffer_data_1[975:968];
        layer3[56][39:32] = buffer_data_1[983:976];
        layer4[56][7:0] = buffer_data_0[951:944];
        layer4[56][15:8] = buffer_data_0[959:952];
        layer4[56][23:16] = buffer_data_0[967:960];
        layer4[56][31:24] = buffer_data_0[975:968];
        layer4[56][39:32] = buffer_data_0[983:976];
        layer0[57][7:0] = buffer_data_4[959:952];
        layer0[57][15:8] = buffer_data_4[967:960];
        layer0[57][23:16] = buffer_data_4[975:968];
        layer0[57][31:24] = buffer_data_4[983:976];
        layer0[57][39:32] = buffer_data_4[991:984];
        layer1[57][7:0] = buffer_data_3[959:952];
        layer1[57][15:8] = buffer_data_3[967:960];
        layer1[57][23:16] = buffer_data_3[975:968];
        layer1[57][31:24] = buffer_data_3[983:976];
        layer1[57][39:32] = buffer_data_3[991:984];
        layer2[57][7:0] = buffer_data_2[959:952];
        layer2[57][15:8] = buffer_data_2[967:960];
        layer2[57][23:16] = buffer_data_2[975:968];
        layer2[57][31:24] = buffer_data_2[983:976];
        layer2[57][39:32] = buffer_data_2[991:984];
        layer3[57][7:0] = buffer_data_1[959:952];
        layer3[57][15:8] = buffer_data_1[967:960];
        layer3[57][23:16] = buffer_data_1[975:968];
        layer3[57][31:24] = buffer_data_1[983:976];
        layer3[57][39:32] = buffer_data_1[991:984];
        layer4[57][7:0] = buffer_data_0[959:952];
        layer4[57][15:8] = buffer_data_0[967:960];
        layer4[57][23:16] = buffer_data_0[975:968];
        layer4[57][31:24] = buffer_data_0[983:976];
        layer4[57][39:32] = buffer_data_0[991:984];
        layer0[58][7:0] = buffer_data_4[967:960];
        layer0[58][15:8] = buffer_data_4[975:968];
        layer0[58][23:16] = buffer_data_4[983:976];
        layer0[58][31:24] = buffer_data_4[991:984];
        layer0[58][39:32] = buffer_data_4[999:992];
        layer1[58][7:0] = buffer_data_3[967:960];
        layer1[58][15:8] = buffer_data_3[975:968];
        layer1[58][23:16] = buffer_data_3[983:976];
        layer1[58][31:24] = buffer_data_3[991:984];
        layer1[58][39:32] = buffer_data_3[999:992];
        layer2[58][7:0] = buffer_data_2[967:960];
        layer2[58][15:8] = buffer_data_2[975:968];
        layer2[58][23:16] = buffer_data_2[983:976];
        layer2[58][31:24] = buffer_data_2[991:984];
        layer2[58][39:32] = buffer_data_2[999:992];
        layer3[58][7:0] = buffer_data_1[967:960];
        layer3[58][15:8] = buffer_data_1[975:968];
        layer3[58][23:16] = buffer_data_1[983:976];
        layer3[58][31:24] = buffer_data_1[991:984];
        layer3[58][39:32] = buffer_data_1[999:992];
        layer4[58][7:0] = buffer_data_0[967:960];
        layer4[58][15:8] = buffer_data_0[975:968];
        layer4[58][23:16] = buffer_data_0[983:976];
        layer4[58][31:24] = buffer_data_0[991:984];
        layer4[58][39:32] = buffer_data_0[999:992];
        layer0[59][7:0] = buffer_data_4[975:968];
        layer0[59][15:8] = buffer_data_4[983:976];
        layer0[59][23:16] = buffer_data_4[991:984];
        layer0[59][31:24] = buffer_data_4[999:992];
        layer0[59][39:32] = buffer_data_4[1007:1000];
        layer1[59][7:0] = buffer_data_3[975:968];
        layer1[59][15:8] = buffer_data_3[983:976];
        layer1[59][23:16] = buffer_data_3[991:984];
        layer1[59][31:24] = buffer_data_3[999:992];
        layer1[59][39:32] = buffer_data_3[1007:1000];
        layer2[59][7:0] = buffer_data_2[975:968];
        layer2[59][15:8] = buffer_data_2[983:976];
        layer2[59][23:16] = buffer_data_2[991:984];
        layer2[59][31:24] = buffer_data_2[999:992];
        layer2[59][39:32] = buffer_data_2[1007:1000];
        layer3[59][7:0] = buffer_data_1[975:968];
        layer3[59][15:8] = buffer_data_1[983:976];
        layer3[59][23:16] = buffer_data_1[991:984];
        layer3[59][31:24] = buffer_data_1[999:992];
        layer3[59][39:32] = buffer_data_1[1007:1000];
        layer4[59][7:0] = buffer_data_0[975:968];
        layer4[59][15:8] = buffer_data_0[983:976];
        layer4[59][23:16] = buffer_data_0[991:984];
        layer4[59][31:24] = buffer_data_0[999:992];
        layer4[59][39:32] = buffer_data_0[1007:1000];
        layer0[60][7:0] = buffer_data_4[983:976];
        layer0[60][15:8] = buffer_data_4[991:984];
        layer0[60][23:16] = buffer_data_4[999:992];
        layer0[60][31:24] = buffer_data_4[1007:1000];
        layer0[60][39:32] = buffer_data_4[1015:1008];
        layer1[60][7:0] = buffer_data_3[983:976];
        layer1[60][15:8] = buffer_data_3[991:984];
        layer1[60][23:16] = buffer_data_3[999:992];
        layer1[60][31:24] = buffer_data_3[1007:1000];
        layer1[60][39:32] = buffer_data_3[1015:1008];
        layer2[60][7:0] = buffer_data_2[983:976];
        layer2[60][15:8] = buffer_data_2[991:984];
        layer2[60][23:16] = buffer_data_2[999:992];
        layer2[60][31:24] = buffer_data_2[1007:1000];
        layer2[60][39:32] = buffer_data_2[1015:1008];
        layer3[60][7:0] = buffer_data_1[983:976];
        layer3[60][15:8] = buffer_data_1[991:984];
        layer3[60][23:16] = buffer_data_1[999:992];
        layer3[60][31:24] = buffer_data_1[1007:1000];
        layer3[60][39:32] = buffer_data_1[1015:1008];
        layer4[60][7:0] = buffer_data_0[983:976];
        layer4[60][15:8] = buffer_data_0[991:984];
        layer4[60][23:16] = buffer_data_0[999:992];
        layer4[60][31:24] = buffer_data_0[1007:1000];
        layer4[60][39:32] = buffer_data_0[1015:1008];
        layer0[61][7:0] = buffer_data_4[991:984];
        layer0[61][15:8] = buffer_data_4[999:992];
        layer0[61][23:16] = buffer_data_4[1007:1000];
        layer0[61][31:24] = buffer_data_4[1015:1008];
        layer0[61][39:32] = buffer_data_4[1023:1016];
        layer1[61][7:0] = buffer_data_3[991:984];
        layer1[61][15:8] = buffer_data_3[999:992];
        layer1[61][23:16] = buffer_data_3[1007:1000];
        layer1[61][31:24] = buffer_data_3[1015:1008];
        layer1[61][39:32] = buffer_data_3[1023:1016];
        layer2[61][7:0] = buffer_data_2[991:984];
        layer2[61][15:8] = buffer_data_2[999:992];
        layer2[61][23:16] = buffer_data_2[1007:1000];
        layer2[61][31:24] = buffer_data_2[1015:1008];
        layer2[61][39:32] = buffer_data_2[1023:1016];
        layer3[61][7:0] = buffer_data_1[991:984];
        layer3[61][15:8] = buffer_data_1[999:992];
        layer3[61][23:16] = buffer_data_1[1007:1000];
        layer3[61][31:24] = buffer_data_1[1015:1008];
        layer3[61][39:32] = buffer_data_1[1023:1016];
        layer4[61][7:0] = buffer_data_0[991:984];
        layer4[61][15:8] = buffer_data_0[999:992];
        layer4[61][23:16] = buffer_data_0[1007:1000];
        layer4[61][31:24] = buffer_data_0[1015:1008];
        layer4[61][39:32] = buffer_data_0[1023:1016];
        layer0[62][7:0] = buffer_data_4[999:992];
        layer0[62][15:8] = buffer_data_4[1007:1000];
        layer0[62][23:16] = buffer_data_4[1015:1008];
        layer0[62][31:24] = buffer_data_4[1023:1016];
        layer0[62][39:32] = buffer_data_4[1031:1024];
        layer1[62][7:0] = buffer_data_3[999:992];
        layer1[62][15:8] = buffer_data_3[1007:1000];
        layer1[62][23:16] = buffer_data_3[1015:1008];
        layer1[62][31:24] = buffer_data_3[1023:1016];
        layer1[62][39:32] = buffer_data_3[1031:1024];
        layer2[62][7:0] = buffer_data_2[999:992];
        layer2[62][15:8] = buffer_data_2[1007:1000];
        layer2[62][23:16] = buffer_data_2[1015:1008];
        layer2[62][31:24] = buffer_data_2[1023:1016];
        layer2[62][39:32] = buffer_data_2[1031:1024];
        layer3[62][7:0] = buffer_data_1[999:992];
        layer3[62][15:8] = buffer_data_1[1007:1000];
        layer3[62][23:16] = buffer_data_1[1015:1008];
        layer3[62][31:24] = buffer_data_1[1023:1016];
        layer3[62][39:32] = buffer_data_1[1031:1024];
        layer4[62][7:0] = buffer_data_0[999:992];
        layer4[62][15:8] = buffer_data_0[1007:1000];
        layer4[62][23:16] = buffer_data_0[1015:1008];
        layer4[62][31:24] = buffer_data_0[1023:1016];
        layer4[62][39:32] = buffer_data_0[1031:1024];
        layer0[63][7:0] = buffer_data_4[1007:1000];
        layer0[63][15:8] = buffer_data_4[1015:1008];
        layer0[63][23:16] = buffer_data_4[1023:1016];
        layer0[63][31:24] = buffer_data_4[1031:1024];
        layer0[63][39:32] = buffer_data_4[1039:1032];
        layer1[63][7:0] = buffer_data_3[1007:1000];
        layer1[63][15:8] = buffer_data_3[1015:1008];
        layer1[63][23:16] = buffer_data_3[1023:1016];
        layer1[63][31:24] = buffer_data_3[1031:1024];
        layer1[63][39:32] = buffer_data_3[1039:1032];
        layer2[63][7:0] = buffer_data_2[1007:1000];
        layer2[63][15:8] = buffer_data_2[1015:1008];
        layer2[63][23:16] = buffer_data_2[1023:1016];
        layer2[63][31:24] = buffer_data_2[1031:1024];
        layer2[63][39:32] = buffer_data_2[1039:1032];
        layer3[63][7:0] = buffer_data_1[1007:1000];
        layer3[63][15:8] = buffer_data_1[1015:1008];
        layer3[63][23:16] = buffer_data_1[1023:1016];
        layer3[63][31:24] = buffer_data_1[1031:1024];
        layer3[63][39:32] = buffer_data_1[1039:1032];
        layer4[63][7:0] = buffer_data_0[1007:1000];
        layer4[63][15:8] = buffer_data_0[1015:1008];
        layer4[63][23:16] = buffer_data_0[1023:1016];
        layer4[63][31:24] = buffer_data_0[1031:1024];
        layer4[63][39:32] = buffer_data_0[1039:1032];
    end
    ST_GAUSSIAN_2: begin
        layer0[0][7:0] = buffer_data_4[1015:1008];
        layer0[0][15:8] = buffer_data_4[1023:1016];
        layer0[0][23:16] = buffer_data_4[1031:1024];
        layer0[0][31:24] = buffer_data_4[1039:1032];
        layer0[0][39:32] = buffer_data_4[1047:1040];
        layer1[0][7:0] = buffer_data_3[1015:1008];
        layer1[0][15:8] = buffer_data_3[1023:1016];
        layer1[0][23:16] = buffer_data_3[1031:1024];
        layer1[0][31:24] = buffer_data_3[1039:1032];
        layer1[0][39:32] = buffer_data_3[1047:1040];
        layer2[0][7:0] = buffer_data_2[1015:1008];
        layer2[0][15:8] = buffer_data_2[1023:1016];
        layer2[0][23:16] = buffer_data_2[1031:1024];
        layer2[0][31:24] = buffer_data_2[1039:1032];
        layer2[0][39:32] = buffer_data_2[1047:1040];
        layer3[0][7:0] = buffer_data_1[1015:1008];
        layer3[0][15:8] = buffer_data_1[1023:1016];
        layer3[0][23:16] = buffer_data_1[1031:1024];
        layer3[0][31:24] = buffer_data_1[1039:1032];
        layer3[0][39:32] = buffer_data_1[1047:1040];
        layer4[0][7:0] = buffer_data_0[1015:1008];
        layer4[0][15:8] = buffer_data_0[1023:1016];
        layer4[0][23:16] = buffer_data_0[1031:1024];
        layer4[0][31:24] = buffer_data_0[1039:1032];
        layer4[0][39:32] = buffer_data_0[1047:1040];
        layer0[1][7:0] = buffer_data_4[1023:1016];
        layer0[1][15:8] = buffer_data_4[1031:1024];
        layer0[1][23:16] = buffer_data_4[1039:1032];
        layer0[1][31:24] = buffer_data_4[1047:1040];
        layer0[1][39:32] = buffer_data_4[1055:1048];
        layer1[1][7:0] = buffer_data_3[1023:1016];
        layer1[1][15:8] = buffer_data_3[1031:1024];
        layer1[1][23:16] = buffer_data_3[1039:1032];
        layer1[1][31:24] = buffer_data_3[1047:1040];
        layer1[1][39:32] = buffer_data_3[1055:1048];
        layer2[1][7:0] = buffer_data_2[1023:1016];
        layer2[1][15:8] = buffer_data_2[1031:1024];
        layer2[1][23:16] = buffer_data_2[1039:1032];
        layer2[1][31:24] = buffer_data_2[1047:1040];
        layer2[1][39:32] = buffer_data_2[1055:1048];
        layer3[1][7:0] = buffer_data_1[1023:1016];
        layer3[1][15:8] = buffer_data_1[1031:1024];
        layer3[1][23:16] = buffer_data_1[1039:1032];
        layer3[1][31:24] = buffer_data_1[1047:1040];
        layer3[1][39:32] = buffer_data_1[1055:1048];
        layer4[1][7:0] = buffer_data_0[1023:1016];
        layer4[1][15:8] = buffer_data_0[1031:1024];
        layer4[1][23:16] = buffer_data_0[1039:1032];
        layer4[1][31:24] = buffer_data_0[1047:1040];
        layer4[1][39:32] = buffer_data_0[1055:1048];
        layer0[2][7:0] = buffer_data_4[1031:1024];
        layer0[2][15:8] = buffer_data_4[1039:1032];
        layer0[2][23:16] = buffer_data_4[1047:1040];
        layer0[2][31:24] = buffer_data_4[1055:1048];
        layer0[2][39:32] = buffer_data_4[1063:1056];
        layer1[2][7:0] = buffer_data_3[1031:1024];
        layer1[2][15:8] = buffer_data_3[1039:1032];
        layer1[2][23:16] = buffer_data_3[1047:1040];
        layer1[2][31:24] = buffer_data_3[1055:1048];
        layer1[2][39:32] = buffer_data_3[1063:1056];
        layer2[2][7:0] = buffer_data_2[1031:1024];
        layer2[2][15:8] = buffer_data_2[1039:1032];
        layer2[2][23:16] = buffer_data_2[1047:1040];
        layer2[2][31:24] = buffer_data_2[1055:1048];
        layer2[2][39:32] = buffer_data_2[1063:1056];
        layer3[2][7:0] = buffer_data_1[1031:1024];
        layer3[2][15:8] = buffer_data_1[1039:1032];
        layer3[2][23:16] = buffer_data_1[1047:1040];
        layer3[2][31:24] = buffer_data_1[1055:1048];
        layer3[2][39:32] = buffer_data_1[1063:1056];
        layer4[2][7:0] = buffer_data_0[1031:1024];
        layer4[2][15:8] = buffer_data_0[1039:1032];
        layer4[2][23:16] = buffer_data_0[1047:1040];
        layer4[2][31:24] = buffer_data_0[1055:1048];
        layer4[2][39:32] = buffer_data_0[1063:1056];
        layer0[3][7:0] = buffer_data_4[1039:1032];
        layer0[3][15:8] = buffer_data_4[1047:1040];
        layer0[3][23:16] = buffer_data_4[1055:1048];
        layer0[3][31:24] = buffer_data_4[1063:1056];
        layer0[3][39:32] = buffer_data_4[1071:1064];
        layer1[3][7:0] = buffer_data_3[1039:1032];
        layer1[3][15:8] = buffer_data_3[1047:1040];
        layer1[3][23:16] = buffer_data_3[1055:1048];
        layer1[3][31:24] = buffer_data_3[1063:1056];
        layer1[3][39:32] = buffer_data_3[1071:1064];
        layer2[3][7:0] = buffer_data_2[1039:1032];
        layer2[3][15:8] = buffer_data_2[1047:1040];
        layer2[3][23:16] = buffer_data_2[1055:1048];
        layer2[3][31:24] = buffer_data_2[1063:1056];
        layer2[3][39:32] = buffer_data_2[1071:1064];
        layer3[3][7:0] = buffer_data_1[1039:1032];
        layer3[3][15:8] = buffer_data_1[1047:1040];
        layer3[3][23:16] = buffer_data_1[1055:1048];
        layer3[3][31:24] = buffer_data_1[1063:1056];
        layer3[3][39:32] = buffer_data_1[1071:1064];
        layer4[3][7:0] = buffer_data_0[1039:1032];
        layer4[3][15:8] = buffer_data_0[1047:1040];
        layer4[3][23:16] = buffer_data_0[1055:1048];
        layer4[3][31:24] = buffer_data_0[1063:1056];
        layer4[3][39:32] = buffer_data_0[1071:1064];
        layer0[4][7:0] = buffer_data_4[1047:1040];
        layer0[4][15:8] = buffer_data_4[1055:1048];
        layer0[4][23:16] = buffer_data_4[1063:1056];
        layer0[4][31:24] = buffer_data_4[1071:1064];
        layer0[4][39:32] = buffer_data_4[1079:1072];
        layer1[4][7:0] = buffer_data_3[1047:1040];
        layer1[4][15:8] = buffer_data_3[1055:1048];
        layer1[4][23:16] = buffer_data_3[1063:1056];
        layer1[4][31:24] = buffer_data_3[1071:1064];
        layer1[4][39:32] = buffer_data_3[1079:1072];
        layer2[4][7:0] = buffer_data_2[1047:1040];
        layer2[4][15:8] = buffer_data_2[1055:1048];
        layer2[4][23:16] = buffer_data_2[1063:1056];
        layer2[4][31:24] = buffer_data_2[1071:1064];
        layer2[4][39:32] = buffer_data_2[1079:1072];
        layer3[4][7:0] = buffer_data_1[1047:1040];
        layer3[4][15:8] = buffer_data_1[1055:1048];
        layer3[4][23:16] = buffer_data_1[1063:1056];
        layer3[4][31:24] = buffer_data_1[1071:1064];
        layer3[4][39:32] = buffer_data_1[1079:1072];
        layer4[4][7:0] = buffer_data_0[1047:1040];
        layer4[4][15:8] = buffer_data_0[1055:1048];
        layer4[4][23:16] = buffer_data_0[1063:1056];
        layer4[4][31:24] = buffer_data_0[1071:1064];
        layer4[4][39:32] = buffer_data_0[1079:1072];
        layer0[5][7:0] = buffer_data_4[1055:1048];
        layer0[5][15:8] = buffer_data_4[1063:1056];
        layer0[5][23:16] = buffer_data_4[1071:1064];
        layer0[5][31:24] = buffer_data_4[1079:1072];
        layer0[5][39:32] = buffer_data_4[1087:1080];
        layer1[5][7:0] = buffer_data_3[1055:1048];
        layer1[5][15:8] = buffer_data_3[1063:1056];
        layer1[5][23:16] = buffer_data_3[1071:1064];
        layer1[5][31:24] = buffer_data_3[1079:1072];
        layer1[5][39:32] = buffer_data_3[1087:1080];
        layer2[5][7:0] = buffer_data_2[1055:1048];
        layer2[5][15:8] = buffer_data_2[1063:1056];
        layer2[5][23:16] = buffer_data_2[1071:1064];
        layer2[5][31:24] = buffer_data_2[1079:1072];
        layer2[5][39:32] = buffer_data_2[1087:1080];
        layer3[5][7:0] = buffer_data_1[1055:1048];
        layer3[5][15:8] = buffer_data_1[1063:1056];
        layer3[5][23:16] = buffer_data_1[1071:1064];
        layer3[5][31:24] = buffer_data_1[1079:1072];
        layer3[5][39:32] = buffer_data_1[1087:1080];
        layer4[5][7:0] = buffer_data_0[1055:1048];
        layer4[5][15:8] = buffer_data_0[1063:1056];
        layer4[5][23:16] = buffer_data_0[1071:1064];
        layer4[5][31:24] = buffer_data_0[1079:1072];
        layer4[5][39:32] = buffer_data_0[1087:1080];
        layer0[6][7:0] = buffer_data_4[1063:1056];
        layer0[6][15:8] = buffer_data_4[1071:1064];
        layer0[6][23:16] = buffer_data_4[1079:1072];
        layer0[6][31:24] = buffer_data_4[1087:1080];
        layer0[6][39:32] = buffer_data_4[1095:1088];
        layer1[6][7:0] = buffer_data_3[1063:1056];
        layer1[6][15:8] = buffer_data_3[1071:1064];
        layer1[6][23:16] = buffer_data_3[1079:1072];
        layer1[6][31:24] = buffer_data_3[1087:1080];
        layer1[6][39:32] = buffer_data_3[1095:1088];
        layer2[6][7:0] = buffer_data_2[1063:1056];
        layer2[6][15:8] = buffer_data_2[1071:1064];
        layer2[6][23:16] = buffer_data_2[1079:1072];
        layer2[6][31:24] = buffer_data_2[1087:1080];
        layer2[6][39:32] = buffer_data_2[1095:1088];
        layer3[6][7:0] = buffer_data_1[1063:1056];
        layer3[6][15:8] = buffer_data_1[1071:1064];
        layer3[6][23:16] = buffer_data_1[1079:1072];
        layer3[6][31:24] = buffer_data_1[1087:1080];
        layer3[6][39:32] = buffer_data_1[1095:1088];
        layer4[6][7:0] = buffer_data_0[1063:1056];
        layer4[6][15:8] = buffer_data_0[1071:1064];
        layer4[6][23:16] = buffer_data_0[1079:1072];
        layer4[6][31:24] = buffer_data_0[1087:1080];
        layer4[6][39:32] = buffer_data_0[1095:1088];
        layer0[7][7:0] = buffer_data_4[1071:1064];
        layer0[7][15:8] = buffer_data_4[1079:1072];
        layer0[7][23:16] = buffer_data_4[1087:1080];
        layer0[7][31:24] = buffer_data_4[1095:1088];
        layer0[7][39:32] = buffer_data_4[1103:1096];
        layer1[7][7:0] = buffer_data_3[1071:1064];
        layer1[7][15:8] = buffer_data_3[1079:1072];
        layer1[7][23:16] = buffer_data_3[1087:1080];
        layer1[7][31:24] = buffer_data_3[1095:1088];
        layer1[7][39:32] = buffer_data_3[1103:1096];
        layer2[7][7:0] = buffer_data_2[1071:1064];
        layer2[7][15:8] = buffer_data_2[1079:1072];
        layer2[7][23:16] = buffer_data_2[1087:1080];
        layer2[7][31:24] = buffer_data_2[1095:1088];
        layer2[7][39:32] = buffer_data_2[1103:1096];
        layer3[7][7:0] = buffer_data_1[1071:1064];
        layer3[7][15:8] = buffer_data_1[1079:1072];
        layer3[7][23:16] = buffer_data_1[1087:1080];
        layer3[7][31:24] = buffer_data_1[1095:1088];
        layer3[7][39:32] = buffer_data_1[1103:1096];
        layer4[7][7:0] = buffer_data_0[1071:1064];
        layer4[7][15:8] = buffer_data_0[1079:1072];
        layer4[7][23:16] = buffer_data_0[1087:1080];
        layer4[7][31:24] = buffer_data_0[1095:1088];
        layer4[7][39:32] = buffer_data_0[1103:1096];
        layer0[8][7:0] = buffer_data_4[1079:1072];
        layer0[8][15:8] = buffer_data_4[1087:1080];
        layer0[8][23:16] = buffer_data_4[1095:1088];
        layer0[8][31:24] = buffer_data_4[1103:1096];
        layer0[8][39:32] = buffer_data_4[1111:1104];
        layer1[8][7:0] = buffer_data_3[1079:1072];
        layer1[8][15:8] = buffer_data_3[1087:1080];
        layer1[8][23:16] = buffer_data_3[1095:1088];
        layer1[8][31:24] = buffer_data_3[1103:1096];
        layer1[8][39:32] = buffer_data_3[1111:1104];
        layer2[8][7:0] = buffer_data_2[1079:1072];
        layer2[8][15:8] = buffer_data_2[1087:1080];
        layer2[8][23:16] = buffer_data_2[1095:1088];
        layer2[8][31:24] = buffer_data_2[1103:1096];
        layer2[8][39:32] = buffer_data_2[1111:1104];
        layer3[8][7:0] = buffer_data_1[1079:1072];
        layer3[8][15:8] = buffer_data_1[1087:1080];
        layer3[8][23:16] = buffer_data_1[1095:1088];
        layer3[8][31:24] = buffer_data_1[1103:1096];
        layer3[8][39:32] = buffer_data_1[1111:1104];
        layer4[8][7:0] = buffer_data_0[1079:1072];
        layer4[8][15:8] = buffer_data_0[1087:1080];
        layer4[8][23:16] = buffer_data_0[1095:1088];
        layer4[8][31:24] = buffer_data_0[1103:1096];
        layer4[8][39:32] = buffer_data_0[1111:1104];
        layer0[9][7:0] = buffer_data_4[1087:1080];
        layer0[9][15:8] = buffer_data_4[1095:1088];
        layer0[9][23:16] = buffer_data_4[1103:1096];
        layer0[9][31:24] = buffer_data_4[1111:1104];
        layer0[9][39:32] = buffer_data_4[1119:1112];
        layer1[9][7:0] = buffer_data_3[1087:1080];
        layer1[9][15:8] = buffer_data_3[1095:1088];
        layer1[9][23:16] = buffer_data_3[1103:1096];
        layer1[9][31:24] = buffer_data_3[1111:1104];
        layer1[9][39:32] = buffer_data_3[1119:1112];
        layer2[9][7:0] = buffer_data_2[1087:1080];
        layer2[9][15:8] = buffer_data_2[1095:1088];
        layer2[9][23:16] = buffer_data_2[1103:1096];
        layer2[9][31:24] = buffer_data_2[1111:1104];
        layer2[9][39:32] = buffer_data_2[1119:1112];
        layer3[9][7:0] = buffer_data_1[1087:1080];
        layer3[9][15:8] = buffer_data_1[1095:1088];
        layer3[9][23:16] = buffer_data_1[1103:1096];
        layer3[9][31:24] = buffer_data_1[1111:1104];
        layer3[9][39:32] = buffer_data_1[1119:1112];
        layer4[9][7:0] = buffer_data_0[1087:1080];
        layer4[9][15:8] = buffer_data_0[1095:1088];
        layer4[9][23:16] = buffer_data_0[1103:1096];
        layer4[9][31:24] = buffer_data_0[1111:1104];
        layer4[9][39:32] = buffer_data_0[1119:1112];
        layer0[10][7:0] = buffer_data_4[1095:1088];
        layer0[10][15:8] = buffer_data_4[1103:1096];
        layer0[10][23:16] = buffer_data_4[1111:1104];
        layer0[10][31:24] = buffer_data_4[1119:1112];
        layer0[10][39:32] = buffer_data_4[1127:1120];
        layer1[10][7:0] = buffer_data_3[1095:1088];
        layer1[10][15:8] = buffer_data_3[1103:1096];
        layer1[10][23:16] = buffer_data_3[1111:1104];
        layer1[10][31:24] = buffer_data_3[1119:1112];
        layer1[10][39:32] = buffer_data_3[1127:1120];
        layer2[10][7:0] = buffer_data_2[1095:1088];
        layer2[10][15:8] = buffer_data_2[1103:1096];
        layer2[10][23:16] = buffer_data_2[1111:1104];
        layer2[10][31:24] = buffer_data_2[1119:1112];
        layer2[10][39:32] = buffer_data_2[1127:1120];
        layer3[10][7:0] = buffer_data_1[1095:1088];
        layer3[10][15:8] = buffer_data_1[1103:1096];
        layer3[10][23:16] = buffer_data_1[1111:1104];
        layer3[10][31:24] = buffer_data_1[1119:1112];
        layer3[10][39:32] = buffer_data_1[1127:1120];
        layer4[10][7:0] = buffer_data_0[1095:1088];
        layer4[10][15:8] = buffer_data_0[1103:1096];
        layer4[10][23:16] = buffer_data_0[1111:1104];
        layer4[10][31:24] = buffer_data_0[1119:1112];
        layer4[10][39:32] = buffer_data_0[1127:1120];
        layer0[11][7:0] = buffer_data_4[1103:1096];
        layer0[11][15:8] = buffer_data_4[1111:1104];
        layer0[11][23:16] = buffer_data_4[1119:1112];
        layer0[11][31:24] = buffer_data_4[1127:1120];
        layer0[11][39:32] = buffer_data_4[1135:1128];
        layer1[11][7:0] = buffer_data_3[1103:1096];
        layer1[11][15:8] = buffer_data_3[1111:1104];
        layer1[11][23:16] = buffer_data_3[1119:1112];
        layer1[11][31:24] = buffer_data_3[1127:1120];
        layer1[11][39:32] = buffer_data_3[1135:1128];
        layer2[11][7:0] = buffer_data_2[1103:1096];
        layer2[11][15:8] = buffer_data_2[1111:1104];
        layer2[11][23:16] = buffer_data_2[1119:1112];
        layer2[11][31:24] = buffer_data_2[1127:1120];
        layer2[11][39:32] = buffer_data_2[1135:1128];
        layer3[11][7:0] = buffer_data_1[1103:1096];
        layer3[11][15:8] = buffer_data_1[1111:1104];
        layer3[11][23:16] = buffer_data_1[1119:1112];
        layer3[11][31:24] = buffer_data_1[1127:1120];
        layer3[11][39:32] = buffer_data_1[1135:1128];
        layer4[11][7:0] = buffer_data_0[1103:1096];
        layer4[11][15:8] = buffer_data_0[1111:1104];
        layer4[11][23:16] = buffer_data_0[1119:1112];
        layer4[11][31:24] = buffer_data_0[1127:1120];
        layer4[11][39:32] = buffer_data_0[1135:1128];
        layer0[12][7:0] = buffer_data_4[1111:1104];
        layer0[12][15:8] = buffer_data_4[1119:1112];
        layer0[12][23:16] = buffer_data_4[1127:1120];
        layer0[12][31:24] = buffer_data_4[1135:1128];
        layer0[12][39:32] = buffer_data_4[1143:1136];
        layer1[12][7:0] = buffer_data_3[1111:1104];
        layer1[12][15:8] = buffer_data_3[1119:1112];
        layer1[12][23:16] = buffer_data_3[1127:1120];
        layer1[12][31:24] = buffer_data_3[1135:1128];
        layer1[12][39:32] = buffer_data_3[1143:1136];
        layer2[12][7:0] = buffer_data_2[1111:1104];
        layer2[12][15:8] = buffer_data_2[1119:1112];
        layer2[12][23:16] = buffer_data_2[1127:1120];
        layer2[12][31:24] = buffer_data_2[1135:1128];
        layer2[12][39:32] = buffer_data_2[1143:1136];
        layer3[12][7:0] = buffer_data_1[1111:1104];
        layer3[12][15:8] = buffer_data_1[1119:1112];
        layer3[12][23:16] = buffer_data_1[1127:1120];
        layer3[12][31:24] = buffer_data_1[1135:1128];
        layer3[12][39:32] = buffer_data_1[1143:1136];
        layer4[12][7:0] = buffer_data_0[1111:1104];
        layer4[12][15:8] = buffer_data_0[1119:1112];
        layer4[12][23:16] = buffer_data_0[1127:1120];
        layer4[12][31:24] = buffer_data_0[1135:1128];
        layer4[12][39:32] = buffer_data_0[1143:1136];
        layer0[13][7:0] = buffer_data_4[1119:1112];
        layer0[13][15:8] = buffer_data_4[1127:1120];
        layer0[13][23:16] = buffer_data_4[1135:1128];
        layer0[13][31:24] = buffer_data_4[1143:1136];
        layer0[13][39:32] = buffer_data_4[1151:1144];
        layer1[13][7:0] = buffer_data_3[1119:1112];
        layer1[13][15:8] = buffer_data_3[1127:1120];
        layer1[13][23:16] = buffer_data_3[1135:1128];
        layer1[13][31:24] = buffer_data_3[1143:1136];
        layer1[13][39:32] = buffer_data_3[1151:1144];
        layer2[13][7:0] = buffer_data_2[1119:1112];
        layer2[13][15:8] = buffer_data_2[1127:1120];
        layer2[13][23:16] = buffer_data_2[1135:1128];
        layer2[13][31:24] = buffer_data_2[1143:1136];
        layer2[13][39:32] = buffer_data_2[1151:1144];
        layer3[13][7:0] = buffer_data_1[1119:1112];
        layer3[13][15:8] = buffer_data_1[1127:1120];
        layer3[13][23:16] = buffer_data_1[1135:1128];
        layer3[13][31:24] = buffer_data_1[1143:1136];
        layer3[13][39:32] = buffer_data_1[1151:1144];
        layer4[13][7:0] = buffer_data_0[1119:1112];
        layer4[13][15:8] = buffer_data_0[1127:1120];
        layer4[13][23:16] = buffer_data_0[1135:1128];
        layer4[13][31:24] = buffer_data_0[1143:1136];
        layer4[13][39:32] = buffer_data_0[1151:1144];
        layer0[14][7:0] = buffer_data_4[1127:1120];
        layer0[14][15:8] = buffer_data_4[1135:1128];
        layer0[14][23:16] = buffer_data_4[1143:1136];
        layer0[14][31:24] = buffer_data_4[1151:1144];
        layer0[14][39:32] = buffer_data_4[1159:1152];
        layer1[14][7:0] = buffer_data_3[1127:1120];
        layer1[14][15:8] = buffer_data_3[1135:1128];
        layer1[14][23:16] = buffer_data_3[1143:1136];
        layer1[14][31:24] = buffer_data_3[1151:1144];
        layer1[14][39:32] = buffer_data_3[1159:1152];
        layer2[14][7:0] = buffer_data_2[1127:1120];
        layer2[14][15:8] = buffer_data_2[1135:1128];
        layer2[14][23:16] = buffer_data_2[1143:1136];
        layer2[14][31:24] = buffer_data_2[1151:1144];
        layer2[14][39:32] = buffer_data_2[1159:1152];
        layer3[14][7:0] = buffer_data_1[1127:1120];
        layer3[14][15:8] = buffer_data_1[1135:1128];
        layer3[14][23:16] = buffer_data_1[1143:1136];
        layer3[14][31:24] = buffer_data_1[1151:1144];
        layer3[14][39:32] = buffer_data_1[1159:1152];
        layer4[14][7:0] = buffer_data_0[1127:1120];
        layer4[14][15:8] = buffer_data_0[1135:1128];
        layer4[14][23:16] = buffer_data_0[1143:1136];
        layer4[14][31:24] = buffer_data_0[1151:1144];
        layer4[14][39:32] = buffer_data_0[1159:1152];
        layer0[15][7:0] = buffer_data_4[1135:1128];
        layer0[15][15:8] = buffer_data_4[1143:1136];
        layer0[15][23:16] = buffer_data_4[1151:1144];
        layer0[15][31:24] = buffer_data_4[1159:1152];
        layer0[15][39:32] = buffer_data_4[1167:1160];
        layer1[15][7:0] = buffer_data_3[1135:1128];
        layer1[15][15:8] = buffer_data_3[1143:1136];
        layer1[15][23:16] = buffer_data_3[1151:1144];
        layer1[15][31:24] = buffer_data_3[1159:1152];
        layer1[15][39:32] = buffer_data_3[1167:1160];
        layer2[15][7:0] = buffer_data_2[1135:1128];
        layer2[15][15:8] = buffer_data_2[1143:1136];
        layer2[15][23:16] = buffer_data_2[1151:1144];
        layer2[15][31:24] = buffer_data_2[1159:1152];
        layer2[15][39:32] = buffer_data_2[1167:1160];
        layer3[15][7:0] = buffer_data_1[1135:1128];
        layer3[15][15:8] = buffer_data_1[1143:1136];
        layer3[15][23:16] = buffer_data_1[1151:1144];
        layer3[15][31:24] = buffer_data_1[1159:1152];
        layer3[15][39:32] = buffer_data_1[1167:1160];
        layer4[15][7:0] = buffer_data_0[1135:1128];
        layer4[15][15:8] = buffer_data_0[1143:1136];
        layer4[15][23:16] = buffer_data_0[1151:1144];
        layer4[15][31:24] = buffer_data_0[1159:1152];
        layer4[15][39:32] = buffer_data_0[1167:1160];
        layer0[16][7:0] = buffer_data_4[1143:1136];
        layer0[16][15:8] = buffer_data_4[1151:1144];
        layer0[16][23:16] = buffer_data_4[1159:1152];
        layer0[16][31:24] = buffer_data_4[1167:1160];
        layer0[16][39:32] = buffer_data_4[1175:1168];
        layer1[16][7:0] = buffer_data_3[1143:1136];
        layer1[16][15:8] = buffer_data_3[1151:1144];
        layer1[16][23:16] = buffer_data_3[1159:1152];
        layer1[16][31:24] = buffer_data_3[1167:1160];
        layer1[16][39:32] = buffer_data_3[1175:1168];
        layer2[16][7:0] = buffer_data_2[1143:1136];
        layer2[16][15:8] = buffer_data_2[1151:1144];
        layer2[16][23:16] = buffer_data_2[1159:1152];
        layer2[16][31:24] = buffer_data_2[1167:1160];
        layer2[16][39:32] = buffer_data_2[1175:1168];
        layer3[16][7:0] = buffer_data_1[1143:1136];
        layer3[16][15:8] = buffer_data_1[1151:1144];
        layer3[16][23:16] = buffer_data_1[1159:1152];
        layer3[16][31:24] = buffer_data_1[1167:1160];
        layer3[16][39:32] = buffer_data_1[1175:1168];
        layer4[16][7:0] = buffer_data_0[1143:1136];
        layer4[16][15:8] = buffer_data_0[1151:1144];
        layer4[16][23:16] = buffer_data_0[1159:1152];
        layer4[16][31:24] = buffer_data_0[1167:1160];
        layer4[16][39:32] = buffer_data_0[1175:1168];
        layer0[17][7:0] = buffer_data_4[1151:1144];
        layer0[17][15:8] = buffer_data_4[1159:1152];
        layer0[17][23:16] = buffer_data_4[1167:1160];
        layer0[17][31:24] = buffer_data_4[1175:1168];
        layer0[17][39:32] = buffer_data_4[1183:1176];
        layer1[17][7:0] = buffer_data_3[1151:1144];
        layer1[17][15:8] = buffer_data_3[1159:1152];
        layer1[17][23:16] = buffer_data_3[1167:1160];
        layer1[17][31:24] = buffer_data_3[1175:1168];
        layer1[17][39:32] = buffer_data_3[1183:1176];
        layer2[17][7:0] = buffer_data_2[1151:1144];
        layer2[17][15:8] = buffer_data_2[1159:1152];
        layer2[17][23:16] = buffer_data_2[1167:1160];
        layer2[17][31:24] = buffer_data_2[1175:1168];
        layer2[17][39:32] = buffer_data_2[1183:1176];
        layer3[17][7:0] = buffer_data_1[1151:1144];
        layer3[17][15:8] = buffer_data_1[1159:1152];
        layer3[17][23:16] = buffer_data_1[1167:1160];
        layer3[17][31:24] = buffer_data_1[1175:1168];
        layer3[17][39:32] = buffer_data_1[1183:1176];
        layer4[17][7:0] = buffer_data_0[1151:1144];
        layer4[17][15:8] = buffer_data_0[1159:1152];
        layer4[17][23:16] = buffer_data_0[1167:1160];
        layer4[17][31:24] = buffer_data_0[1175:1168];
        layer4[17][39:32] = buffer_data_0[1183:1176];
        layer0[18][7:0] = buffer_data_4[1159:1152];
        layer0[18][15:8] = buffer_data_4[1167:1160];
        layer0[18][23:16] = buffer_data_4[1175:1168];
        layer0[18][31:24] = buffer_data_4[1183:1176];
        layer0[18][39:32] = buffer_data_4[1191:1184];
        layer1[18][7:0] = buffer_data_3[1159:1152];
        layer1[18][15:8] = buffer_data_3[1167:1160];
        layer1[18][23:16] = buffer_data_3[1175:1168];
        layer1[18][31:24] = buffer_data_3[1183:1176];
        layer1[18][39:32] = buffer_data_3[1191:1184];
        layer2[18][7:0] = buffer_data_2[1159:1152];
        layer2[18][15:8] = buffer_data_2[1167:1160];
        layer2[18][23:16] = buffer_data_2[1175:1168];
        layer2[18][31:24] = buffer_data_2[1183:1176];
        layer2[18][39:32] = buffer_data_2[1191:1184];
        layer3[18][7:0] = buffer_data_1[1159:1152];
        layer3[18][15:8] = buffer_data_1[1167:1160];
        layer3[18][23:16] = buffer_data_1[1175:1168];
        layer3[18][31:24] = buffer_data_1[1183:1176];
        layer3[18][39:32] = buffer_data_1[1191:1184];
        layer4[18][7:0] = buffer_data_0[1159:1152];
        layer4[18][15:8] = buffer_data_0[1167:1160];
        layer4[18][23:16] = buffer_data_0[1175:1168];
        layer4[18][31:24] = buffer_data_0[1183:1176];
        layer4[18][39:32] = buffer_data_0[1191:1184];
        layer0[19][7:0] = buffer_data_4[1167:1160];
        layer0[19][15:8] = buffer_data_4[1175:1168];
        layer0[19][23:16] = buffer_data_4[1183:1176];
        layer0[19][31:24] = buffer_data_4[1191:1184];
        layer0[19][39:32] = buffer_data_4[1199:1192];
        layer1[19][7:0] = buffer_data_3[1167:1160];
        layer1[19][15:8] = buffer_data_3[1175:1168];
        layer1[19][23:16] = buffer_data_3[1183:1176];
        layer1[19][31:24] = buffer_data_3[1191:1184];
        layer1[19][39:32] = buffer_data_3[1199:1192];
        layer2[19][7:0] = buffer_data_2[1167:1160];
        layer2[19][15:8] = buffer_data_2[1175:1168];
        layer2[19][23:16] = buffer_data_2[1183:1176];
        layer2[19][31:24] = buffer_data_2[1191:1184];
        layer2[19][39:32] = buffer_data_2[1199:1192];
        layer3[19][7:0] = buffer_data_1[1167:1160];
        layer3[19][15:8] = buffer_data_1[1175:1168];
        layer3[19][23:16] = buffer_data_1[1183:1176];
        layer3[19][31:24] = buffer_data_1[1191:1184];
        layer3[19][39:32] = buffer_data_1[1199:1192];
        layer4[19][7:0] = buffer_data_0[1167:1160];
        layer4[19][15:8] = buffer_data_0[1175:1168];
        layer4[19][23:16] = buffer_data_0[1183:1176];
        layer4[19][31:24] = buffer_data_0[1191:1184];
        layer4[19][39:32] = buffer_data_0[1199:1192];
        layer0[20][7:0] = buffer_data_4[1175:1168];
        layer0[20][15:8] = buffer_data_4[1183:1176];
        layer0[20][23:16] = buffer_data_4[1191:1184];
        layer0[20][31:24] = buffer_data_4[1199:1192];
        layer0[20][39:32] = buffer_data_4[1207:1200];
        layer1[20][7:0] = buffer_data_3[1175:1168];
        layer1[20][15:8] = buffer_data_3[1183:1176];
        layer1[20][23:16] = buffer_data_3[1191:1184];
        layer1[20][31:24] = buffer_data_3[1199:1192];
        layer1[20][39:32] = buffer_data_3[1207:1200];
        layer2[20][7:0] = buffer_data_2[1175:1168];
        layer2[20][15:8] = buffer_data_2[1183:1176];
        layer2[20][23:16] = buffer_data_2[1191:1184];
        layer2[20][31:24] = buffer_data_2[1199:1192];
        layer2[20][39:32] = buffer_data_2[1207:1200];
        layer3[20][7:0] = buffer_data_1[1175:1168];
        layer3[20][15:8] = buffer_data_1[1183:1176];
        layer3[20][23:16] = buffer_data_1[1191:1184];
        layer3[20][31:24] = buffer_data_1[1199:1192];
        layer3[20][39:32] = buffer_data_1[1207:1200];
        layer4[20][7:0] = buffer_data_0[1175:1168];
        layer4[20][15:8] = buffer_data_0[1183:1176];
        layer4[20][23:16] = buffer_data_0[1191:1184];
        layer4[20][31:24] = buffer_data_0[1199:1192];
        layer4[20][39:32] = buffer_data_0[1207:1200];
        layer0[21][7:0] = buffer_data_4[1183:1176];
        layer0[21][15:8] = buffer_data_4[1191:1184];
        layer0[21][23:16] = buffer_data_4[1199:1192];
        layer0[21][31:24] = buffer_data_4[1207:1200];
        layer0[21][39:32] = buffer_data_4[1215:1208];
        layer1[21][7:0] = buffer_data_3[1183:1176];
        layer1[21][15:8] = buffer_data_3[1191:1184];
        layer1[21][23:16] = buffer_data_3[1199:1192];
        layer1[21][31:24] = buffer_data_3[1207:1200];
        layer1[21][39:32] = buffer_data_3[1215:1208];
        layer2[21][7:0] = buffer_data_2[1183:1176];
        layer2[21][15:8] = buffer_data_2[1191:1184];
        layer2[21][23:16] = buffer_data_2[1199:1192];
        layer2[21][31:24] = buffer_data_2[1207:1200];
        layer2[21][39:32] = buffer_data_2[1215:1208];
        layer3[21][7:0] = buffer_data_1[1183:1176];
        layer3[21][15:8] = buffer_data_1[1191:1184];
        layer3[21][23:16] = buffer_data_1[1199:1192];
        layer3[21][31:24] = buffer_data_1[1207:1200];
        layer3[21][39:32] = buffer_data_1[1215:1208];
        layer4[21][7:0] = buffer_data_0[1183:1176];
        layer4[21][15:8] = buffer_data_0[1191:1184];
        layer4[21][23:16] = buffer_data_0[1199:1192];
        layer4[21][31:24] = buffer_data_0[1207:1200];
        layer4[21][39:32] = buffer_data_0[1215:1208];
        layer0[22][7:0] = buffer_data_4[1191:1184];
        layer0[22][15:8] = buffer_data_4[1199:1192];
        layer0[22][23:16] = buffer_data_4[1207:1200];
        layer0[22][31:24] = buffer_data_4[1215:1208];
        layer0[22][39:32] = buffer_data_4[1223:1216];
        layer1[22][7:0] = buffer_data_3[1191:1184];
        layer1[22][15:8] = buffer_data_3[1199:1192];
        layer1[22][23:16] = buffer_data_3[1207:1200];
        layer1[22][31:24] = buffer_data_3[1215:1208];
        layer1[22][39:32] = buffer_data_3[1223:1216];
        layer2[22][7:0] = buffer_data_2[1191:1184];
        layer2[22][15:8] = buffer_data_2[1199:1192];
        layer2[22][23:16] = buffer_data_2[1207:1200];
        layer2[22][31:24] = buffer_data_2[1215:1208];
        layer2[22][39:32] = buffer_data_2[1223:1216];
        layer3[22][7:0] = buffer_data_1[1191:1184];
        layer3[22][15:8] = buffer_data_1[1199:1192];
        layer3[22][23:16] = buffer_data_1[1207:1200];
        layer3[22][31:24] = buffer_data_1[1215:1208];
        layer3[22][39:32] = buffer_data_1[1223:1216];
        layer4[22][7:0] = buffer_data_0[1191:1184];
        layer4[22][15:8] = buffer_data_0[1199:1192];
        layer4[22][23:16] = buffer_data_0[1207:1200];
        layer4[22][31:24] = buffer_data_0[1215:1208];
        layer4[22][39:32] = buffer_data_0[1223:1216];
        layer0[23][7:0] = buffer_data_4[1199:1192];
        layer0[23][15:8] = buffer_data_4[1207:1200];
        layer0[23][23:16] = buffer_data_4[1215:1208];
        layer0[23][31:24] = buffer_data_4[1223:1216];
        layer0[23][39:32] = buffer_data_4[1231:1224];
        layer1[23][7:0] = buffer_data_3[1199:1192];
        layer1[23][15:8] = buffer_data_3[1207:1200];
        layer1[23][23:16] = buffer_data_3[1215:1208];
        layer1[23][31:24] = buffer_data_3[1223:1216];
        layer1[23][39:32] = buffer_data_3[1231:1224];
        layer2[23][7:0] = buffer_data_2[1199:1192];
        layer2[23][15:8] = buffer_data_2[1207:1200];
        layer2[23][23:16] = buffer_data_2[1215:1208];
        layer2[23][31:24] = buffer_data_2[1223:1216];
        layer2[23][39:32] = buffer_data_2[1231:1224];
        layer3[23][7:0] = buffer_data_1[1199:1192];
        layer3[23][15:8] = buffer_data_1[1207:1200];
        layer3[23][23:16] = buffer_data_1[1215:1208];
        layer3[23][31:24] = buffer_data_1[1223:1216];
        layer3[23][39:32] = buffer_data_1[1231:1224];
        layer4[23][7:0] = buffer_data_0[1199:1192];
        layer4[23][15:8] = buffer_data_0[1207:1200];
        layer4[23][23:16] = buffer_data_0[1215:1208];
        layer4[23][31:24] = buffer_data_0[1223:1216];
        layer4[23][39:32] = buffer_data_0[1231:1224];
        layer0[24][7:0] = buffer_data_4[1207:1200];
        layer0[24][15:8] = buffer_data_4[1215:1208];
        layer0[24][23:16] = buffer_data_4[1223:1216];
        layer0[24][31:24] = buffer_data_4[1231:1224];
        layer0[24][39:32] = buffer_data_4[1239:1232];
        layer1[24][7:0] = buffer_data_3[1207:1200];
        layer1[24][15:8] = buffer_data_3[1215:1208];
        layer1[24][23:16] = buffer_data_3[1223:1216];
        layer1[24][31:24] = buffer_data_3[1231:1224];
        layer1[24][39:32] = buffer_data_3[1239:1232];
        layer2[24][7:0] = buffer_data_2[1207:1200];
        layer2[24][15:8] = buffer_data_2[1215:1208];
        layer2[24][23:16] = buffer_data_2[1223:1216];
        layer2[24][31:24] = buffer_data_2[1231:1224];
        layer2[24][39:32] = buffer_data_2[1239:1232];
        layer3[24][7:0] = buffer_data_1[1207:1200];
        layer3[24][15:8] = buffer_data_1[1215:1208];
        layer3[24][23:16] = buffer_data_1[1223:1216];
        layer3[24][31:24] = buffer_data_1[1231:1224];
        layer3[24][39:32] = buffer_data_1[1239:1232];
        layer4[24][7:0] = buffer_data_0[1207:1200];
        layer4[24][15:8] = buffer_data_0[1215:1208];
        layer4[24][23:16] = buffer_data_0[1223:1216];
        layer4[24][31:24] = buffer_data_0[1231:1224];
        layer4[24][39:32] = buffer_data_0[1239:1232];
        layer0[25][7:0] = buffer_data_4[1215:1208];
        layer0[25][15:8] = buffer_data_4[1223:1216];
        layer0[25][23:16] = buffer_data_4[1231:1224];
        layer0[25][31:24] = buffer_data_4[1239:1232];
        layer0[25][39:32] = buffer_data_4[1247:1240];
        layer1[25][7:0] = buffer_data_3[1215:1208];
        layer1[25][15:8] = buffer_data_3[1223:1216];
        layer1[25][23:16] = buffer_data_3[1231:1224];
        layer1[25][31:24] = buffer_data_3[1239:1232];
        layer1[25][39:32] = buffer_data_3[1247:1240];
        layer2[25][7:0] = buffer_data_2[1215:1208];
        layer2[25][15:8] = buffer_data_2[1223:1216];
        layer2[25][23:16] = buffer_data_2[1231:1224];
        layer2[25][31:24] = buffer_data_2[1239:1232];
        layer2[25][39:32] = buffer_data_2[1247:1240];
        layer3[25][7:0] = buffer_data_1[1215:1208];
        layer3[25][15:8] = buffer_data_1[1223:1216];
        layer3[25][23:16] = buffer_data_1[1231:1224];
        layer3[25][31:24] = buffer_data_1[1239:1232];
        layer3[25][39:32] = buffer_data_1[1247:1240];
        layer4[25][7:0] = buffer_data_0[1215:1208];
        layer4[25][15:8] = buffer_data_0[1223:1216];
        layer4[25][23:16] = buffer_data_0[1231:1224];
        layer4[25][31:24] = buffer_data_0[1239:1232];
        layer4[25][39:32] = buffer_data_0[1247:1240];
        layer0[26][7:0] = buffer_data_4[1223:1216];
        layer0[26][15:8] = buffer_data_4[1231:1224];
        layer0[26][23:16] = buffer_data_4[1239:1232];
        layer0[26][31:24] = buffer_data_4[1247:1240];
        layer0[26][39:32] = buffer_data_4[1255:1248];
        layer1[26][7:0] = buffer_data_3[1223:1216];
        layer1[26][15:8] = buffer_data_3[1231:1224];
        layer1[26][23:16] = buffer_data_3[1239:1232];
        layer1[26][31:24] = buffer_data_3[1247:1240];
        layer1[26][39:32] = buffer_data_3[1255:1248];
        layer2[26][7:0] = buffer_data_2[1223:1216];
        layer2[26][15:8] = buffer_data_2[1231:1224];
        layer2[26][23:16] = buffer_data_2[1239:1232];
        layer2[26][31:24] = buffer_data_2[1247:1240];
        layer2[26][39:32] = buffer_data_2[1255:1248];
        layer3[26][7:0] = buffer_data_1[1223:1216];
        layer3[26][15:8] = buffer_data_1[1231:1224];
        layer3[26][23:16] = buffer_data_1[1239:1232];
        layer3[26][31:24] = buffer_data_1[1247:1240];
        layer3[26][39:32] = buffer_data_1[1255:1248];
        layer4[26][7:0] = buffer_data_0[1223:1216];
        layer4[26][15:8] = buffer_data_0[1231:1224];
        layer4[26][23:16] = buffer_data_0[1239:1232];
        layer4[26][31:24] = buffer_data_0[1247:1240];
        layer4[26][39:32] = buffer_data_0[1255:1248];
        layer0[27][7:0] = buffer_data_4[1231:1224];
        layer0[27][15:8] = buffer_data_4[1239:1232];
        layer0[27][23:16] = buffer_data_4[1247:1240];
        layer0[27][31:24] = buffer_data_4[1255:1248];
        layer0[27][39:32] = buffer_data_4[1263:1256];
        layer1[27][7:0] = buffer_data_3[1231:1224];
        layer1[27][15:8] = buffer_data_3[1239:1232];
        layer1[27][23:16] = buffer_data_3[1247:1240];
        layer1[27][31:24] = buffer_data_3[1255:1248];
        layer1[27][39:32] = buffer_data_3[1263:1256];
        layer2[27][7:0] = buffer_data_2[1231:1224];
        layer2[27][15:8] = buffer_data_2[1239:1232];
        layer2[27][23:16] = buffer_data_2[1247:1240];
        layer2[27][31:24] = buffer_data_2[1255:1248];
        layer2[27][39:32] = buffer_data_2[1263:1256];
        layer3[27][7:0] = buffer_data_1[1231:1224];
        layer3[27][15:8] = buffer_data_1[1239:1232];
        layer3[27][23:16] = buffer_data_1[1247:1240];
        layer3[27][31:24] = buffer_data_1[1255:1248];
        layer3[27][39:32] = buffer_data_1[1263:1256];
        layer4[27][7:0] = buffer_data_0[1231:1224];
        layer4[27][15:8] = buffer_data_0[1239:1232];
        layer4[27][23:16] = buffer_data_0[1247:1240];
        layer4[27][31:24] = buffer_data_0[1255:1248];
        layer4[27][39:32] = buffer_data_0[1263:1256];
        layer0[28][7:0] = buffer_data_4[1239:1232];
        layer0[28][15:8] = buffer_data_4[1247:1240];
        layer0[28][23:16] = buffer_data_4[1255:1248];
        layer0[28][31:24] = buffer_data_4[1263:1256];
        layer0[28][39:32] = buffer_data_4[1271:1264];
        layer1[28][7:0] = buffer_data_3[1239:1232];
        layer1[28][15:8] = buffer_data_3[1247:1240];
        layer1[28][23:16] = buffer_data_3[1255:1248];
        layer1[28][31:24] = buffer_data_3[1263:1256];
        layer1[28][39:32] = buffer_data_3[1271:1264];
        layer2[28][7:0] = buffer_data_2[1239:1232];
        layer2[28][15:8] = buffer_data_2[1247:1240];
        layer2[28][23:16] = buffer_data_2[1255:1248];
        layer2[28][31:24] = buffer_data_2[1263:1256];
        layer2[28][39:32] = buffer_data_2[1271:1264];
        layer3[28][7:0] = buffer_data_1[1239:1232];
        layer3[28][15:8] = buffer_data_1[1247:1240];
        layer3[28][23:16] = buffer_data_1[1255:1248];
        layer3[28][31:24] = buffer_data_1[1263:1256];
        layer3[28][39:32] = buffer_data_1[1271:1264];
        layer4[28][7:0] = buffer_data_0[1239:1232];
        layer4[28][15:8] = buffer_data_0[1247:1240];
        layer4[28][23:16] = buffer_data_0[1255:1248];
        layer4[28][31:24] = buffer_data_0[1263:1256];
        layer4[28][39:32] = buffer_data_0[1271:1264];
        layer0[29][7:0] = buffer_data_4[1247:1240];
        layer0[29][15:8] = buffer_data_4[1255:1248];
        layer0[29][23:16] = buffer_data_4[1263:1256];
        layer0[29][31:24] = buffer_data_4[1271:1264];
        layer0[29][39:32] = buffer_data_4[1279:1272];
        layer1[29][7:0] = buffer_data_3[1247:1240];
        layer1[29][15:8] = buffer_data_3[1255:1248];
        layer1[29][23:16] = buffer_data_3[1263:1256];
        layer1[29][31:24] = buffer_data_3[1271:1264];
        layer1[29][39:32] = buffer_data_3[1279:1272];
        layer2[29][7:0] = buffer_data_2[1247:1240];
        layer2[29][15:8] = buffer_data_2[1255:1248];
        layer2[29][23:16] = buffer_data_2[1263:1256];
        layer2[29][31:24] = buffer_data_2[1271:1264];
        layer2[29][39:32] = buffer_data_2[1279:1272];
        layer3[29][7:0] = buffer_data_1[1247:1240];
        layer3[29][15:8] = buffer_data_1[1255:1248];
        layer3[29][23:16] = buffer_data_1[1263:1256];
        layer3[29][31:24] = buffer_data_1[1271:1264];
        layer3[29][39:32] = buffer_data_1[1279:1272];
        layer4[29][7:0] = buffer_data_0[1247:1240];
        layer4[29][15:8] = buffer_data_0[1255:1248];
        layer4[29][23:16] = buffer_data_0[1263:1256];
        layer4[29][31:24] = buffer_data_0[1271:1264];
        layer4[29][39:32] = buffer_data_0[1279:1272];
        layer0[30][7:0] = buffer_data_4[1255:1248];
        layer0[30][15:8] = buffer_data_4[1263:1256];
        layer0[30][23:16] = buffer_data_4[1271:1264];
        layer0[30][31:24] = buffer_data_4[1279:1272];
        layer0[30][39:32] = buffer_data_4[1287:1280];
        layer1[30][7:0] = buffer_data_3[1255:1248];
        layer1[30][15:8] = buffer_data_3[1263:1256];
        layer1[30][23:16] = buffer_data_3[1271:1264];
        layer1[30][31:24] = buffer_data_3[1279:1272];
        layer1[30][39:32] = buffer_data_3[1287:1280];
        layer2[30][7:0] = buffer_data_2[1255:1248];
        layer2[30][15:8] = buffer_data_2[1263:1256];
        layer2[30][23:16] = buffer_data_2[1271:1264];
        layer2[30][31:24] = buffer_data_2[1279:1272];
        layer2[30][39:32] = buffer_data_2[1287:1280];
        layer3[30][7:0] = buffer_data_1[1255:1248];
        layer3[30][15:8] = buffer_data_1[1263:1256];
        layer3[30][23:16] = buffer_data_1[1271:1264];
        layer3[30][31:24] = buffer_data_1[1279:1272];
        layer3[30][39:32] = buffer_data_1[1287:1280];
        layer4[30][7:0] = buffer_data_0[1255:1248];
        layer4[30][15:8] = buffer_data_0[1263:1256];
        layer4[30][23:16] = buffer_data_0[1271:1264];
        layer4[30][31:24] = buffer_data_0[1279:1272];
        layer4[30][39:32] = buffer_data_0[1287:1280];
        layer0[31][7:0] = buffer_data_4[1263:1256];
        layer0[31][15:8] = buffer_data_4[1271:1264];
        layer0[31][23:16] = buffer_data_4[1279:1272];
        layer0[31][31:24] = buffer_data_4[1287:1280];
        layer0[31][39:32] = buffer_data_4[1295:1288];
        layer1[31][7:0] = buffer_data_3[1263:1256];
        layer1[31][15:8] = buffer_data_3[1271:1264];
        layer1[31][23:16] = buffer_data_3[1279:1272];
        layer1[31][31:24] = buffer_data_3[1287:1280];
        layer1[31][39:32] = buffer_data_3[1295:1288];
        layer2[31][7:0] = buffer_data_2[1263:1256];
        layer2[31][15:8] = buffer_data_2[1271:1264];
        layer2[31][23:16] = buffer_data_2[1279:1272];
        layer2[31][31:24] = buffer_data_2[1287:1280];
        layer2[31][39:32] = buffer_data_2[1295:1288];
        layer3[31][7:0] = buffer_data_1[1263:1256];
        layer3[31][15:8] = buffer_data_1[1271:1264];
        layer3[31][23:16] = buffer_data_1[1279:1272];
        layer3[31][31:24] = buffer_data_1[1287:1280];
        layer3[31][39:32] = buffer_data_1[1295:1288];
        layer4[31][7:0] = buffer_data_0[1263:1256];
        layer4[31][15:8] = buffer_data_0[1271:1264];
        layer4[31][23:16] = buffer_data_0[1279:1272];
        layer4[31][31:24] = buffer_data_0[1287:1280];
        layer4[31][39:32] = buffer_data_0[1295:1288];
        layer0[32][7:0] = buffer_data_4[1271:1264];
        layer0[32][15:8] = buffer_data_4[1279:1272];
        layer0[32][23:16] = buffer_data_4[1287:1280];
        layer0[32][31:24] = buffer_data_4[1295:1288];
        layer0[32][39:32] = buffer_data_4[1303:1296];
        layer1[32][7:0] = buffer_data_3[1271:1264];
        layer1[32][15:8] = buffer_data_3[1279:1272];
        layer1[32][23:16] = buffer_data_3[1287:1280];
        layer1[32][31:24] = buffer_data_3[1295:1288];
        layer1[32][39:32] = buffer_data_3[1303:1296];
        layer2[32][7:0] = buffer_data_2[1271:1264];
        layer2[32][15:8] = buffer_data_2[1279:1272];
        layer2[32][23:16] = buffer_data_2[1287:1280];
        layer2[32][31:24] = buffer_data_2[1295:1288];
        layer2[32][39:32] = buffer_data_2[1303:1296];
        layer3[32][7:0] = buffer_data_1[1271:1264];
        layer3[32][15:8] = buffer_data_1[1279:1272];
        layer3[32][23:16] = buffer_data_1[1287:1280];
        layer3[32][31:24] = buffer_data_1[1295:1288];
        layer3[32][39:32] = buffer_data_1[1303:1296];
        layer4[32][7:0] = buffer_data_0[1271:1264];
        layer4[32][15:8] = buffer_data_0[1279:1272];
        layer4[32][23:16] = buffer_data_0[1287:1280];
        layer4[32][31:24] = buffer_data_0[1295:1288];
        layer4[32][39:32] = buffer_data_0[1303:1296];
        layer0[33][7:0] = buffer_data_4[1279:1272];
        layer0[33][15:8] = buffer_data_4[1287:1280];
        layer0[33][23:16] = buffer_data_4[1295:1288];
        layer0[33][31:24] = buffer_data_4[1303:1296];
        layer0[33][39:32] = buffer_data_4[1311:1304];
        layer1[33][7:0] = buffer_data_3[1279:1272];
        layer1[33][15:8] = buffer_data_3[1287:1280];
        layer1[33][23:16] = buffer_data_3[1295:1288];
        layer1[33][31:24] = buffer_data_3[1303:1296];
        layer1[33][39:32] = buffer_data_3[1311:1304];
        layer2[33][7:0] = buffer_data_2[1279:1272];
        layer2[33][15:8] = buffer_data_2[1287:1280];
        layer2[33][23:16] = buffer_data_2[1295:1288];
        layer2[33][31:24] = buffer_data_2[1303:1296];
        layer2[33][39:32] = buffer_data_2[1311:1304];
        layer3[33][7:0] = buffer_data_1[1279:1272];
        layer3[33][15:8] = buffer_data_1[1287:1280];
        layer3[33][23:16] = buffer_data_1[1295:1288];
        layer3[33][31:24] = buffer_data_1[1303:1296];
        layer3[33][39:32] = buffer_data_1[1311:1304];
        layer4[33][7:0] = buffer_data_0[1279:1272];
        layer4[33][15:8] = buffer_data_0[1287:1280];
        layer4[33][23:16] = buffer_data_0[1295:1288];
        layer4[33][31:24] = buffer_data_0[1303:1296];
        layer4[33][39:32] = buffer_data_0[1311:1304];
        layer0[34][7:0] = buffer_data_4[1287:1280];
        layer0[34][15:8] = buffer_data_4[1295:1288];
        layer0[34][23:16] = buffer_data_4[1303:1296];
        layer0[34][31:24] = buffer_data_4[1311:1304];
        layer0[34][39:32] = buffer_data_4[1319:1312];
        layer1[34][7:0] = buffer_data_3[1287:1280];
        layer1[34][15:8] = buffer_data_3[1295:1288];
        layer1[34][23:16] = buffer_data_3[1303:1296];
        layer1[34][31:24] = buffer_data_3[1311:1304];
        layer1[34][39:32] = buffer_data_3[1319:1312];
        layer2[34][7:0] = buffer_data_2[1287:1280];
        layer2[34][15:8] = buffer_data_2[1295:1288];
        layer2[34][23:16] = buffer_data_2[1303:1296];
        layer2[34][31:24] = buffer_data_2[1311:1304];
        layer2[34][39:32] = buffer_data_2[1319:1312];
        layer3[34][7:0] = buffer_data_1[1287:1280];
        layer3[34][15:8] = buffer_data_1[1295:1288];
        layer3[34][23:16] = buffer_data_1[1303:1296];
        layer3[34][31:24] = buffer_data_1[1311:1304];
        layer3[34][39:32] = buffer_data_1[1319:1312];
        layer4[34][7:0] = buffer_data_0[1287:1280];
        layer4[34][15:8] = buffer_data_0[1295:1288];
        layer4[34][23:16] = buffer_data_0[1303:1296];
        layer4[34][31:24] = buffer_data_0[1311:1304];
        layer4[34][39:32] = buffer_data_0[1319:1312];
        layer0[35][7:0] = buffer_data_4[1295:1288];
        layer0[35][15:8] = buffer_data_4[1303:1296];
        layer0[35][23:16] = buffer_data_4[1311:1304];
        layer0[35][31:24] = buffer_data_4[1319:1312];
        layer0[35][39:32] = buffer_data_4[1327:1320];
        layer1[35][7:0] = buffer_data_3[1295:1288];
        layer1[35][15:8] = buffer_data_3[1303:1296];
        layer1[35][23:16] = buffer_data_3[1311:1304];
        layer1[35][31:24] = buffer_data_3[1319:1312];
        layer1[35][39:32] = buffer_data_3[1327:1320];
        layer2[35][7:0] = buffer_data_2[1295:1288];
        layer2[35][15:8] = buffer_data_2[1303:1296];
        layer2[35][23:16] = buffer_data_2[1311:1304];
        layer2[35][31:24] = buffer_data_2[1319:1312];
        layer2[35][39:32] = buffer_data_2[1327:1320];
        layer3[35][7:0] = buffer_data_1[1295:1288];
        layer3[35][15:8] = buffer_data_1[1303:1296];
        layer3[35][23:16] = buffer_data_1[1311:1304];
        layer3[35][31:24] = buffer_data_1[1319:1312];
        layer3[35][39:32] = buffer_data_1[1327:1320];
        layer4[35][7:0] = buffer_data_0[1295:1288];
        layer4[35][15:8] = buffer_data_0[1303:1296];
        layer4[35][23:16] = buffer_data_0[1311:1304];
        layer4[35][31:24] = buffer_data_0[1319:1312];
        layer4[35][39:32] = buffer_data_0[1327:1320];
        layer0[36][7:0] = buffer_data_4[1303:1296];
        layer0[36][15:8] = buffer_data_4[1311:1304];
        layer0[36][23:16] = buffer_data_4[1319:1312];
        layer0[36][31:24] = buffer_data_4[1327:1320];
        layer0[36][39:32] = buffer_data_4[1335:1328];
        layer1[36][7:0] = buffer_data_3[1303:1296];
        layer1[36][15:8] = buffer_data_3[1311:1304];
        layer1[36][23:16] = buffer_data_3[1319:1312];
        layer1[36][31:24] = buffer_data_3[1327:1320];
        layer1[36][39:32] = buffer_data_3[1335:1328];
        layer2[36][7:0] = buffer_data_2[1303:1296];
        layer2[36][15:8] = buffer_data_2[1311:1304];
        layer2[36][23:16] = buffer_data_2[1319:1312];
        layer2[36][31:24] = buffer_data_2[1327:1320];
        layer2[36][39:32] = buffer_data_2[1335:1328];
        layer3[36][7:0] = buffer_data_1[1303:1296];
        layer3[36][15:8] = buffer_data_1[1311:1304];
        layer3[36][23:16] = buffer_data_1[1319:1312];
        layer3[36][31:24] = buffer_data_1[1327:1320];
        layer3[36][39:32] = buffer_data_1[1335:1328];
        layer4[36][7:0] = buffer_data_0[1303:1296];
        layer4[36][15:8] = buffer_data_0[1311:1304];
        layer4[36][23:16] = buffer_data_0[1319:1312];
        layer4[36][31:24] = buffer_data_0[1327:1320];
        layer4[36][39:32] = buffer_data_0[1335:1328];
        layer0[37][7:0] = buffer_data_4[1311:1304];
        layer0[37][15:8] = buffer_data_4[1319:1312];
        layer0[37][23:16] = buffer_data_4[1327:1320];
        layer0[37][31:24] = buffer_data_4[1335:1328];
        layer0[37][39:32] = buffer_data_4[1343:1336];
        layer1[37][7:0] = buffer_data_3[1311:1304];
        layer1[37][15:8] = buffer_data_3[1319:1312];
        layer1[37][23:16] = buffer_data_3[1327:1320];
        layer1[37][31:24] = buffer_data_3[1335:1328];
        layer1[37][39:32] = buffer_data_3[1343:1336];
        layer2[37][7:0] = buffer_data_2[1311:1304];
        layer2[37][15:8] = buffer_data_2[1319:1312];
        layer2[37][23:16] = buffer_data_2[1327:1320];
        layer2[37][31:24] = buffer_data_2[1335:1328];
        layer2[37][39:32] = buffer_data_2[1343:1336];
        layer3[37][7:0] = buffer_data_1[1311:1304];
        layer3[37][15:8] = buffer_data_1[1319:1312];
        layer3[37][23:16] = buffer_data_1[1327:1320];
        layer3[37][31:24] = buffer_data_1[1335:1328];
        layer3[37][39:32] = buffer_data_1[1343:1336];
        layer4[37][7:0] = buffer_data_0[1311:1304];
        layer4[37][15:8] = buffer_data_0[1319:1312];
        layer4[37][23:16] = buffer_data_0[1327:1320];
        layer4[37][31:24] = buffer_data_0[1335:1328];
        layer4[37][39:32] = buffer_data_0[1343:1336];
        layer0[38][7:0] = buffer_data_4[1319:1312];
        layer0[38][15:8] = buffer_data_4[1327:1320];
        layer0[38][23:16] = buffer_data_4[1335:1328];
        layer0[38][31:24] = buffer_data_4[1343:1336];
        layer0[38][39:32] = buffer_data_4[1351:1344];
        layer1[38][7:0] = buffer_data_3[1319:1312];
        layer1[38][15:8] = buffer_data_3[1327:1320];
        layer1[38][23:16] = buffer_data_3[1335:1328];
        layer1[38][31:24] = buffer_data_3[1343:1336];
        layer1[38][39:32] = buffer_data_3[1351:1344];
        layer2[38][7:0] = buffer_data_2[1319:1312];
        layer2[38][15:8] = buffer_data_2[1327:1320];
        layer2[38][23:16] = buffer_data_2[1335:1328];
        layer2[38][31:24] = buffer_data_2[1343:1336];
        layer2[38][39:32] = buffer_data_2[1351:1344];
        layer3[38][7:0] = buffer_data_1[1319:1312];
        layer3[38][15:8] = buffer_data_1[1327:1320];
        layer3[38][23:16] = buffer_data_1[1335:1328];
        layer3[38][31:24] = buffer_data_1[1343:1336];
        layer3[38][39:32] = buffer_data_1[1351:1344];
        layer4[38][7:0] = buffer_data_0[1319:1312];
        layer4[38][15:8] = buffer_data_0[1327:1320];
        layer4[38][23:16] = buffer_data_0[1335:1328];
        layer4[38][31:24] = buffer_data_0[1343:1336];
        layer4[38][39:32] = buffer_data_0[1351:1344];
        layer0[39][7:0] = buffer_data_4[1327:1320];
        layer0[39][15:8] = buffer_data_4[1335:1328];
        layer0[39][23:16] = buffer_data_4[1343:1336];
        layer0[39][31:24] = buffer_data_4[1351:1344];
        layer0[39][39:32] = buffer_data_4[1359:1352];
        layer1[39][7:0] = buffer_data_3[1327:1320];
        layer1[39][15:8] = buffer_data_3[1335:1328];
        layer1[39][23:16] = buffer_data_3[1343:1336];
        layer1[39][31:24] = buffer_data_3[1351:1344];
        layer1[39][39:32] = buffer_data_3[1359:1352];
        layer2[39][7:0] = buffer_data_2[1327:1320];
        layer2[39][15:8] = buffer_data_2[1335:1328];
        layer2[39][23:16] = buffer_data_2[1343:1336];
        layer2[39][31:24] = buffer_data_2[1351:1344];
        layer2[39][39:32] = buffer_data_2[1359:1352];
        layer3[39][7:0] = buffer_data_1[1327:1320];
        layer3[39][15:8] = buffer_data_1[1335:1328];
        layer3[39][23:16] = buffer_data_1[1343:1336];
        layer3[39][31:24] = buffer_data_1[1351:1344];
        layer3[39][39:32] = buffer_data_1[1359:1352];
        layer4[39][7:0] = buffer_data_0[1327:1320];
        layer4[39][15:8] = buffer_data_0[1335:1328];
        layer4[39][23:16] = buffer_data_0[1343:1336];
        layer4[39][31:24] = buffer_data_0[1351:1344];
        layer4[39][39:32] = buffer_data_0[1359:1352];
        layer0[40][7:0] = buffer_data_4[1335:1328];
        layer0[40][15:8] = buffer_data_4[1343:1336];
        layer0[40][23:16] = buffer_data_4[1351:1344];
        layer0[40][31:24] = buffer_data_4[1359:1352];
        layer0[40][39:32] = buffer_data_4[1367:1360];
        layer1[40][7:0] = buffer_data_3[1335:1328];
        layer1[40][15:8] = buffer_data_3[1343:1336];
        layer1[40][23:16] = buffer_data_3[1351:1344];
        layer1[40][31:24] = buffer_data_3[1359:1352];
        layer1[40][39:32] = buffer_data_3[1367:1360];
        layer2[40][7:0] = buffer_data_2[1335:1328];
        layer2[40][15:8] = buffer_data_2[1343:1336];
        layer2[40][23:16] = buffer_data_2[1351:1344];
        layer2[40][31:24] = buffer_data_2[1359:1352];
        layer2[40][39:32] = buffer_data_2[1367:1360];
        layer3[40][7:0] = buffer_data_1[1335:1328];
        layer3[40][15:8] = buffer_data_1[1343:1336];
        layer3[40][23:16] = buffer_data_1[1351:1344];
        layer3[40][31:24] = buffer_data_1[1359:1352];
        layer3[40][39:32] = buffer_data_1[1367:1360];
        layer4[40][7:0] = buffer_data_0[1335:1328];
        layer4[40][15:8] = buffer_data_0[1343:1336];
        layer4[40][23:16] = buffer_data_0[1351:1344];
        layer4[40][31:24] = buffer_data_0[1359:1352];
        layer4[40][39:32] = buffer_data_0[1367:1360];
        layer0[41][7:0] = buffer_data_4[1343:1336];
        layer0[41][15:8] = buffer_data_4[1351:1344];
        layer0[41][23:16] = buffer_data_4[1359:1352];
        layer0[41][31:24] = buffer_data_4[1367:1360];
        layer0[41][39:32] = buffer_data_4[1375:1368];
        layer1[41][7:0] = buffer_data_3[1343:1336];
        layer1[41][15:8] = buffer_data_3[1351:1344];
        layer1[41][23:16] = buffer_data_3[1359:1352];
        layer1[41][31:24] = buffer_data_3[1367:1360];
        layer1[41][39:32] = buffer_data_3[1375:1368];
        layer2[41][7:0] = buffer_data_2[1343:1336];
        layer2[41][15:8] = buffer_data_2[1351:1344];
        layer2[41][23:16] = buffer_data_2[1359:1352];
        layer2[41][31:24] = buffer_data_2[1367:1360];
        layer2[41][39:32] = buffer_data_2[1375:1368];
        layer3[41][7:0] = buffer_data_1[1343:1336];
        layer3[41][15:8] = buffer_data_1[1351:1344];
        layer3[41][23:16] = buffer_data_1[1359:1352];
        layer3[41][31:24] = buffer_data_1[1367:1360];
        layer3[41][39:32] = buffer_data_1[1375:1368];
        layer4[41][7:0] = buffer_data_0[1343:1336];
        layer4[41][15:8] = buffer_data_0[1351:1344];
        layer4[41][23:16] = buffer_data_0[1359:1352];
        layer4[41][31:24] = buffer_data_0[1367:1360];
        layer4[41][39:32] = buffer_data_0[1375:1368];
        layer0[42][7:0] = buffer_data_4[1351:1344];
        layer0[42][15:8] = buffer_data_4[1359:1352];
        layer0[42][23:16] = buffer_data_4[1367:1360];
        layer0[42][31:24] = buffer_data_4[1375:1368];
        layer0[42][39:32] = buffer_data_4[1383:1376];
        layer1[42][7:0] = buffer_data_3[1351:1344];
        layer1[42][15:8] = buffer_data_3[1359:1352];
        layer1[42][23:16] = buffer_data_3[1367:1360];
        layer1[42][31:24] = buffer_data_3[1375:1368];
        layer1[42][39:32] = buffer_data_3[1383:1376];
        layer2[42][7:0] = buffer_data_2[1351:1344];
        layer2[42][15:8] = buffer_data_2[1359:1352];
        layer2[42][23:16] = buffer_data_2[1367:1360];
        layer2[42][31:24] = buffer_data_2[1375:1368];
        layer2[42][39:32] = buffer_data_2[1383:1376];
        layer3[42][7:0] = buffer_data_1[1351:1344];
        layer3[42][15:8] = buffer_data_1[1359:1352];
        layer3[42][23:16] = buffer_data_1[1367:1360];
        layer3[42][31:24] = buffer_data_1[1375:1368];
        layer3[42][39:32] = buffer_data_1[1383:1376];
        layer4[42][7:0] = buffer_data_0[1351:1344];
        layer4[42][15:8] = buffer_data_0[1359:1352];
        layer4[42][23:16] = buffer_data_0[1367:1360];
        layer4[42][31:24] = buffer_data_0[1375:1368];
        layer4[42][39:32] = buffer_data_0[1383:1376];
        layer0[43][7:0] = buffer_data_4[1359:1352];
        layer0[43][15:8] = buffer_data_4[1367:1360];
        layer0[43][23:16] = buffer_data_4[1375:1368];
        layer0[43][31:24] = buffer_data_4[1383:1376];
        layer0[43][39:32] = buffer_data_4[1391:1384];
        layer1[43][7:0] = buffer_data_3[1359:1352];
        layer1[43][15:8] = buffer_data_3[1367:1360];
        layer1[43][23:16] = buffer_data_3[1375:1368];
        layer1[43][31:24] = buffer_data_3[1383:1376];
        layer1[43][39:32] = buffer_data_3[1391:1384];
        layer2[43][7:0] = buffer_data_2[1359:1352];
        layer2[43][15:8] = buffer_data_2[1367:1360];
        layer2[43][23:16] = buffer_data_2[1375:1368];
        layer2[43][31:24] = buffer_data_2[1383:1376];
        layer2[43][39:32] = buffer_data_2[1391:1384];
        layer3[43][7:0] = buffer_data_1[1359:1352];
        layer3[43][15:8] = buffer_data_1[1367:1360];
        layer3[43][23:16] = buffer_data_1[1375:1368];
        layer3[43][31:24] = buffer_data_1[1383:1376];
        layer3[43][39:32] = buffer_data_1[1391:1384];
        layer4[43][7:0] = buffer_data_0[1359:1352];
        layer4[43][15:8] = buffer_data_0[1367:1360];
        layer4[43][23:16] = buffer_data_0[1375:1368];
        layer4[43][31:24] = buffer_data_0[1383:1376];
        layer4[43][39:32] = buffer_data_0[1391:1384];
        layer0[44][7:0] = buffer_data_4[1367:1360];
        layer0[44][15:8] = buffer_data_4[1375:1368];
        layer0[44][23:16] = buffer_data_4[1383:1376];
        layer0[44][31:24] = buffer_data_4[1391:1384];
        layer0[44][39:32] = buffer_data_4[1399:1392];
        layer1[44][7:0] = buffer_data_3[1367:1360];
        layer1[44][15:8] = buffer_data_3[1375:1368];
        layer1[44][23:16] = buffer_data_3[1383:1376];
        layer1[44][31:24] = buffer_data_3[1391:1384];
        layer1[44][39:32] = buffer_data_3[1399:1392];
        layer2[44][7:0] = buffer_data_2[1367:1360];
        layer2[44][15:8] = buffer_data_2[1375:1368];
        layer2[44][23:16] = buffer_data_2[1383:1376];
        layer2[44][31:24] = buffer_data_2[1391:1384];
        layer2[44][39:32] = buffer_data_2[1399:1392];
        layer3[44][7:0] = buffer_data_1[1367:1360];
        layer3[44][15:8] = buffer_data_1[1375:1368];
        layer3[44][23:16] = buffer_data_1[1383:1376];
        layer3[44][31:24] = buffer_data_1[1391:1384];
        layer3[44][39:32] = buffer_data_1[1399:1392];
        layer4[44][7:0] = buffer_data_0[1367:1360];
        layer4[44][15:8] = buffer_data_0[1375:1368];
        layer4[44][23:16] = buffer_data_0[1383:1376];
        layer4[44][31:24] = buffer_data_0[1391:1384];
        layer4[44][39:32] = buffer_data_0[1399:1392];
        layer0[45][7:0] = buffer_data_4[1375:1368];
        layer0[45][15:8] = buffer_data_4[1383:1376];
        layer0[45][23:16] = buffer_data_4[1391:1384];
        layer0[45][31:24] = buffer_data_4[1399:1392];
        layer0[45][39:32] = buffer_data_4[1407:1400];
        layer1[45][7:0] = buffer_data_3[1375:1368];
        layer1[45][15:8] = buffer_data_3[1383:1376];
        layer1[45][23:16] = buffer_data_3[1391:1384];
        layer1[45][31:24] = buffer_data_3[1399:1392];
        layer1[45][39:32] = buffer_data_3[1407:1400];
        layer2[45][7:0] = buffer_data_2[1375:1368];
        layer2[45][15:8] = buffer_data_2[1383:1376];
        layer2[45][23:16] = buffer_data_2[1391:1384];
        layer2[45][31:24] = buffer_data_2[1399:1392];
        layer2[45][39:32] = buffer_data_2[1407:1400];
        layer3[45][7:0] = buffer_data_1[1375:1368];
        layer3[45][15:8] = buffer_data_1[1383:1376];
        layer3[45][23:16] = buffer_data_1[1391:1384];
        layer3[45][31:24] = buffer_data_1[1399:1392];
        layer3[45][39:32] = buffer_data_1[1407:1400];
        layer4[45][7:0] = buffer_data_0[1375:1368];
        layer4[45][15:8] = buffer_data_0[1383:1376];
        layer4[45][23:16] = buffer_data_0[1391:1384];
        layer4[45][31:24] = buffer_data_0[1399:1392];
        layer4[45][39:32] = buffer_data_0[1407:1400];
        layer0[46][7:0] = buffer_data_4[1383:1376];
        layer0[46][15:8] = buffer_data_4[1391:1384];
        layer0[46][23:16] = buffer_data_4[1399:1392];
        layer0[46][31:24] = buffer_data_4[1407:1400];
        layer0[46][39:32] = buffer_data_4[1415:1408];
        layer1[46][7:0] = buffer_data_3[1383:1376];
        layer1[46][15:8] = buffer_data_3[1391:1384];
        layer1[46][23:16] = buffer_data_3[1399:1392];
        layer1[46][31:24] = buffer_data_3[1407:1400];
        layer1[46][39:32] = buffer_data_3[1415:1408];
        layer2[46][7:0] = buffer_data_2[1383:1376];
        layer2[46][15:8] = buffer_data_2[1391:1384];
        layer2[46][23:16] = buffer_data_2[1399:1392];
        layer2[46][31:24] = buffer_data_2[1407:1400];
        layer2[46][39:32] = buffer_data_2[1415:1408];
        layer3[46][7:0] = buffer_data_1[1383:1376];
        layer3[46][15:8] = buffer_data_1[1391:1384];
        layer3[46][23:16] = buffer_data_1[1399:1392];
        layer3[46][31:24] = buffer_data_1[1407:1400];
        layer3[46][39:32] = buffer_data_1[1415:1408];
        layer4[46][7:0] = buffer_data_0[1383:1376];
        layer4[46][15:8] = buffer_data_0[1391:1384];
        layer4[46][23:16] = buffer_data_0[1399:1392];
        layer4[46][31:24] = buffer_data_0[1407:1400];
        layer4[46][39:32] = buffer_data_0[1415:1408];
        layer0[47][7:0] = buffer_data_4[1391:1384];
        layer0[47][15:8] = buffer_data_4[1399:1392];
        layer0[47][23:16] = buffer_data_4[1407:1400];
        layer0[47][31:24] = buffer_data_4[1415:1408];
        layer0[47][39:32] = buffer_data_4[1423:1416];
        layer1[47][7:0] = buffer_data_3[1391:1384];
        layer1[47][15:8] = buffer_data_3[1399:1392];
        layer1[47][23:16] = buffer_data_3[1407:1400];
        layer1[47][31:24] = buffer_data_3[1415:1408];
        layer1[47][39:32] = buffer_data_3[1423:1416];
        layer2[47][7:0] = buffer_data_2[1391:1384];
        layer2[47][15:8] = buffer_data_2[1399:1392];
        layer2[47][23:16] = buffer_data_2[1407:1400];
        layer2[47][31:24] = buffer_data_2[1415:1408];
        layer2[47][39:32] = buffer_data_2[1423:1416];
        layer3[47][7:0] = buffer_data_1[1391:1384];
        layer3[47][15:8] = buffer_data_1[1399:1392];
        layer3[47][23:16] = buffer_data_1[1407:1400];
        layer3[47][31:24] = buffer_data_1[1415:1408];
        layer3[47][39:32] = buffer_data_1[1423:1416];
        layer4[47][7:0] = buffer_data_0[1391:1384];
        layer4[47][15:8] = buffer_data_0[1399:1392];
        layer4[47][23:16] = buffer_data_0[1407:1400];
        layer4[47][31:24] = buffer_data_0[1415:1408];
        layer4[47][39:32] = buffer_data_0[1423:1416];
        layer0[48][7:0] = buffer_data_4[1399:1392];
        layer0[48][15:8] = buffer_data_4[1407:1400];
        layer0[48][23:16] = buffer_data_4[1415:1408];
        layer0[48][31:24] = buffer_data_4[1423:1416];
        layer0[48][39:32] = buffer_data_4[1431:1424];
        layer1[48][7:0] = buffer_data_3[1399:1392];
        layer1[48][15:8] = buffer_data_3[1407:1400];
        layer1[48][23:16] = buffer_data_3[1415:1408];
        layer1[48][31:24] = buffer_data_3[1423:1416];
        layer1[48][39:32] = buffer_data_3[1431:1424];
        layer2[48][7:0] = buffer_data_2[1399:1392];
        layer2[48][15:8] = buffer_data_2[1407:1400];
        layer2[48][23:16] = buffer_data_2[1415:1408];
        layer2[48][31:24] = buffer_data_2[1423:1416];
        layer2[48][39:32] = buffer_data_2[1431:1424];
        layer3[48][7:0] = buffer_data_1[1399:1392];
        layer3[48][15:8] = buffer_data_1[1407:1400];
        layer3[48][23:16] = buffer_data_1[1415:1408];
        layer3[48][31:24] = buffer_data_1[1423:1416];
        layer3[48][39:32] = buffer_data_1[1431:1424];
        layer4[48][7:0] = buffer_data_0[1399:1392];
        layer4[48][15:8] = buffer_data_0[1407:1400];
        layer4[48][23:16] = buffer_data_0[1415:1408];
        layer4[48][31:24] = buffer_data_0[1423:1416];
        layer4[48][39:32] = buffer_data_0[1431:1424];
        layer0[49][7:0] = buffer_data_4[1407:1400];
        layer0[49][15:8] = buffer_data_4[1415:1408];
        layer0[49][23:16] = buffer_data_4[1423:1416];
        layer0[49][31:24] = buffer_data_4[1431:1424];
        layer0[49][39:32] = buffer_data_4[1439:1432];
        layer1[49][7:0] = buffer_data_3[1407:1400];
        layer1[49][15:8] = buffer_data_3[1415:1408];
        layer1[49][23:16] = buffer_data_3[1423:1416];
        layer1[49][31:24] = buffer_data_3[1431:1424];
        layer1[49][39:32] = buffer_data_3[1439:1432];
        layer2[49][7:0] = buffer_data_2[1407:1400];
        layer2[49][15:8] = buffer_data_2[1415:1408];
        layer2[49][23:16] = buffer_data_2[1423:1416];
        layer2[49][31:24] = buffer_data_2[1431:1424];
        layer2[49][39:32] = buffer_data_2[1439:1432];
        layer3[49][7:0] = buffer_data_1[1407:1400];
        layer3[49][15:8] = buffer_data_1[1415:1408];
        layer3[49][23:16] = buffer_data_1[1423:1416];
        layer3[49][31:24] = buffer_data_1[1431:1424];
        layer3[49][39:32] = buffer_data_1[1439:1432];
        layer4[49][7:0] = buffer_data_0[1407:1400];
        layer4[49][15:8] = buffer_data_0[1415:1408];
        layer4[49][23:16] = buffer_data_0[1423:1416];
        layer4[49][31:24] = buffer_data_0[1431:1424];
        layer4[49][39:32] = buffer_data_0[1439:1432];
        layer0[50][7:0] = buffer_data_4[1415:1408];
        layer0[50][15:8] = buffer_data_4[1423:1416];
        layer0[50][23:16] = buffer_data_4[1431:1424];
        layer0[50][31:24] = buffer_data_4[1439:1432];
        layer0[50][39:32] = buffer_data_4[1447:1440];
        layer1[50][7:0] = buffer_data_3[1415:1408];
        layer1[50][15:8] = buffer_data_3[1423:1416];
        layer1[50][23:16] = buffer_data_3[1431:1424];
        layer1[50][31:24] = buffer_data_3[1439:1432];
        layer1[50][39:32] = buffer_data_3[1447:1440];
        layer2[50][7:0] = buffer_data_2[1415:1408];
        layer2[50][15:8] = buffer_data_2[1423:1416];
        layer2[50][23:16] = buffer_data_2[1431:1424];
        layer2[50][31:24] = buffer_data_2[1439:1432];
        layer2[50][39:32] = buffer_data_2[1447:1440];
        layer3[50][7:0] = buffer_data_1[1415:1408];
        layer3[50][15:8] = buffer_data_1[1423:1416];
        layer3[50][23:16] = buffer_data_1[1431:1424];
        layer3[50][31:24] = buffer_data_1[1439:1432];
        layer3[50][39:32] = buffer_data_1[1447:1440];
        layer4[50][7:0] = buffer_data_0[1415:1408];
        layer4[50][15:8] = buffer_data_0[1423:1416];
        layer4[50][23:16] = buffer_data_0[1431:1424];
        layer4[50][31:24] = buffer_data_0[1439:1432];
        layer4[50][39:32] = buffer_data_0[1447:1440];
        layer0[51][7:0] = buffer_data_4[1423:1416];
        layer0[51][15:8] = buffer_data_4[1431:1424];
        layer0[51][23:16] = buffer_data_4[1439:1432];
        layer0[51][31:24] = buffer_data_4[1447:1440];
        layer0[51][39:32] = buffer_data_4[1455:1448];
        layer1[51][7:0] = buffer_data_3[1423:1416];
        layer1[51][15:8] = buffer_data_3[1431:1424];
        layer1[51][23:16] = buffer_data_3[1439:1432];
        layer1[51][31:24] = buffer_data_3[1447:1440];
        layer1[51][39:32] = buffer_data_3[1455:1448];
        layer2[51][7:0] = buffer_data_2[1423:1416];
        layer2[51][15:8] = buffer_data_2[1431:1424];
        layer2[51][23:16] = buffer_data_2[1439:1432];
        layer2[51][31:24] = buffer_data_2[1447:1440];
        layer2[51][39:32] = buffer_data_2[1455:1448];
        layer3[51][7:0] = buffer_data_1[1423:1416];
        layer3[51][15:8] = buffer_data_1[1431:1424];
        layer3[51][23:16] = buffer_data_1[1439:1432];
        layer3[51][31:24] = buffer_data_1[1447:1440];
        layer3[51][39:32] = buffer_data_1[1455:1448];
        layer4[51][7:0] = buffer_data_0[1423:1416];
        layer4[51][15:8] = buffer_data_0[1431:1424];
        layer4[51][23:16] = buffer_data_0[1439:1432];
        layer4[51][31:24] = buffer_data_0[1447:1440];
        layer4[51][39:32] = buffer_data_0[1455:1448];
        layer0[52][7:0] = buffer_data_4[1431:1424];
        layer0[52][15:8] = buffer_data_4[1439:1432];
        layer0[52][23:16] = buffer_data_4[1447:1440];
        layer0[52][31:24] = buffer_data_4[1455:1448];
        layer0[52][39:32] = buffer_data_4[1463:1456];
        layer1[52][7:0] = buffer_data_3[1431:1424];
        layer1[52][15:8] = buffer_data_3[1439:1432];
        layer1[52][23:16] = buffer_data_3[1447:1440];
        layer1[52][31:24] = buffer_data_3[1455:1448];
        layer1[52][39:32] = buffer_data_3[1463:1456];
        layer2[52][7:0] = buffer_data_2[1431:1424];
        layer2[52][15:8] = buffer_data_2[1439:1432];
        layer2[52][23:16] = buffer_data_2[1447:1440];
        layer2[52][31:24] = buffer_data_2[1455:1448];
        layer2[52][39:32] = buffer_data_2[1463:1456];
        layer3[52][7:0] = buffer_data_1[1431:1424];
        layer3[52][15:8] = buffer_data_1[1439:1432];
        layer3[52][23:16] = buffer_data_1[1447:1440];
        layer3[52][31:24] = buffer_data_1[1455:1448];
        layer3[52][39:32] = buffer_data_1[1463:1456];
        layer4[52][7:0] = buffer_data_0[1431:1424];
        layer4[52][15:8] = buffer_data_0[1439:1432];
        layer4[52][23:16] = buffer_data_0[1447:1440];
        layer4[52][31:24] = buffer_data_0[1455:1448];
        layer4[52][39:32] = buffer_data_0[1463:1456];
        layer0[53][7:0] = buffer_data_4[1439:1432];
        layer0[53][15:8] = buffer_data_4[1447:1440];
        layer0[53][23:16] = buffer_data_4[1455:1448];
        layer0[53][31:24] = buffer_data_4[1463:1456];
        layer0[53][39:32] = buffer_data_4[1471:1464];
        layer1[53][7:0] = buffer_data_3[1439:1432];
        layer1[53][15:8] = buffer_data_3[1447:1440];
        layer1[53][23:16] = buffer_data_3[1455:1448];
        layer1[53][31:24] = buffer_data_3[1463:1456];
        layer1[53][39:32] = buffer_data_3[1471:1464];
        layer2[53][7:0] = buffer_data_2[1439:1432];
        layer2[53][15:8] = buffer_data_2[1447:1440];
        layer2[53][23:16] = buffer_data_2[1455:1448];
        layer2[53][31:24] = buffer_data_2[1463:1456];
        layer2[53][39:32] = buffer_data_2[1471:1464];
        layer3[53][7:0] = buffer_data_1[1439:1432];
        layer3[53][15:8] = buffer_data_1[1447:1440];
        layer3[53][23:16] = buffer_data_1[1455:1448];
        layer3[53][31:24] = buffer_data_1[1463:1456];
        layer3[53][39:32] = buffer_data_1[1471:1464];
        layer4[53][7:0] = buffer_data_0[1439:1432];
        layer4[53][15:8] = buffer_data_0[1447:1440];
        layer4[53][23:16] = buffer_data_0[1455:1448];
        layer4[53][31:24] = buffer_data_0[1463:1456];
        layer4[53][39:32] = buffer_data_0[1471:1464];
        layer0[54][7:0] = buffer_data_4[1447:1440];
        layer0[54][15:8] = buffer_data_4[1455:1448];
        layer0[54][23:16] = buffer_data_4[1463:1456];
        layer0[54][31:24] = buffer_data_4[1471:1464];
        layer0[54][39:32] = buffer_data_4[1479:1472];
        layer1[54][7:0] = buffer_data_3[1447:1440];
        layer1[54][15:8] = buffer_data_3[1455:1448];
        layer1[54][23:16] = buffer_data_3[1463:1456];
        layer1[54][31:24] = buffer_data_3[1471:1464];
        layer1[54][39:32] = buffer_data_3[1479:1472];
        layer2[54][7:0] = buffer_data_2[1447:1440];
        layer2[54][15:8] = buffer_data_2[1455:1448];
        layer2[54][23:16] = buffer_data_2[1463:1456];
        layer2[54][31:24] = buffer_data_2[1471:1464];
        layer2[54][39:32] = buffer_data_2[1479:1472];
        layer3[54][7:0] = buffer_data_1[1447:1440];
        layer3[54][15:8] = buffer_data_1[1455:1448];
        layer3[54][23:16] = buffer_data_1[1463:1456];
        layer3[54][31:24] = buffer_data_1[1471:1464];
        layer3[54][39:32] = buffer_data_1[1479:1472];
        layer4[54][7:0] = buffer_data_0[1447:1440];
        layer4[54][15:8] = buffer_data_0[1455:1448];
        layer4[54][23:16] = buffer_data_0[1463:1456];
        layer4[54][31:24] = buffer_data_0[1471:1464];
        layer4[54][39:32] = buffer_data_0[1479:1472];
        layer0[55][7:0] = buffer_data_4[1455:1448];
        layer0[55][15:8] = buffer_data_4[1463:1456];
        layer0[55][23:16] = buffer_data_4[1471:1464];
        layer0[55][31:24] = buffer_data_4[1479:1472];
        layer0[55][39:32] = buffer_data_4[1487:1480];
        layer1[55][7:0] = buffer_data_3[1455:1448];
        layer1[55][15:8] = buffer_data_3[1463:1456];
        layer1[55][23:16] = buffer_data_3[1471:1464];
        layer1[55][31:24] = buffer_data_3[1479:1472];
        layer1[55][39:32] = buffer_data_3[1487:1480];
        layer2[55][7:0] = buffer_data_2[1455:1448];
        layer2[55][15:8] = buffer_data_2[1463:1456];
        layer2[55][23:16] = buffer_data_2[1471:1464];
        layer2[55][31:24] = buffer_data_2[1479:1472];
        layer2[55][39:32] = buffer_data_2[1487:1480];
        layer3[55][7:0] = buffer_data_1[1455:1448];
        layer3[55][15:8] = buffer_data_1[1463:1456];
        layer3[55][23:16] = buffer_data_1[1471:1464];
        layer3[55][31:24] = buffer_data_1[1479:1472];
        layer3[55][39:32] = buffer_data_1[1487:1480];
        layer4[55][7:0] = buffer_data_0[1455:1448];
        layer4[55][15:8] = buffer_data_0[1463:1456];
        layer4[55][23:16] = buffer_data_0[1471:1464];
        layer4[55][31:24] = buffer_data_0[1479:1472];
        layer4[55][39:32] = buffer_data_0[1487:1480];
        layer0[56][7:0] = buffer_data_4[1463:1456];
        layer0[56][15:8] = buffer_data_4[1471:1464];
        layer0[56][23:16] = buffer_data_4[1479:1472];
        layer0[56][31:24] = buffer_data_4[1487:1480];
        layer0[56][39:32] = buffer_data_4[1495:1488];
        layer1[56][7:0] = buffer_data_3[1463:1456];
        layer1[56][15:8] = buffer_data_3[1471:1464];
        layer1[56][23:16] = buffer_data_3[1479:1472];
        layer1[56][31:24] = buffer_data_3[1487:1480];
        layer1[56][39:32] = buffer_data_3[1495:1488];
        layer2[56][7:0] = buffer_data_2[1463:1456];
        layer2[56][15:8] = buffer_data_2[1471:1464];
        layer2[56][23:16] = buffer_data_2[1479:1472];
        layer2[56][31:24] = buffer_data_2[1487:1480];
        layer2[56][39:32] = buffer_data_2[1495:1488];
        layer3[56][7:0] = buffer_data_1[1463:1456];
        layer3[56][15:8] = buffer_data_1[1471:1464];
        layer3[56][23:16] = buffer_data_1[1479:1472];
        layer3[56][31:24] = buffer_data_1[1487:1480];
        layer3[56][39:32] = buffer_data_1[1495:1488];
        layer4[56][7:0] = buffer_data_0[1463:1456];
        layer4[56][15:8] = buffer_data_0[1471:1464];
        layer4[56][23:16] = buffer_data_0[1479:1472];
        layer4[56][31:24] = buffer_data_0[1487:1480];
        layer4[56][39:32] = buffer_data_0[1495:1488];
        layer0[57][7:0] = buffer_data_4[1471:1464];
        layer0[57][15:8] = buffer_data_4[1479:1472];
        layer0[57][23:16] = buffer_data_4[1487:1480];
        layer0[57][31:24] = buffer_data_4[1495:1488];
        layer0[57][39:32] = buffer_data_4[1503:1496];
        layer1[57][7:0] = buffer_data_3[1471:1464];
        layer1[57][15:8] = buffer_data_3[1479:1472];
        layer1[57][23:16] = buffer_data_3[1487:1480];
        layer1[57][31:24] = buffer_data_3[1495:1488];
        layer1[57][39:32] = buffer_data_3[1503:1496];
        layer2[57][7:0] = buffer_data_2[1471:1464];
        layer2[57][15:8] = buffer_data_2[1479:1472];
        layer2[57][23:16] = buffer_data_2[1487:1480];
        layer2[57][31:24] = buffer_data_2[1495:1488];
        layer2[57][39:32] = buffer_data_2[1503:1496];
        layer3[57][7:0] = buffer_data_1[1471:1464];
        layer3[57][15:8] = buffer_data_1[1479:1472];
        layer3[57][23:16] = buffer_data_1[1487:1480];
        layer3[57][31:24] = buffer_data_1[1495:1488];
        layer3[57][39:32] = buffer_data_1[1503:1496];
        layer4[57][7:0] = buffer_data_0[1471:1464];
        layer4[57][15:8] = buffer_data_0[1479:1472];
        layer4[57][23:16] = buffer_data_0[1487:1480];
        layer4[57][31:24] = buffer_data_0[1495:1488];
        layer4[57][39:32] = buffer_data_0[1503:1496];
        layer0[58][7:0] = buffer_data_4[1479:1472];
        layer0[58][15:8] = buffer_data_4[1487:1480];
        layer0[58][23:16] = buffer_data_4[1495:1488];
        layer0[58][31:24] = buffer_data_4[1503:1496];
        layer0[58][39:32] = buffer_data_4[1511:1504];
        layer1[58][7:0] = buffer_data_3[1479:1472];
        layer1[58][15:8] = buffer_data_3[1487:1480];
        layer1[58][23:16] = buffer_data_3[1495:1488];
        layer1[58][31:24] = buffer_data_3[1503:1496];
        layer1[58][39:32] = buffer_data_3[1511:1504];
        layer2[58][7:0] = buffer_data_2[1479:1472];
        layer2[58][15:8] = buffer_data_2[1487:1480];
        layer2[58][23:16] = buffer_data_2[1495:1488];
        layer2[58][31:24] = buffer_data_2[1503:1496];
        layer2[58][39:32] = buffer_data_2[1511:1504];
        layer3[58][7:0] = buffer_data_1[1479:1472];
        layer3[58][15:8] = buffer_data_1[1487:1480];
        layer3[58][23:16] = buffer_data_1[1495:1488];
        layer3[58][31:24] = buffer_data_1[1503:1496];
        layer3[58][39:32] = buffer_data_1[1511:1504];
        layer4[58][7:0] = buffer_data_0[1479:1472];
        layer4[58][15:8] = buffer_data_0[1487:1480];
        layer4[58][23:16] = buffer_data_0[1495:1488];
        layer4[58][31:24] = buffer_data_0[1503:1496];
        layer4[58][39:32] = buffer_data_0[1511:1504];
        layer0[59][7:0] = buffer_data_4[1487:1480];
        layer0[59][15:8] = buffer_data_4[1495:1488];
        layer0[59][23:16] = buffer_data_4[1503:1496];
        layer0[59][31:24] = buffer_data_4[1511:1504];
        layer0[59][39:32] = buffer_data_4[1519:1512];
        layer1[59][7:0] = buffer_data_3[1487:1480];
        layer1[59][15:8] = buffer_data_3[1495:1488];
        layer1[59][23:16] = buffer_data_3[1503:1496];
        layer1[59][31:24] = buffer_data_3[1511:1504];
        layer1[59][39:32] = buffer_data_3[1519:1512];
        layer2[59][7:0] = buffer_data_2[1487:1480];
        layer2[59][15:8] = buffer_data_2[1495:1488];
        layer2[59][23:16] = buffer_data_2[1503:1496];
        layer2[59][31:24] = buffer_data_2[1511:1504];
        layer2[59][39:32] = buffer_data_2[1519:1512];
        layer3[59][7:0] = buffer_data_1[1487:1480];
        layer3[59][15:8] = buffer_data_1[1495:1488];
        layer3[59][23:16] = buffer_data_1[1503:1496];
        layer3[59][31:24] = buffer_data_1[1511:1504];
        layer3[59][39:32] = buffer_data_1[1519:1512];
        layer4[59][7:0] = buffer_data_0[1487:1480];
        layer4[59][15:8] = buffer_data_0[1495:1488];
        layer4[59][23:16] = buffer_data_0[1503:1496];
        layer4[59][31:24] = buffer_data_0[1511:1504];
        layer4[59][39:32] = buffer_data_0[1519:1512];
        layer0[60][7:0] = buffer_data_4[1495:1488];
        layer0[60][15:8] = buffer_data_4[1503:1496];
        layer0[60][23:16] = buffer_data_4[1511:1504];
        layer0[60][31:24] = buffer_data_4[1519:1512];
        layer0[60][39:32] = buffer_data_4[1527:1520];
        layer1[60][7:0] = buffer_data_3[1495:1488];
        layer1[60][15:8] = buffer_data_3[1503:1496];
        layer1[60][23:16] = buffer_data_3[1511:1504];
        layer1[60][31:24] = buffer_data_3[1519:1512];
        layer1[60][39:32] = buffer_data_3[1527:1520];
        layer2[60][7:0] = buffer_data_2[1495:1488];
        layer2[60][15:8] = buffer_data_2[1503:1496];
        layer2[60][23:16] = buffer_data_2[1511:1504];
        layer2[60][31:24] = buffer_data_2[1519:1512];
        layer2[60][39:32] = buffer_data_2[1527:1520];
        layer3[60][7:0] = buffer_data_1[1495:1488];
        layer3[60][15:8] = buffer_data_1[1503:1496];
        layer3[60][23:16] = buffer_data_1[1511:1504];
        layer3[60][31:24] = buffer_data_1[1519:1512];
        layer3[60][39:32] = buffer_data_1[1527:1520];
        layer4[60][7:0] = buffer_data_0[1495:1488];
        layer4[60][15:8] = buffer_data_0[1503:1496];
        layer4[60][23:16] = buffer_data_0[1511:1504];
        layer4[60][31:24] = buffer_data_0[1519:1512];
        layer4[60][39:32] = buffer_data_0[1527:1520];
        layer0[61][7:0] = buffer_data_4[1503:1496];
        layer0[61][15:8] = buffer_data_4[1511:1504];
        layer0[61][23:16] = buffer_data_4[1519:1512];
        layer0[61][31:24] = buffer_data_4[1527:1520];
        layer0[61][39:32] = buffer_data_4[1535:1528];
        layer1[61][7:0] = buffer_data_3[1503:1496];
        layer1[61][15:8] = buffer_data_3[1511:1504];
        layer1[61][23:16] = buffer_data_3[1519:1512];
        layer1[61][31:24] = buffer_data_3[1527:1520];
        layer1[61][39:32] = buffer_data_3[1535:1528];
        layer2[61][7:0] = buffer_data_2[1503:1496];
        layer2[61][15:8] = buffer_data_2[1511:1504];
        layer2[61][23:16] = buffer_data_2[1519:1512];
        layer2[61][31:24] = buffer_data_2[1527:1520];
        layer2[61][39:32] = buffer_data_2[1535:1528];
        layer3[61][7:0] = buffer_data_1[1503:1496];
        layer3[61][15:8] = buffer_data_1[1511:1504];
        layer3[61][23:16] = buffer_data_1[1519:1512];
        layer3[61][31:24] = buffer_data_1[1527:1520];
        layer3[61][39:32] = buffer_data_1[1535:1528];
        layer4[61][7:0] = buffer_data_0[1503:1496];
        layer4[61][15:8] = buffer_data_0[1511:1504];
        layer4[61][23:16] = buffer_data_0[1519:1512];
        layer4[61][31:24] = buffer_data_0[1527:1520];
        layer4[61][39:32] = buffer_data_0[1535:1528];
        layer0[62][7:0] = buffer_data_4[1511:1504];
        layer0[62][15:8] = buffer_data_4[1519:1512];
        layer0[62][23:16] = buffer_data_4[1527:1520];
        layer0[62][31:24] = buffer_data_4[1535:1528];
        layer0[62][39:32] = buffer_data_4[1543:1536];
        layer1[62][7:0] = buffer_data_3[1511:1504];
        layer1[62][15:8] = buffer_data_3[1519:1512];
        layer1[62][23:16] = buffer_data_3[1527:1520];
        layer1[62][31:24] = buffer_data_3[1535:1528];
        layer1[62][39:32] = buffer_data_3[1543:1536];
        layer2[62][7:0] = buffer_data_2[1511:1504];
        layer2[62][15:8] = buffer_data_2[1519:1512];
        layer2[62][23:16] = buffer_data_2[1527:1520];
        layer2[62][31:24] = buffer_data_2[1535:1528];
        layer2[62][39:32] = buffer_data_2[1543:1536];
        layer3[62][7:0] = buffer_data_1[1511:1504];
        layer3[62][15:8] = buffer_data_1[1519:1512];
        layer3[62][23:16] = buffer_data_1[1527:1520];
        layer3[62][31:24] = buffer_data_1[1535:1528];
        layer3[62][39:32] = buffer_data_1[1543:1536];
        layer4[62][7:0] = buffer_data_0[1511:1504];
        layer4[62][15:8] = buffer_data_0[1519:1512];
        layer4[62][23:16] = buffer_data_0[1527:1520];
        layer4[62][31:24] = buffer_data_0[1535:1528];
        layer4[62][39:32] = buffer_data_0[1543:1536];
        layer0[63][7:0] = buffer_data_4[1519:1512];
        layer0[63][15:8] = buffer_data_4[1527:1520];
        layer0[63][23:16] = buffer_data_4[1535:1528];
        layer0[63][31:24] = buffer_data_4[1543:1536];
        layer0[63][39:32] = buffer_data_4[1551:1544];
        layer1[63][7:0] = buffer_data_3[1519:1512];
        layer1[63][15:8] = buffer_data_3[1527:1520];
        layer1[63][23:16] = buffer_data_3[1535:1528];
        layer1[63][31:24] = buffer_data_3[1543:1536];
        layer1[63][39:32] = buffer_data_3[1551:1544];
        layer2[63][7:0] = buffer_data_2[1519:1512];
        layer2[63][15:8] = buffer_data_2[1527:1520];
        layer2[63][23:16] = buffer_data_2[1535:1528];
        layer2[63][31:24] = buffer_data_2[1543:1536];
        layer2[63][39:32] = buffer_data_2[1551:1544];
        layer3[63][7:0] = buffer_data_1[1519:1512];
        layer3[63][15:8] = buffer_data_1[1527:1520];
        layer3[63][23:16] = buffer_data_1[1535:1528];
        layer3[63][31:24] = buffer_data_1[1543:1536];
        layer3[63][39:32] = buffer_data_1[1551:1544];
        layer4[63][7:0] = buffer_data_0[1519:1512];
        layer4[63][15:8] = buffer_data_0[1527:1520];
        layer4[63][23:16] = buffer_data_0[1535:1528];
        layer4[63][31:24] = buffer_data_0[1543:1536];
        layer4[63][39:32] = buffer_data_0[1551:1544];
    end
    ST_GAUSSIAN_3: begin
        layer0[0][7:0] = buffer_data_4[1527:1520];
        layer0[0][15:8] = buffer_data_4[1535:1528];
        layer0[0][23:16] = buffer_data_4[1543:1536];
        layer0[0][31:24] = buffer_data_4[1551:1544];
        layer0[0][39:32] = buffer_data_4[1559:1552];
        layer1[0][7:0] = buffer_data_3[1527:1520];
        layer1[0][15:8] = buffer_data_3[1535:1528];
        layer1[0][23:16] = buffer_data_3[1543:1536];
        layer1[0][31:24] = buffer_data_3[1551:1544];
        layer1[0][39:32] = buffer_data_3[1559:1552];
        layer2[0][7:0] = buffer_data_2[1527:1520];
        layer2[0][15:8] = buffer_data_2[1535:1528];
        layer2[0][23:16] = buffer_data_2[1543:1536];
        layer2[0][31:24] = buffer_data_2[1551:1544];
        layer2[0][39:32] = buffer_data_2[1559:1552];
        layer3[0][7:0] = buffer_data_1[1527:1520];
        layer3[0][15:8] = buffer_data_1[1535:1528];
        layer3[0][23:16] = buffer_data_1[1543:1536];
        layer3[0][31:24] = buffer_data_1[1551:1544];
        layer3[0][39:32] = buffer_data_1[1559:1552];
        layer4[0][7:0] = buffer_data_0[1527:1520];
        layer4[0][15:8] = buffer_data_0[1535:1528];
        layer4[0][23:16] = buffer_data_0[1543:1536];
        layer4[0][31:24] = buffer_data_0[1551:1544];
        layer4[0][39:32] = buffer_data_0[1559:1552];
        layer0[1][7:0] = buffer_data_4[1535:1528];
        layer0[1][15:8] = buffer_data_4[1543:1536];
        layer0[1][23:16] = buffer_data_4[1551:1544];
        layer0[1][31:24] = buffer_data_4[1559:1552];
        layer0[1][39:32] = buffer_data_4[1567:1560];
        layer1[1][7:0] = buffer_data_3[1535:1528];
        layer1[1][15:8] = buffer_data_3[1543:1536];
        layer1[1][23:16] = buffer_data_3[1551:1544];
        layer1[1][31:24] = buffer_data_3[1559:1552];
        layer1[1][39:32] = buffer_data_3[1567:1560];
        layer2[1][7:0] = buffer_data_2[1535:1528];
        layer2[1][15:8] = buffer_data_2[1543:1536];
        layer2[1][23:16] = buffer_data_2[1551:1544];
        layer2[1][31:24] = buffer_data_2[1559:1552];
        layer2[1][39:32] = buffer_data_2[1567:1560];
        layer3[1][7:0] = buffer_data_1[1535:1528];
        layer3[1][15:8] = buffer_data_1[1543:1536];
        layer3[1][23:16] = buffer_data_1[1551:1544];
        layer3[1][31:24] = buffer_data_1[1559:1552];
        layer3[1][39:32] = buffer_data_1[1567:1560];
        layer4[1][7:0] = buffer_data_0[1535:1528];
        layer4[1][15:8] = buffer_data_0[1543:1536];
        layer4[1][23:16] = buffer_data_0[1551:1544];
        layer4[1][31:24] = buffer_data_0[1559:1552];
        layer4[1][39:32] = buffer_data_0[1567:1560];
        layer0[2][7:0] = buffer_data_4[1543:1536];
        layer0[2][15:8] = buffer_data_4[1551:1544];
        layer0[2][23:16] = buffer_data_4[1559:1552];
        layer0[2][31:24] = buffer_data_4[1567:1560];
        layer0[2][39:32] = buffer_data_4[1575:1568];
        layer1[2][7:0] = buffer_data_3[1543:1536];
        layer1[2][15:8] = buffer_data_3[1551:1544];
        layer1[2][23:16] = buffer_data_3[1559:1552];
        layer1[2][31:24] = buffer_data_3[1567:1560];
        layer1[2][39:32] = buffer_data_3[1575:1568];
        layer2[2][7:0] = buffer_data_2[1543:1536];
        layer2[2][15:8] = buffer_data_2[1551:1544];
        layer2[2][23:16] = buffer_data_2[1559:1552];
        layer2[2][31:24] = buffer_data_2[1567:1560];
        layer2[2][39:32] = buffer_data_2[1575:1568];
        layer3[2][7:0] = buffer_data_1[1543:1536];
        layer3[2][15:8] = buffer_data_1[1551:1544];
        layer3[2][23:16] = buffer_data_1[1559:1552];
        layer3[2][31:24] = buffer_data_1[1567:1560];
        layer3[2][39:32] = buffer_data_1[1575:1568];
        layer4[2][7:0] = buffer_data_0[1543:1536];
        layer4[2][15:8] = buffer_data_0[1551:1544];
        layer4[2][23:16] = buffer_data_0[1559:1552];
        layer4[2][31:24] = buffer_data_0[1567:1560];
        layer4[2][39:32] = buffer_data_0[1575:1568];
        layer0[3][7:0] = buffer_data_4[1551:1544];
        layer0[3][15:8] = buffer_data_4[1559:1552];
        layer0[3][23:16] = buffer_data_4[1567:1560];
        layer0[3][31:24] = buffer_data_4[1575:1568];
        layer0[3][39:32] = buffer_data_4[1583:1576];
        layer1[3][7:0] = buffer_data_3[1551:1544];
        layer1[3][15:8] = buffer_data_3[1559:1552];
        layer1[3][23:16] = buffer_data_3[1567:1560];
        layer1[3][31:24] = buffer_data_3[1575:1568];
        layer1[3][39:32] = buffer_data_3[1583:1576];
        layer2[3][7:0] = buffer_data_2[1551:1544];
        layer2[3][15:8] = buffer_data_2[1559:1552];
        layer2[3][23:16] = buffer_data_2[1567:1560];
        layer2[3][31:24] = buffer_data_2[1575:1568];
        layer2[3][39:32] = buffer_data_2[1583:1576];
        layer3[3][7:0] = buffer_data_1[1551:1544];
        layer3[3][15:8] = buffer_data_1[1559:1552];
        layer3[3][23:16] = buffer_data_1[1567:1560];
        layer3[3][31:24] = buffer_data_1[1575:1568];
        layer3[3][39:32] = buffer_data_1[1583:1576];
        layer4[3][7:0] = buffer_data_0[1551:1544];
        layer4[3][15:8] = buffer_data_0[1559:1552];
        layer4[3][23:16] = buffer_data_0[1567:1560];
        layer4[3][31:24] = buffer_data_0[1575:1568];
        layer4[3][39:32] = buffer_data_0[1583:1576];
        layer0[4][7:0] = buffer_data_4[1559:1552];
        layer0[4][15:8] = buffer_data_4[1567:1560];
        layer0[4][23:16] = buffer_data_4[1575:1568];
        layer0[4][31:24] = buffer_data_4[1583:1576];
        layer0[4][39:32] = buffer_data_4[1591:1584];
        layer1[4][7:0] = buffer_data_3[1559:1552];
        layer1[4][15:8] = buffer_data_3[1567:1560];
        layer1[4][23:16] = buffer_data_3[1575:1568];
        layer1[4][31:24] = buffer_data_3[1583:1576];
        layer1[4][39:32] = buffer_data_3[1591:1584];
        layer2[4][7:0] = buffer_data_2[1559:1552];
        layer2[4][15:8] = buffer_data_2[1567:1560];
        layer2[4][23:16] = buffer_data_2[1575:1568];
        layer2[4][31:24] = buffer_data_2[1583:1576];
        layer2[4][39:32] = buffer_data_2[1591:1584];
        layer3[4][7:0] = buffer_data_1[1559:1552];
        layer3[4][15:8] = buffer_data_1[1567:1560];
        layer3[4][23:16] = buffer_data_1[1575:1568];
        layer3[4][31:24] = buffer_data_1[1583:1576];
        layer3[4][39:32] = buffer_data_1[1591:1584];
        layer4[4][7:0] = buffer_data_0[1559:1552];
        layer4[4][15:8] = buffer_data_0[1567:1560];
        layer4[4][23:16] = buffer_data_0[1575:1568];
        layer4[4][31:24] = buffer_data_0[1583:1576];
        layer4[4][39:32] = buffer_data_0[1591:1584];
        layer0[5][7:0] = buffer_data_4[1567:1560];
        layer0[5][15:8] = buffer_data_4[1575:1568];
        layer0[5][23:16] = buffer_data_4[1583:1576];
        layer0[5][31:24] = buffer_data_4[1591:1584];
        layer0[5][39:32] = buffer_data_4[1599:1592];
        layer1[5][7:0] = buffer_data_3[1567:1560];
        layer1[5][15:8] = buffer_data_3[1575:1568];
        layer1[5][23:16] = buffer_data_3[1583:1576];
        layer1[5][31:24] = buffer_data_3[1591:1584];
        layer1[5][39:32] = buffer_data_3[1599:1592];
        layer2[5][7:0] = buffer_data_2[1567:1560];
        layer2[5][15:8] = buffer_data_2[1575:1568];
        layer2[5][23:16] = buffer_data_2[1583:1576];
        layer2[5][31:24] = buffer_data_2[1591:1584];
        layer2[5][39:32] = buffer_data_2[1599:1592];
        layer3[5][7:0] = buffer_data_1[1567:1560];
        layer3[5][15:8] = buffer_data_1[1575:1568];
        layer3[5][23:16] = buffer_data_1[1583:1576];
        layer3[5][31:24] = buffer_data_1[1591:1584];
        layer3[5][39:32] = buffer_data_1[1599:1592];
        layer4[5][7:0] = buffer_data_0[1567:1560];
        layer4[5][15:8] = buffer_data_0[1575:1568];
        layer4[5][23:16] = buffer_data_0[1583:1576];
        layer4[5][31:24] = buffer_data_0[1591:1584];
        layer4[5][39:32] = buffer_data_0[1599:1592];
        layer0[6][7:0] = buffer_data_4[1575:1568];
        layer0[6][15:8] = buffer_data_4[1583:1576];
        layer0[6][23:16] = buffer_data_4[1591:1584];
        layer0[6][31:24] = buffer_data_4[1599:1592];
        layer0[6][39:32] = buffer_data_4[1607:1600];
        layer1[6][7:0] = buffer_data_3[1575:1568];
        layer1[6][15:8] = buffer_data_3[1583:1576];
        layer1[6][23:16] = buffer_data_3[1591:1584];
        layer1[6][31:24] = buffer_data_3[1599:1592];
        layer1[6][39:32] = buffer_data_3[1607:1600];
        layer2[6][7:0] = buffer_data_2[1575:1568];
        layer2[6][15:8] = buffer_data_2[1583:1576];
        layer2[6][23:16] = buffer_data_2[1591:1584];
        layer2[6][31:24] = buffer_data_2[1599:1592];
        layer2[6][39:32] = buffer_data_2[1607:1600];
        layer3[6][7:0] = buffer_data_1[1575:1568];
        layer3[6][15:8] = buffer_data_1[1583:1576];
        layer3[6][23:16] = buffer_data_1[1591:1584];
        layer3[6][31:24] = buffer_data_1[1599:1592];
        layer3[6][39:32] = buffer_data_1[1607:1600];
        layer4[6][7:0] = buffer_data_0[1575:1568];
        layer4[6][15:8] = buffer_data_0[1583:1576];
        layer4[6][23:16] = buffer_data_0[1591:1584];
        layer4[6][31:24] = buffer_data_0[1599:1592];
        layer4[6][39:32] = buffer_data_0[1607:1600];
        layer0[7][7:0] = buffer_data_4[1583:1576];
        layer0[7][15:8] = buffer_data_4[1591:1584];
        layer0[7][23:16] = buffer_data_4[1599:1592];
        layer0[7][31:24] = buffer_data_4[1607:1600];
        layer0[7][39:32] = buffer_data_4[1615:1608];
        layer1[7][7:0] = buffer_data_3[1583:1576];
        layer1[7][15:8] = buffer_data_3[1591:1584];
        layer1[7][23:16] = buffer_data_3[1599:1592];
        layer1[7][31:24] = buffer_data_3[1607:1600];
        layer1[7][39:32] = buffer_data_3[1615:1608];
        layer2[7][7:0] = buffer_data_2[1583:1576];
        layer2[7][15:8] = buffer_data_2[1591:1584];
        layer2[7][23:16] = buffer_data_2[1599:1592];
        layer2[7][31:24] = buffer_data_2[1607:1600];
        layer2[7][39:32] = buffer_data_2[1615:1608];
        layer3[7][7:0] = buffer_data_1[1583:1576];
        layer3[7][15:8] = buffer_data_1[1591:1584];
        layer3[7][23:16] = buffer_data_1[1599:1592];
        layer3[7][31:24] = buffer_data_1[1607:1600];
        layer3[7][39:32] = buffer_data_1[1615:1608];
        layer4[7][7:0] = buffer_data_0[1583:1576];
        layer4[7][15:8] = buffer_data_0[1591:1584];
        layer4[7][23:16] = buffer_data_0[1599:1592];
        layer4[7][31:24] = buffer_data_0[1607:1600];
        layer4[7][39:32] = buffer_data_0[1615:1608];
        layer0[8][7:0] = buffer_data_4[1591:1584];
        layer0[8][15:8] = buffer_data_4[1599:1592];
        layer0[8][23:16] = buffer_data_4[1607:1600];
        layer0[8][31:24] = buffer_data_4[1615:1608];
        layer0[8][39:32] = buffer_data_4[1623:1616];
        layer1[8][7:0] = buffer_data_3[1591:1584];
        layer1[8][15:8] = buffer_data_3[1599:1592];
        layer1[8][23:16] = buffer_data_3[1607:1600];
        layer1[8][31:24] = buffer_data_3[1615:1608];
        layer1[8][39:32] = buffer_data_3[1623:1616];
        layer2[8][7:0] = buffer_data_2[1591:1584];
        layer2[8][15:8] = buffer_data_2[1599:1592];
        layer2[8][23:16] = buffer_data_2[1607:1600];
        layer2[8][31:24] = buffer_data_2[1615:1608];
        layer2[8][39:32] = buffer_data_2[1623:1616];
        layer3[8][7:0] = buffer_data_1[1591:1584];
        layer3[8][15:8] = buffer_data_1[1599:1592];
        layer3[8][23:16] = buffer_data_1[1607:1600];
        layer3[8][31:24] = buffer_data_1[1615:1608];
        layer3[8][39:32] = buffer_data_1[1623:1616];
        layer4[8][7:0] = buffer_data_0[1591:1584];
        layer4[8][15:8] = buffer_data_0[1599:1592];
        layer4[8][23:16] = buffer_data_0[1607:1600];
        layer4[8][31:24] = buffer_data_0[1615:1608];
        layer4[8][39:32] = buffer_data_0[1623:1616];
        layer0[9][7:0] = buffer_data_4[1599:1592];
        layer0[9][15:8] = buffer_data_4[1607:1600];
        layer0[9][23:16] = buffer_data_4[1615:1608];
        layer0[9][31:24] = buffer_data_4[1623:1616];
        layer0[9][39:32] = buffer_data_4[1631:1624];
        layer1[9][7:0] = buffer_data_3[1599:1592];
        layer1[9][15:8] = buffer_data_3[1607:1600];
        layer1[9][23:16] = buffer_data_3[1615:1608];
        layer1[9][31:24] = buffer_data_3[1623:1616];
        layer1[9][39:32] = buffer_data_3[1631:1624];
        layer2[9][7:0] = buffer_data_2[1599:1592];
        layer2[9][15:8] = buffer_data_2[1607:1600];
        layer2[9][23:16] = buffer_data_2[1615:1608];
        layer2[9][31:24] = buffer_data_2[1623:1616];
        layer2[9][39:32] = buffer_data_2[1631:1624];
        layer3[9][7:0] = buffer_data_1[1599:1592];
        layer3[9][15:8] = buffer_data_1[1607:1600];
        layer3[9][23:16] = buffer_data_1[1615:1608];
        layer3[9][31:24] = buffer_data_1[1623:1616];
        layer3[9][39:32] = buffer_data_1[1631:1624];
        layer4[9][7:0] = buffer_data_0[1599:1592];
        layer4[9][15:8] = buffer_data_0[1607:1600];
        layer4[9][23:16] = buffer_data_0[1615:1608];
        layer4[9][31:24] = buffer_data_0[1623:1616];
        layer4[9][39:32] = buffer_data_0[1631:1624];
        layer0[10][7:0] = buffer_data_4[1607:1600];
        layer0[10][15:8] = buffer_data_4[1615:1608];
        layer0[10][23:16] = buffer_data_4[1623:1616];
        layer0[10][31:24] = buffer_data_4[1631:1624];
        layer0[10][39:32] = buffer_data_4[1639:1632];
        layer1[10][7:0] = buffer_data_3[1607:1600];
        layer1[10][15:8] = buffer_data_3[1615:1608];
        layer1[10][23:16] = buffer_data_3[1623:1616];
        layer1[10][31:24] = buffer_data_3[1631:1624];
        layer1[10][39:32] = buffer_data_3[1639:1632];
        layer2[10][7:0] = buffer_data_2[1607:1600];
        layer2[10][15:8] = buffer_data_2[1615:1608];
        layer2[10][23:16] = buffer_data_2[1623:1616];
        layer2[10][31:24] = buffer_data_2[1631:1624];
        layer2[10][39:32] = buffer_data_2[1639:1632];
        layer3[10][7:0] = buffer_data_1[1607:1600];
        layer3[10][15:8] = buffer_data_1[1615:1608];
        layer3[10][23:16] = buffer_data_1[1623:1616];
        layer3[10][31:24] = buffer_data_1[1631:1624];
        layer3[10][39:32] = buffer_data_1[1639:1632];
        layer4[10][7:0] = buffer_data_0[1607:1600];
        layer4[10][15:8] = buffer_data_0[1615:1608];
        layer4[10][23:16] = buffer_data_0[1623:1616];
        layer4[10][31:24] = buffer_data_0[1631:1624];
        layer4[10][39:32] = buffer_data_0[1639:1632];
        layer0[11][7:0] = buffer_data_4[1615:1608];
        layer0[11][15:8] = buffer_data_4[1623:1616];
        layer0[11][23:16] = buffer_data_4[1631:1624];
        layer0[11][31:24] = buffer_data_4[1639:1632];
        layer0[11][39:32] = buffer_data_4[1647:1640];
        layer1[11][7:0] = buffer_data_3[1615:1608];
        layer1[11][15:8] = buffer_data_3[1623:1616];
        layer1[11][23:16] = buffer_data_3[1631:1624];
        layer1[11][31:24] = buffer_data_3[1639:1632];
        layer1[11][39:32] = buffer_data_3[1647:1640];
        layer2[11][7:0] = buffer_data_2[1615:1608];
        layer2[11][15:8] = buffer_data_2[1623:1616];
        layer2[11][23:16] = buffer_data_2[1631:1624];
        layer2[11][31:24] = buffer_data_2[1639:1632];
        layer2[11][39:32] = buffer_data_2[1647:1640];
        layer3[11][7:0] = buffer_data_1[1615:1608];
        layer3[11][15:8] = buffer_data_1[1623:1616];
        layer3[11][23:16] = buffer_data_1[1631:1624];
        layer3[11][31:24] = buffer_data_1[1639:1632];
        layer3[11][39:32] = buffer_data_1[1647:1640];
        layer4[11][7:0] = buffer_data_0[1615:1608];
        layer4[11][15:8] = buffer_data_0[1623:1616];
        layer4[11][23:16] = buffer_data_0[1631:1624];
        layer4[11][31:24] = buffer_data_0[1639:1632];
        layer4[11][39:32] = buffer_data_0[1647:1640];
        layer0[12][7:0] = buffer_data_4[1623:1616];
        layer0[12][15:8] = buffer_data_4[1631:1624];
        layer0[12][23:16] = buffer_data_4[1639:1632];
        layer0[12][31:24] = buffer_data_4[1647:1640];
        layer0[12][39:32] = buffer_data_4[1655:1648];
        layer1[12][7:0] = buffer_data_3[1623:1616];
        layer1[12][15:8] = buffer_data_3[1631:1624];
        layer1[12][23:16] = buffer_data_3[1639:1632];
        layer1[12][31:24] = buffer_data_3[1647:1640];
        layer1[12][39:32] = buffer_data_3[1655:1648];
        layer2[12][7:0] = buffer_data_2[1623:1616];
        layer2[12][15:8] = buffer_data_2[1631:1624];
        layer2[12][23:16] = buffer_data_2[1639:1632];
        layer2[12][31:24] = buffer_data_2[1647:1640];
        layer2[12][39:32] = buffer_data_2[1655:1648];
        layer3[12][7:0] = buffer_data_1[1623:1616];
        layer3[12][15:8] = buffer_data_1[1631:1624];
        layer3[12][23:16] = buffer_data_1[1639:1632];
        layer3[12][31:24] = buffer_data_1[1647:1640];
        layer3[12][39:32] = buffer_data_1[1655:1648];
        layer4[12][7:0] = buffer_data_0[1623:1616];
        layer4[12][15:8] = buffer_data_0[1631:1624];
        layer4[12][23:16] = buffer_data_0[1639:1632];
        layer4[12][31:24] = buffer_data_0[1647:1640];
        layer4[12][39:32] = buffer_data_0[1655:1648];
        layer0[13][7:0] = buffer_data_4[1631:1624];
        layer0[13][15:8] = buffer_data_4[1639:1632];
        layer0[13][23:16] = buffer_data_4[1647:1640];
        layer0[13][31:24] = buffer_data_4[1655:1648];
        layer0[13][39:32] = buffer_data_4[1663:1656];
        layer1[13][7:0] = buffer_data_3[1631:1624];
        layer1[13][15:8] = buffer_data_3[1639:1632];
        layer1[13][23:16] = buffer_data_3[1647:1640];
        layer1[13][31:24] = buffer_data_3[1655:1648];
        layer1[13][39:32] = buffer_data_3[1663:1656];
        layer2[13][7:0] = buffer_data_2[1631:1624];
        layer2[13][15:8] = buffer_data_2[1639:1632];
        layer2[13][23:16] = buffer_data_2[1647:1640];
        layer2[13][31:24] = buffer_data_2[1655:1648];
        layer2[13][39:32] = buffer_data_2[1663:1656];
        layer3[13][7:0] = buffer_data_1[1631:1624];
        layer3[13][15:8] = buffer_data_1[1639:1632];
        layer3[13][23:16] = buffer_data_1[1647:1640];
        layer3[13][31:24] = buffer_data_1[1655:1648];
        layer3[13][39:32] = buffer_data_1[1663:1656];
        layer4[13][7:0] = buffer_data_0[1631:1624];
        layer4[13][15:8] = buffer_data_0[1639:1632];
        layer4[13][23:16] = buffer_data_0[1647:1640];
        layer4[13][31:24] = buffer_data_0[1655:1648];
        layer4[13][39:32] = buffer_data_0[1663:1656];
        layer0[14][7:0] = buffer_data_4[1639:1632];
        layer0[14][15:8] = buffer_data_4[1647:1640];
        layer0[14][23:16] = buffer_data_4[1655:1648];
        layer0[14][31:24] = buffer_data_4[1663:1656];
        layer0[14][39:32] = buffer_data_4[1671:1664];
        layer1[14][7:0] = buffer_data_3[1639:1632];
        layer1[14][15:8] = buffer_data_3[1647:1640];
        layer1[14][23:16] = buffer_data_3[1655:1648];
        layer1[14][31:24] = buffer_data_3[1663:1656];
        layer1[14][39:32] = buffer_data_3[1671:1664];
        layer2[14][7:0] = buffer_data_2[1639:1632];
        layer2[14][15:8] = buffer_data_2[1647:1640];
        layer2[14][23:16] = buffer_data_2[1655:1648];
        layer2[14][31:24] = buffer_data_2[1663:1656];
        layer2[14][39:32] = buffer_data_2[1671:1664];
        layer3[14][7:0] = buffer_data_1[1639:1632];
        layer3[14][15:8] = buffer_data_1[1647:1640];
        layer3[14][23:16] = buffer_data_1[1655:1648];
        layer3[14][31:24] = buffer_data_1[1663:1656];
        layer3[14][39:32] = buffer_data_1[1671:1664];
        layer4[14][7:0] = buffer_data_0[1639:1632];
        layer4[14][15:8] = buffer_data_0[1647:1640];
        layer4[14][23:16] = buffer_data_0[1655:1648];
        layer4[14][31:24] = buffer_data_0[1663:1656];
        layer4[14][39:32] = buffer_data_0[1671:1664];
        layer0[15][7:0] = buffer_data_4[1647:1640];
        layer0[15][15:8] = buffer_data_4[1655:1648];
        layer0[15][23:16] = buffer_data_4[1663:1656];
        layer0[15][31:24] = buffer_data_4[1671:1664];
        layer0[15][39:32] = buffer_data_4[1679:1672];
        layer1[15][7:0] = buffer_data_3[1647:1640];
        layer1[15][15:8] = buffer_data_3[1655:1648];
        layer1[15][23:16] = buffer_data_3[1663:1656];
        layer1[15][31:24] = buffer_data_3[1671:1664];
        layer1[15][39:32] = buffer_data_3[1679:1672];
        layer2[15][7:0] = buffer_data_2[1647:1640];
        layer2[15][15:8] = buffer_data_2[1655:1648];
        layer2[15][23:16] = buffer_data_2[1663:1656];
        layer2[15][31:24] = buffer_data_2[1671:1664];
        layer2[15][39:32] = buffer_data_2[1679:1672];
        layer3[15][7:0] = buffer_data_1[1647:1640];
        layer3[15][15:8] = buffer_data_1[1655:1648];
        layer3[15][23:16] = buffer_data_1[1663:1656];
        layer3[15][31:24] = buffer_data_1[1671:1664];
        layer3[15][39:32] = buffer_data_1[1679:1672];
        layer4[15][7:0] = buffer_data_0[1647:1640];
        layer4[15][15:8] = buffer_data_0[1655:1648];
        layer4[15][23:16] = buffer_data_0[1663:1656];
        layer4[15][31:24] = buffer_data_0[1671:1664];
        layer4[15][39:32] = buffer_data_0[1679:1672];
        layer0[16][7:0] = buffer_data_4[1655:1648];
        layer0[16][15:8] = buffer_data_4[1663:1656];
        layer0[16][23:16] = buffer_data_4[1671:1664];
        layer0[16][31:24] = buffer_data_4[1679:1672];
        layer0[16][39:32] = buffer_data_4[1687:1680];
        layer1[16][7:0] = buffer_data_3[1655:1648];
        layer1[16][15:8] = buffer_data_3[1663:1656];
        layer1[16][23:16] = buffer_data_3[1671:1664];
        layer1[16][31:24] = buffer_data_3[1679:1672];
        layer1[16][39:32] = buffer_data_3[1687:1680];
        layer2[16][7:0] = buffer_data_2[1655:1648];
        layer2[16][15:8] = buffer_data_2[1663:1656];
        layer2[16][23:16] = buffer_data_2[1671:1664];
        layer2[16][31:24] = buffer_data_2[1679:1672];
        layer2[16][39:32] = buffer_data_2[1687:1680];
        layer3[16][7:0] = buffer_data_1[1655:1648];
        layer3[16][15:8] = buffer_data_1[1663:1656];
        layer3[16][23:16] = buffer_data_1[1671:1664];
        layer3[16][31:24] = buffer_data_1[1679:1672];
        layer3[16][39:32] = buffer_data_1[1687:1680];
        layer4[16][7:0] = buffer_data_0[1655:1648];
        layer4[16][15:8] = buffer_data_0[1663:1656];
        layer4[16][23:16] = buffer_data_0[1671:1664];
        layer4[16][31:24] = buffer_data_0[1679:1672];
        layer4[16][39:32] = buffer_data_0[1687:1680];
        layer0[17][7:0] = buffer_data_4[1663:1656];
        layer0[17][15:8] = buffer_data_4[1671:1664];
        layer0[17][23:16] = buffer_data_4[1679:1672];
        layer0[17][31:24] = buffer_data_4[1687:1680];
        layer0[17][39:32] = buffer_data_4[1695:1688];
        layer1[17][7:0] = buffer_data_3[1663:1656];
        layer1[17][15:8] = buffer_data_3[1671:1664];
        layer1[17][23:16] = buffer_data_3[1679:1672];
        layer1[17][31:24] = buffer_data_3[1687:1680];
        layer1[17][39:32] = buffer_data_3[1695:1688];
        layer2[17][7:0] = buffer_data_2[1663:1656];
        layer2[17][15:8] = buffer_data_2[1671:1664];
        layer2[17][23:16] = buffer_data_2[1679:1672];
        layer2[17][31:24] = buffer_data_2[1687:1680];
        layer2[17][39:32] = buffer_data_2[1695:1688];
        layer3[17][7:0] = buffer_data_1[1663:1656];
        layer3[17][15:8] = buffer_data_1[1671:1664];
        layer3[17][23:16] = buffer_data_1[1679:1672];
        layer3[17][31:24] = buffer_data_1[1687:1680];
        layer3[17][39:32] = buffer_data_1[1695:1688];
        layer4[17][7:0] = buffer_data_0[1663:1656];
        layer4[17][15:8] = buffer_data_0[1671:1664];
        layer4[17][23:16] = buffer_data_0[1679:1672];
        layer4[17][31:24] = buffer_data_0[1687:1680];
        layer4[17][39:32] = buffer_data_0[1695:1688];
        layer0[18][7:0] = buffer_data_4[1671:1664];
        layer0[18][15:8] = buffer_data_4[1679:1672];
        layer0[18][23:16] = buffer_data_4[1687:1680];
        layer0[18][31:24] = buffer_data_4[1695:1688];
        layer0[18][39:32] = buffer_data_4[1703:1696];
        layer1[18][7:0] = buffer_data_3[1671:1664];
        layer1[18][15:8] = buffer_data_3[1679:1672];
        layer1[18][23:16] = buffer_data_3[1687:1680];
        layer1[18][31:24] = buffer_data_3[1695:1688];
        layer1[18][39:32] = buffer_data_3[1703:1696];
        layer2[18][7:0] = buffer_data_2[1671:1664];
        layer2[18][15:8] = buffer_data_2[1679:1672];
        layer2[18][23:16] = buffer_data_2[1687:1680];
        layer2[18][31:24] = buffer_data_2[1695:1688];
        layer2[18][39:32] = buffer_data_2[1703:1696];
        layer3[18][7:0] = buffer_data_1[1671:1664];
        layer3[18][15:8] = buffer_data_1[1679:1672];
        layer3[18][23:16] = buffer_data_1[1687:1680];
        layer3[18][31:24] = buffer_data_1[1695:1688];
        layer3[18][39:32] = buffer_data_1[1703:1696];
        layer4[18][7:0] = buffer_data_0[1671:1664];
        layer4[18][15:8] = buffer_data_0[1679:1672];
        layer4[18][23:16] = buffer_data_0[1687:1680];
        layer4[18][31:24] = buffer_data_0[1695:1688];
        layer4[18][39:32] = buffer_data_0[1703:1696];
        layer0[19][7:0] = buffer_data_4[1679:1672];
        layer0[19][15:8] = buffer_data_4[1687:1680];
        layer0[19][23:16] = buffer_data_4[1695:1688];
        layer0[19][31:24] = buffer_data_4[1703:1696];
        layer0[19][39:32] = buffer_data_4[1711:1704];
        layer1[19][7:0] = buffer_data_3[1679:1672];
        layer1[19][15:8] = buffer_data_3[1687:1680];
        layer1[19][23:16] = buffer_data_3[1695:1688];
        layer1[19][31:24] = buffer_data_3[1703:1696];
        layer1[19][39:32] = buffer_data_3[1711:1704];
        layer2[19][7:0] = buffer_data_2[1679:1672];
        layer2[19][15:8] = buffer_data_2[1687:1680];
        layer2[19][23:16] = buffer_data_2[1695:1688];
        layer2[19][31:24] = buffer_data_2[1703:1696];
        layer2[19][39:32] = buffer_data_2[1711:1704];
        layer3[19][7:0] = buffer_data_1[1679:1672];
        layer3[19][15:8] = buffer_data_1[1687:1680];
        layer3[19][23:16] = buffer_data_1[1695:1688];
        layer3[19][31:24] = buffer_data_1[1703:1696];
        layer3[19][39:32] = buffer_data_1[1711:1704];
        layer4[19][7:0] = buffer_data_0[1679:1672];
        layer4[19][15:8] = buffer_data_0[1687:1680];
        layer4[19][23:16] = buffer_data_0[1695:1688];
        layer4[19][31:24] = buffer_data_0[1703:1696];
        layer4[19][39:32] = buffer_data_0[1711:1704];
        layer0[20][7:0] = buffer_data_4[1687:1680];
        layer0[20][15:8] = buffer_data_4[1695:1688];
        layer0[20][23:16] = buffer_data_4[1703:1696];
        layer0[20][31:24] = buffer_data_4[1711:1704];
        layer0[20][39:32] = buffer_data_4[1719:1712];
        layer1[20][7:0] = buffer_data_3[1687:1680];
        layer1[20][15:8] = buffer_data_3[1695:1688];
        layer1[20][23:16] = buffer_data_3[1703:1696];
        layer1[20][31:24] = buffer_data_3[1711:1704];
        layer1[20][39:32] = buffer_data_3[1719:1712];
        layer2[20][7:0] = buffer_data_2[1687:1680];
        layer2[20][15:8] = buffer_data_2[1695:1688];
        layer2[20][23:16] = buffer_data_2[1703:1696];
        layer2[20][31:24] = buffer_data_2[1711:1704];
        layer2[20][39:32] = buffer_data_2[1719:1712];
        layer3[20][7:0] = buffer_data_1[1687:1680];
        layer3[20][15:8] = buffer_data_1[1695:1688];
        layer3[20][23:16] = buffer_data_1[1703:1696];
        layer3[20][31:24] = buffer_data_1[1711:1704];
        layer3[20][39:32] = buffer_data_1[1719:1712];
        layer4[20][7:0] = buffer_data_0[1687:1680];
        layer4[20][15:8] = buffer_data_0[1695:1688];
        layer4[20][23:16] = buffer_data_0[1703:1696];
        layer4[20][31:24] = buffer_data_0[1711:1704];
        layer4[20][39:32] = buffer_data_0[1719:1712];
        layer0[21][7:0] = buffer_data_4[1695:1688];
        layer0[21][15:8] = buffer_data_4[1703:1696];
        layer0[21][23:16] = buffer_data_4[1711:1704];
        layer0[21][31:24] = buffer_data_4[1719:1712];
        layer0[21][39:32] = buffer_data_4[1727:1720];
        layer1[21][7:0] = buffer_data_3[1695:1688];
        layer1[21][15:8] = buffer_data_3[1703:1696];
        layer1[21][23:16] = buffer_data_3[1711:1704];
        layer1[21][31:24] = buffer_data_3[1719:1712];
        layer1[21][39:32] = buffer_data_3[1727:1720];
        layer2[21][7:0] = buffer_data_2[1695:1688];
        layer2[21][15:8] = buffer_data_2[1703:1696];
        layer2[21][23:16] = buffer_data_2[1711:1704];
        layer2[21][31:24] = buffer_data_2[1719:1712];
        layer2[21][39:32] = buffer_data_2[1727:1720];
        layer3[21][7:0] = buffer_data_1[1695:1688];
        layer3[21][15:8] = buffer_data_1[1703:1696];
        layer3[21][23:16] = buffer_data_1[1711:1704];
        layer3[21][31:24] = buffer_data_1[1719:1712];
        layer3[21][39:32] = buffer_data_1[1727:1720];
        layer4[21][7:0] = buffer_data_0[1695:1688];
        layer4[21][15:8] = buffer_data_0[1703:1696];
        layer4[21][23:16] = buffer_data_0[1711:1704];
        layer4[21][31:24] = buffer_data_0[1719:1712];
        layer4[21][39:32] = buffer_data_0[1727:1720];
        layer0[22][7:0] = buffer_data_4[1703:1696];
        layer0[22][15:8] = buffer_data_4[1711:1704];
        layer0[22][23:16] = buffer_data_4[1719:1712];
        layer0[22][31:24] = buffer_data_4[1727:1720];
        layer0[22][39:32] = buffer_data_4[1735:1728];
        layer1[22][7:0] = buffer_data_3[1703:1696];
        layer1[22][15:8] = buffer_data_3[1711:1704];
        layer1[22][23:16] = buffer_data_3[1719:1712];
        layer1[22][31:24] = buffer_data_3[1727:1720];
        layer1[22][39:32] = buffer_data_3[1735:1728];
        layer2[22][7:0] = buffer_data_2[1703:1696];
        layer2[22][15:8] = buffer_data_2[1711:1704];
        layer2[22][23:16] = buffer_data_2[1719:1712];
        layer2[22][31:24] = buffer_data_2[1727:1720];
        layer2[22][39:32] = buffer_data_2[1735:1728];
        layer3[22][7:0] = buffer_data_1[1703:1696];
        layer3[22][15:8] = buffer_data_1[1711:1704];
        layer3[22][23:16] = buffer_data_1[1719:1712];
        layer3[22][31:24] = buffer_data_1[1727:1720];
        layer3[22][39:32] = buffer_data_1[1735:1728];
        layer4[22][7:0] = buffer_data_0[1703:1696];
        layer4[22][15:8] = buffer_data_0[1711:1704];
        layer4[22][23:16] = buffer_data_0[1719:1712];
        layer4[22][31:24] = buffer_data_0[1727:1720];
        layer4[22][39:32] = buffer_data_0[1735:1728];
        layer0[23][7:0] = buffer_data_4[1711:1704];
        layer0[23][15:8] = buffer_data_4[1719:1712];
        layer0[23][23:16] = buffer_data_4[1727:1720];
        layer0[23][31:24] = buffer_data_4[1735:1728];
        layer0[23][39:32] = buffer_data_4[1743:1736];
        layer1[23][7:0] = buffer_data_3[1711:1704];
        layer1[23][15:8] = buffer_data_3[1719:1712];
        layer1[23][23:16] = buffer_data_3[1727:1720];
        layer1[23][31:24] = buffer_data_3[1735:1728];
        layer1[23][39:32] = buffer_data_3[1743:1736];
        layer2[23][7:0] = buffer_data_2[1711:1704];
        layer2[23][15:8] = buffer_data_2[1719:1712];
        layer2[23][23:16] = buffer_data_2[1727:1720];
        layer2[23][31:24] = buffer_data_2[1735:1728];
        layer2[23][39:32] = buffer_data_2[1743:1736];
        layer3[23][7:0] = buffer_data_1[1711:1704];
        layer3[23][15:8] = buffer_data_1[1719:1712];
        layer3[23][23:16] = buffer_data_1[1727:1720];
        layer3[23][31:24] = buffer_data_1[1735:1728];
        layer3[23][39:32] = buffer_data_1[1743:1736];
        layer4[23][7:0] = buffer_data_0[1711:1704];
        layer4[23][15:8] = buffer_data_0[1719:1712];
        layer4[23][23:16] = buffer_data_0[1727:1720];
        layer4[23][31:24] = buffer_data_0[1735:1728];
        layer4[23][39:32] = buffer_data_0[1743:1736];
        layer0[24][7:0] = buffer_data_4[1719:1712];
        layer0[24][15:8] = buffer_data_4[1727:1720];
        layer0[24][23:16] = buffer_data_4[1735:1728];
        layer0[24][31:24] = buffer_data_4[1743:1736];
        layer0[24][39:32] = buffer_data_4[1751:1744];
        layer1[24][7:0] = buffer_data_3[1719:1712];
        layer1[24][15:8] = buffer_data_3[1727:1720];
        layer1[24][23:16] = buffer_data_3[1735:1728];
        layer1[24][31:24] = buffer_data_3[1743:1736];
        layer1[24][39:32] = buffer_data_3[1751:1744];
        layer2[24][7:0] = buffer_data_2[1719:1712];
        layer2[24][15:8] = buffer_data_2[1727:1720];
        layer2[24][23:16] = buffer_data_2[1735:1728];
        layer2[24][31:24] = buffer_data_2[1743:1736];
        layer2[24][39:32] = buffer_data_2[1751:1744];
        layer3[24][7:0] = buffer_data_1[1719:1712];
        layer3[24][15:8] = buffer_data_1[1727:1720];
        layer3[24][23:16] = buffer_data_1[1735:1728];
        layer3[24][31:24] = buffer_data_1[1743:1736];
        layer3[24][39:32] = buffer_data_1[1751:1744];
        layer4[24][7:0] = buffer_data_0[1719:1712];
        layer4[24][15:8] = buffer_data_0[1727:1720];
        layer4[24][23:16] = buffer_data_0[1735:1728];
        layer4[24][31:24] = buffer_data_0[1743:1736];
        layer4[24][39:32] = buffer_data_0[1751:1744];
        layer0[25][7:0] = buffer_data_4[1727:1720];
        layer0[25][15:8] = buffer_data_4[1735:1728];
        layer0[25][23:16] = buffer_data_4[1743:1736];
        layer0[25][31:24] = buffer_data_4[1751:1744];
        layer0[25][39:32] = buffer_data_4[1759:1752];
        layer1[25][7:0] = buffer_data_3[1727:1720];
        layer1[25][15:8] = buffer_data_3[1735:1728];
        layer1[25][23:16] = buffer_data_3[1743:1736];
        layer1[25][31:24] = buffer_data_3[1751:1744];
        layer1[25][39:32] = buffer_data_3[1759:1752];
        layer2[25][7:0] = buffer_data_2[1727:1720];
        layer2[25][15:8] = buffer_data_2[1735:1728];
        layer2[25][23:16] = buffer_data_2[1743:1736];
        layer2[25][31:24] = buffer_data_2[1751:1744];
        layer2[25][39:32] = buffer_data_2[1759:1752];
        layer3[25][7:0] = buffer_data_1[1727:1720];
        layer3[25][15:8] = buffer_data_1[1735:1728];
        layer3[25][23:16] = buffer_data_1[1743:1736];
        layer3[25][31:24] = buffer_data_1[1751:1744];
        layer3[25][39:32] = buffer_data_1[1759:1752];
        layer4[25][7:0] = buffer_data_0[1727:1720];
        layer4[25][15:8] = buffer_data_0[1735:1728];
        layer4[25][23:16] = buffer_data_0[1743:1736];
        layer4[25][31:24] = buffer_data_0[1751:1744];
        layer4[25][39:32] = buffer_data_0[1759:1752];
        layer0[26][7:0] = buffer_data_4[1735:1728];
        layer0[26][15:8] = buffer_data_4[1743:1736];
        layer0[26][23:16] = buffer_data_4[1751:1744];
        layer0[26][31:24] = buffer_data_4[1759:1752];
        layer0[26][39:32] = buffer_data_4[1767:1760];
        layer1[26][7:0] = buffer_data_3[1735:1728];
        layer1[26][15:8] = buffer_data_3[1743:1736];
        layer1[26][23:16] = buffer_data_3[1751:1744];
        layer1[26][31:24] = buffer_data_3[1759:1752];
        layer1[26][39:32] = buffer_data_3[1767:1760];
        layer2[26][7:0] = buffer_data_2[1735:1728];
        layer2[26][15:8] = buffer_data_2[1743:1736];
        layer2[26][23:16] = buffer_data_2[1751:1744];
        layer2[26][31:24] = buffer_data_2[1759:1752];
        layer2[26][39:32] = buffer_data_2[1767:1760];
        layer3[26][7:0] = buffer_data_1[1735:1728];
        layer3[26][15:8] = buffer_data_1[1743:1736];
        layer3[26][23:16] = buffer_data_1[1751:1744];
        layer3[26][31:24] = buffer_data_1[1759:1752];
        layer3[26][39:32] = buffer_data_1[1767:1760];
        layer4[26][7:0] = buffer_data_0[1735:1728];
        layer4[26][15:8] = buffer_data_0[1743:1736];
        layer4[26][23:16] = buffer_data_0[1751:1744];
        layer4[26][31:24] = buffer_data_0[1759:1752];
        layer4[26][39:32] = buffer_data_0[1767:1760];
        layer0[27][7:0] = buffer_data_4[1743:1736];
        layer0[27][15:8] = buffer_data_4[1751:1744];
        layer0[27][23:16] = buffer_data_4[1759:1752];
        layer0[27][31:24] = buffer_data_4[1767:1760];
        layer0[27][39:32] = buffer_data_4[1775:1768];
        layer1[27][7:0] = buffer_data_3[1743:1736];
        layer1[27][15:8] = buffer_data_3[1751:1744];
        layer1[27][23:16] = buffer_data_3[1759:1752];
        layer1[27][31:24] = buffer_data_3[1767:1760];
        layer1[27][39:32] = buffer_data_3[1775:1768];
        layer2[27][7:0] = buffer_data_2[1743:1736];
        layer2[27][15:8] = buffer_data_2[1751:1744];
        layer2[27][23:16] = buffer_data_2[1759:1752];
        layer2[27][31:24] = buffer_data_2[1767:1760];
        layer2[27][39:32] = buffer_data_2[1775:1768];
        layer3[27][7:0] = buffer_data_1[1743:1736];
        layer3[27][15:8] = buffer_data_1[1751:1744];
        layer3[27][23:16] = buffer_data_1[1759:1752];
        layer3[27][31:24] = buffer_data_1[1767:1760];
        layer3[27][39:32] = buffer_data_1[1775:1768];
        layer4[27][7:0] = buffer_data_0[1743:1736];
        layer4[27][15:8] = buffer_data_0[1751:1744];
        layer4[27][23:16] = buffer_data_0[1759:1752];
        layer4[27][31:24] = buffer_data_0[1767:1760];
        layer4[27][39:32] = buffer_data_0[1775:1768];
        layer0[28][7:0] = buffer_data_4[1751:1744];
        layer0[28][15:8] = buffer_data_4[1759:1752];
        layer0[28][23:16] = buffer_data_4[1767:1760];
        layer0[28][31:24] = buffer_data_4[1775:1768];
        layer0[28][39:32] = buffer_data_4[1783:1776];
        layer1[28][7:0] = buffer_data_3[1751:1744];
        layer1[28][15:8] = buffer_data_3[1759:1752];
        layer1[28][23:16] = buffer_data_3[1767:1760];
        layer1[28][31:24] = buffer_data_3[1775:1768];
        layer1[28][39:32] = buffer_data_3[1783:1776];
        layer2[28][7:0] = buffer_data_2[1751:1744];
        layer2[28][15:8] = buffer_data_2[1759:1752];
        layer2[28][23:16] = buffer_data_2[1767:1760];
        layer2[28][31:24] = buffer_data_2[1775:1768];
        layer2[28][39:32] = buffer_data_2[1783:1776];
        layer3[28][7:0] = buffer_data_1[1751:1744];
        layer3[28][15:8] = buffer_data_1[1759:1752];
        layer3[28][23:16] = buffer_data_1[1767:1760];
        layer3[28][31:24] = buffer_data_1[1775:1768];
        layer3[28][39:32] = buffer_data_1[1783:1776];
        layer4[28][7:0] = buffer_data_0[1751:1744];
        layer4[28][15:8] = buffer_data_0[1759:1752];
        layer4[28][23:16] = buffer_data_0[1767:1760];
        layer4[28][31:24] = buffer_data_0[1775:1768];
        layer4[28][39:32] = buffer_data_0[1783:1776];
        layer0[29][7:0] = buffer_data_4[1759:1752];
        layer0[29][15:8] = buffer_data_4[1767:1760];
        layer0[29][23:16] = buffer_data_4[1775:1768];
        layer0[29][31:24] = buffer_data_4[1783:1776];
        layer0[29][39:32] = buffer_data_4[1791:1784];
        layer1[29][7:0] = buffer_data_3[1759:1752];
        layer1[29][15:8] = buffer_data_3[1767:1760];
        layer1[29][23:16] = buffer_data_3[1775:1768];
        layer1[29][31:24] = buffer_data_3[1783:1776];
        layer1[29][39:32] = buffer_data_3[1791:1784];
        layer2[29][7:0] = buffer_data_2[1759:1752];
        layer2[29][15:8] = buffer_data_2[1767:1760];
        layer2[29][23:16] = buffer_data_2[1775:1768];
        layer2[29][31:24] = buffer_data_2[1783:1776];
        layer2[29][39:32] = buffer_data_2[1791:1784];
        layer3[29][7:0] = buffer_data_1[1759:1752];
        layer3[29][15:8] = buffer_data_1[1767:1760];
        layer3[29][23:16] = buffer_data_1[1775:1768];
        layer3[29][31:24] = buffer_data_1[1783:1776];
        layer3[29][39:32] = buffer_data_1[1791:1784];
        layer4[29][7:0] = buffer_data_0[1759:1752];
        layer4[29][15:8] = buffer_data_0[1767:1760];
        layer4[29][23:16] = buffer_data_0[1775:1768];
        layer4[29][31:24] = buffer_data_0[1783:1776];
        layer4[29][39:32] = buffer_data_0[1791:1784];
        layer0[30][7:0] = buffer_data_4[1767:1760];
        layer0[30][15:8] = buffer_data_4[1775:1768];
        layer0[30][23:16] = buffer_data_4[1783:1776];
        layer0[30][31:24] = buffer_data_4[1791:1784];
        layer0[30][39:32] = buffer_data_4[1799:1792];
        layer1[30][7:0] = buffer_data_3[1767:1760];
        layer1[30][15:8] = buffer_data_3[1775:1768];
        layer1[30][23:16] = buffer_data_3[1783:1776];
        layer1[30][31:24] = buffer_data_3[1791:1784];
        layer1[30][39:32] = buffer_data_3[1799:1792];
        layer2[30][7:0] = buffer_data_2[1767:1760];
        layer2[30][15:8] = buffer_data_2[1775:1768];
        layer2[30][23:16] = buffer_data_2[1783:1776];
        layer2[30][31:24] = buffer_data_2[1791:1784];
        layer2[30][39:32] = buffer_data_2[1799:1792];
        layer3[30][7:0] = buffer_data_1[1767:1760];
        layer3[30][15:8] = buffer_data_1[1775:1768];
        layer3[30][23:16] = buffer_data_1[1783:1776];
        layer3[30][31:24] = buffer_data_1[1791:1784];
        layer3[30][39:32] = buffer_data_1[1799:1792];
        layer4[30][7:0] = buffer_data_0[1767:1760];
        layer4[30][15:8] = buffer_data_0[1775:1768];
        layer4[30][23:16] = buffer_data_0[1783:1776];
        layer4[30][31:24] = buffer_data_0[1791:1784];
        layer4[30][39:32] = buffer_data_0[1799:1792];
        layer0[31][7:0] = buffer_data_4[1775:1768];
        layer0[31][15:8] = buffer_data_4[1783:1776];
        layer0[31][23:16] = buffer_data_4[1791:1784];
        layer0[31][31:24] = buffer_data_4[1799:1792];
        layer0[31][39:32] = buffer_data_4[1807:1800];
        layer1[31][7:0] = buffer_data_3[1775:1768];
        layer1[31][15:8] = buffer_data_3[1783:1776];
        layer1[31][23:16] = buffer_data_3[1791:1784];
        layer1[31][31:24] = buffer_data_3[1799:1792];
        layer1[31][39:32] = buffer_data_3[1807:1800];
        layer2[31][7:0] = buffer_data_2[1775:1768];
        layer2[31][15:8] = buffer_data_2[1783:1776];
        layer2[31][23:16] = buffer_data_2[1791:1784];
        layer2[31][31:24] = buffer_data_2[1799:1792];
        layer2[31][39:32] = buffer_data_2[1807:1800];
        layer3[31][7:0] = buffer_data_1[1775:1768];
        layer3[31][15:8] = buffer_data_1[1783:1776];
        layer3[31][23:16] = buffer_data_1[1791:1784];
        layer3[31][31:24] = buffer_data_1[1799:1792];
        layer3[31][39:32] = buffer_data_1[1807:1800];
        layer4[31][7:0] = buffer_data_0[1775:1768];
        layer4[31][15:8] = buffer_data_0[1783:1776];
        layer4[31][23:16] = buffer_data_0[1791:1784];
        layer4[31][31:24] = buffer_data_0[1799:1792];
        layer4[31][39:32] = buffer_data_0[1807:1800];
        layer0[32][7:0] = buffer_data_4[1783:1776];
        layer0[32][15:8] = buffer_data_4[1791:1784];
        layer0[32][23:16] = buffer_data_4[1799:1792];
        layer0[32][31:24] = buffer_data_4[1807:1800];
        layer0[32][39:32] = buffer_data_4[1815:1808];
        layer1[32][7:0] = buffer_data_3[1783:1776];
        layer1[32][15:8] = buffer_data_3[1791:1784];
        layer1[32][23:16] = buffer_data_3[1799:1792];
        layer1[32][31:24] = buffer_data_3[1807:1800];
        layer1[32][39:32] = buffer_data_3[1815:1808];
        layer2[32][7:0] = buffer_data_2[1783:1776];
        layer2[32][15:8] = buffer_data_2[1791:1784];
        layer2[32][23:16] = buffer_data_2[1799:1792];
        layer2[32][31:24] = buffer_data_2[1807:1800];
        layer2[32][39:32] = buffer_data_2[1815:1808];
        layer3[32][7:0] = buffer_data_1[1783:1776];
        layer3[32][15:8] = buffer_data_1[1791:1784];
        layer3[32][23:16] = buffer_data_1[1799:1792];
        layer3[32][31:24] = buffer_data_1[1807:1800];
        layer3[32][39:32] = buffer_data_1[1815:1808];
        layer4[32][7:0] = buffer_data_0[1783:1776];
        layer4[32][15:8] = buffer_data_0[1791:1784];
        layer4[32][23:16] = buffer_data_0[1799:1792];
        layer4[32][31:24] = buffer_data_0[1807:1800];
        layer4[32][39:32] = buffer_data_0[1815:1808];
        layer0[33][7:0] = buffer_data_4[1791:1784];
        layer0[33][15:8] = buffer_data_4[1799:1792];
        layer0[33][23:16] = buffer_data_4[1807:1800];
        layer0[33][31:24] = buffer_data_4[1815:1808];
        layer0[33][39:32] = buffer_data_4[1823:1816];
        layer1[33][7:0] = buffer_data_3[1791:1784];
        layer1[33][15:8] = buffer_data_3[1799:1792];
        layer1[33][23:16] = buffer_data_3[1807:1800];
        layer1[33][31:24] = buffer_data_3[1815:1808];
        layer1[33][39:32] = buffer_data_3[1823:1816];
        layer2[33][7:0] = buffer_data_2[1791:1784];
        layer2[33][15:8] = buffer_data_2[1799:1792];
        layer2[33][23:16] = buffer_data_2[1807:1800];
        layer2[33][31:24] = buffer_data_2[1815:1808];
        layer2[33][39:32] = buffer_data_2[1823:1816];
        layer3[33][7:0] = buffer_data_1[1791:1784];
        layer3[33][15:8] = buffer_data_1[1799:1792];
        layer3[33][23:16] = buffer_data_1[1807:1800];
        layer3[33][31:24] = buffer_data_1[1815:1808];
        layer3[33][39:32] = buffer_data_1[1823:1816];
        layer4[33][7:0] = buffer_data_0[1791:1784];
        layer4[33][15:8] = buffer_data_0[1799:1792];
        layer4[33][23:16] = buffer_data_0[1807:1800];
        layer4[33][31:24] = buffer_data_0[1815:1808];
        layer4[33][39:32] = buffer_data_0[1823:1816];
        layer0[34][7:0] = buffer_data_4[1799:1792];
        layer0[34][15:8] = buffer_data_4[1807:1800];
        layer0[34][23:16] = buffer_data_4[1815:1808];
        layer0[34][31:24] = buffer_data_4[1823:1816];
        layer0[34][39:32] = buffer_data_4[1831:1824];
        layer1[34][7:0] = buffer_data_3[1799:1792];
        layer1[34][15:8] = buffer_data_3[1807:1800];
        layer1[34][23:16] = buffer_data_3[1815:1808];
        layer1[34][31:24] = buffer_data_3[1823:1816];
        layer1[34][39:32] = buffer_data_3[1831:1824];
        layer2[34][7:0] = buffer_data_2[1799:1792];
        layer2[34][15:8] = buffer_data_2[1807:1800];
        layer2[34][23:16] = buffer_data_2[1815:1808];
        layer2[34][31:24] = buffer_data_2[1823:1816];
        layer2[34][39:32] = buffer_data_2[1831:1824];
        layer3[34][7:0] = buffer_data_1[1799:1792];
        layer3[34][15:8] = buffer_data_1[1807:1800];
        layer3[34][23:16] = buffer_data_1[1815:1808];
        layer3[34][31:24] = buffer_data_1[1823:1816];
        layer3[34][39:32] = buffer_data_1[1831:1824];
        layer4[34][7:0] = buffer_data_0[1799:1792];
        layer4[34][15:8] = buffer_data_0[1807:1800];
        layer4[34][23:16] = buffer_data_0[1815:1808];
        layer4[34][31:24] = buffer_data_0[1823:1816];
        layer4[34][39:32] = buffer_data_0[1831:1824];
        layer0[35][7:0] = buffer_data_4[1807:1800];
        layer0[35][15:8] = buffer_data_4[1815:1808];
        layer0[35][23:16] = buffer_data_4[1823:1816];
        layer0[35][31:24] = buffer_data_4[1831:1824];
        layer0[35][39:32] = buffer_data_4[1839:1832];
        layer1[35][7:0] = buffer_data_3[1807:1800];
        layer1[35][15:8] = buffer_data_3[1815:1808];
        layer1[35][23:16] = buffer_data_3[1823:1816];
        layer1[35][31:24] = buffer_data_3[1831:1824];
        layer1[35][39:32] = buffer_data_3[1839:1832];
        layer2[35][7:0] = buffer_data_2[1807:1800];
        layer2[35][15:8] = buffer_data_2[1815:1808];
        layer2[35][23:16] = buffer_data_2[1823:1816];
        layer2[35][31:24] = buffer_data_2[1831:1824];
        layer2[35][39:32] = buffer_data_2[1839:1832];
        layer3[35][7:0] = buffer_data_1[1807:1800];
        layer3[35][15:8] = buffer_data_1[1815:1808];
        layer3[35][23:16] = buffer_data_1[1823:1816];
        layer3[35][31:24] = buffer_data_1[1831:1824];
        layer3[35][39:32] = buffer_data_1[1839:1832];
        layer4[35][7:0] = buffer_data_0[1807:1800];
        layer4[35][15:8] = buffer_data_0[1815:1808];
        layer4[35][23:16] = buffer_data_0[1823:1816];
        layer4[35][31:24] = buffer_data_0[1831:1824];
        layer4[35][39:32] = buffer_data_0[1839:1832];
        layer0[36][7:0] = buffer_data_4[1815:1808];
        layer0[36][15:8] = buffer_data_4[1823:1816];
        layer0[36][23:16] = buffer_data_4[1831:1824];
        layer0[36][31:24] = buffer_data_4[1839:1832];
        layer0[36][39:32] = buffer_data_4[1847:1840];
        layer1[36][7:0] = buffer_data_3[1815:1808];
        layer1[36][15:8] = buffer_data_3[1823:1816];
        layer1[36][23:16] = buffer_data_3[1831:1824];
        layer1[36][31:24] = buffer_data_3[1839:1832];
        layer1[36][39:32] = buffer_data_3[1847:1840];
        layer2[36][7:0] = buffer_data_2[1815:1808];
        layer2[36][15:8] = buffer_data_2[1823:1816];
        layer2[36][23:16] = buffer_data_2[1831:1824];
        layer2[36][31:24] = buffer_data_2[1839:1832];
        layer2[36][39:32] = buffer_data_2[1847:1840];
        layer3[36][7:0] = buffer_data_1[1815:1808];
        layer3[36][15:8] = buffer_data_1[1823:1816];
        layer3[36][23:16] = buffer_data_1[1831:1824];
        layer3[36][31:24] = buffer_data_1[1839:1832];
        layer3[36][39:32] = buffer_data_1[1847:1840];
        layer4[36][7:0] = buffer_data_0[1815:1808];
        layer4[36][15:8] = buffer_data_0[1823:1816];
        layer4[36][23:16] = buffer_data_0[1831:1824];
        layer4[36][31:24] = buffer_data_0[1839:1832];
        layer4[36][39:32] = buffer_data_0[1847:1840];
        layer0[37][7:0] = buffer_data_4[1823:1816];
        layer0[37][15:8] = buffer_data_4[1831:1824];
        layer0[37][23:16] = buffer_data_4[1839:1832];
        layer0[37][31:24] = buffer_data_4[1847:1840];
        layer0[37][39:32] = buffer_data_4[1855:1848];
        layer1[37][7:0] = buffer_data_3[1823:1816];
        layer1[37][15:8] = buffer_data_3[1831:1824];
        layer1[37][23:16] = buffer_data_3[1839:1832];
        layer1[37][31:24] = buffer_data_3[1847:1840];
        layer1[37][39:32] = buffer_data_3[1855:1848];
        layer2[37][7:0] = buffer_data_2[1823:1816];
        layer2[37][15:8] = buffer_data_2[1831:1824];
        layer2[37][23:16] = buffer_data_2[1839:1832];
        layer2[37][31:24] = buffer_data_2[1847:1840];
        layer2[37][39:32] = buffer_data_2[1855:1848];
        layer3[37][7:0] = buffer_data_1[1823:1816];
        layer3[37][15:8] = buffer_data_1[1831:1824];
        layer3[37][23:16] = buffer_data_1[1839:1832];
        layer3[37][31:24] = buffer_data_1[1847:1840];
        layer3[37][39:32] = buffer_data_1[1855:1848];
        layer4[37][7:0] = buffer_data_0[1823:1816];
        layer4[37][15:8] = buffer_data_0[1831:1824];
        layer4[37][23:16] = buffer_data_0[1839:1832];
        layer4[37][31:24] = buffer_data_0[1847:1840];
        layer4[37][39:32] = buffer_data_0[1855:1848];
        layer0[38][7:0] = buffer_data_4[1831:1824];
        layer0[38][15:8] = buffer_data_4[1839:1832];
        layer0[38][23:16] = buffer_data_4[1847:1840];
        layer0[38][31:24] = buffer_data_4[1855:1848];
        layer0[38][39:32] = buffer_data_4[1863:1856];
        layer1[38][7:0] = buffer_data_3[1831:1824];
        layer1[38][15:8] = buffer_data_3[1839:1832];
        layer1[38][23:16] = buffer_data_3[1847:1840];
        layer1[38][31:24] = buffer_data_3[1855:1848];
        layer1[38][39:32] = buffer_data_3[1863:1856];
        layer2[38][7:0] = buffer_data_2[1831:1824];
        layer2[38][15:8] = buffer_data_2[1839:1832];
        layer2[38][23:16] = buffer_data_2[1847:1840];
        layer2[38][31:24] = buffer_data_2[1855:1848];
        layer2[38][39:32] = buffer_data_2[1863:1856];
        layer3[38][7:0] = buffer_data_1[1831:1824];
        layer3[38][15:8] = buffer_data_1[1839:1832];
        layer3[38][23:16] = buffer_data_1[1847:1840];
        layer3[38][31:24] = buffer_data_1[1855:1848];
        layer3[38][39:32] = buffer_data_1[1863:1856];
        layer4[38][7:0] = buffer_data_0[1831:1824];
        layer4[38][15:8] = buffer_data_0[1839:1832];
        layer4[38][23:16] = buffer_data_0[1847:1840];
        layer4[38][31:24] = buffer_data_0[1855:1848];
        layer4[38][39:32] = buffer_data_0[1863:1856];
        layer0[39][7:0] = buffer_data_4[1839:1832];
        layer0[39][15:8] = buffer_data_4[1847:1840];
        layer0[39][23:16] = buffer_data_4[1855:1848];
        layer0[39][31:24] = buffer_data_4[1863:1856];
        layer0[39][39:32] = buffer_data_4[1871:1864];
        layer1[39][7:0] = buffer_data_3[1839:1832];
        layer1[39][15:8] = buffer_data_3[1847:1840];
        layer1[39][23:16] = buffer_data_3[1855:1848];
        layer1[39][31:24] = buffer_data_3[1863:1856];
        layer1[39][39:32] = buffer_data_3[1871:1864];
        layer2[39][7:0] = buffer_data_2[1839:1832];
        layer2[39][15:8] = buffer_data_2[1847:1840];
        layer2[39][23:16] = buffer_data_2[1855:1848];
        layer2[39][31:24] = buffer_data_2[1863:1856];
        layer2[39][39:32] = buffer_data_2[1871:1864];
        layer3[39][7:0] = buffer_data_1[1839:1832];
        layer3[39][15:8] = buffer_data_1[1847:1840];
        layer3[39][23:16] = buffer_data_1[1855:1848];
        layer3[39][31:24] = buffer_data_1[1863:1856];
        layer3[39][39:32] = buffer_data_1[1871:1864];
        layer4[39][7:0] = buffer_data_0[1839:1832];
        layer4[39][15:8] = buffer_data_0[1847:1840];
        layer4[39][23:16] = buffer_data_0[1855:1848];
        layer4[39][31:24] = buffer_data_0[1863:1856];
        layer4[39][39:32] = buffer_data_0[1871:1864];
        layer0[40][7:0] = buffer_data_4[1847:1840];
        layer0[40][15:8] = buffer_data_4[1855:1848];
        layer0[40][23:16] = buffer_data_4[1863:1856];
        layer0[40][31:24] = buffer_data_4[1871:1864];
        layer0[40][39:32] = buffer_data_4[1879:1872];
        layer1[40][7:0] = buffer_data_3[1847:1840];
        layer1[40][15:8] = buffer_data_3[1855:1848];
        layer1[40][23:16] = buffer_data_3[1863:1856];
        layer1[40][31:24] = buffer_data_3[1871:1864];
        layer1[40][39:32] = buffer_data_3[1879:1872];
        layer2[40][7:0] = buffer_data_2[1847:1840];
        layer2[40][15:8] = buffer_data_2[1855:1848];
        layer2[40][23:16] = buffer_data_2[1863:1856];
        layer2[40][31:24] = buffer_data_2[1871:1864];
        layer2[40][39:32] = buffer_data_2[1879:1872];
        layer3[40][7:0] = buffer_data_1[1847:1840];
        layer3[40][15:8] = buffer_data_1[1855:1848];
        layer3[40][23:16] = buffer_data_1[1863:1856];
        layer3[40][31:24] = buffer_data_1[1871:1864];
        layer3[40][39:32] = buffer_data_1[1879:1872];
        layer4[40][7:0] = buffer_data_0[1847:1840];
        layer4[40][15:8] = buffer_data_0[1855:1848];
        layer4[40][23:16] = buffer_data_0[1863:1856];
        layer4[40][31:24] = buffer_data_0[1871:1864];
        layer4[40][39:32] = buffer_data_0[1879:1872];
        layer0[41][7:0] = buffer_data_4[1855:1848];
        layer0[41][15:8] = buffer_data_4[1863:1856];
        layer0[41][23:16] = buffer_data_4[1871:1864];
        layer0[41][31:24] = buffer_data_4[1879:1872];
        layer0[41][39:32] = buffer_data_4[1887:1880];
        layer1[41][7:0] = buffer_data_3[1855:1848];
        layer1[41][15:8] = buffer_data_3[1863:1856];
        layer1[41][23:16] = buffer_data_3[1871:1864];
        layer1[41][31:24] = buffer_data_3[1879:1872];
        layer1[41][39:32] = buffer_data_3[1887:1880];
        layer2[41][7:0] = buffer_data_2[1855:1848];
        layer2[41][15:8] = buffer_data_2[1863:1856];
        layer2[41][23:16] = buffer_data_2[1871:1864];
        layer2[41][31:24] = buffer_data_2[1879:1872];
        layer2[41][39:32] = buffer_data_2[1887:1880];
        layer3[41][7:0] = buffer_data_1[1855:1848];
        layer3[41][15:8] = buffer_data_1[1863:1856];
        layer3[41][23:16] = buffer_data_1[1871:1864];
        layer3[41][31:24] = buffer_data_1[1879:1872];
        layer3[41][39:32] = buffer_data_1[1887:1880];
        layer4[41][7:0] = buffer_data_0[1855:1848];
        layer4[41][15:8] = buffer_data_0[1863:1856];
        layer4[41][23:16] = buffer_data_0[1871:1864];
        layer4[41][31:24] = buffer_data_0[1879:1872];
        layer4[41][39:32] = buffer_data_0[1887:1880];
        layer0[42][7:0] = buffer_data_4[1863:1856];
        layer0[42][15:8] = buffer_data_4[1871:1864];
        layer0[42][23:16] = buffer_data_4[1879:1872];
        layer0[42][31:24] = buffer_data_4[1887:1880];
        layer0[42][39:32] = buffer_data_4[1895:1888];
        layer1[42][7:0] = buffer_data_3[1863:1856];
        layer1[42][15:8] = buffer_data_3[1871:1864];
        layer1[42][23:16] = buffer_data_3[1879:1872];
        layer1[42][31:24] = buffer_data_3[1887:1880];
        layer1[42][39:32] = buffer_data_3[1895:1888];
        layer2[42][7:0] = buffer_data_2[1863:1856];
        layer2[42][15:8] = buffer_data_2[1871:1864];
        layer2[42][23:16] = buffer_data_2[1879:1872];
        layer2[42][31:24] = buffer_data_2[1887:1880];
        layer2[42][39:32] = buffer_data_2[1895:1888];
        layer3[42][7:0] = buffer_data_1[1863:1856];
        layer3[42][15:8] = buffer_data_1[1871:1864];
        layer3[42][23:16] = buffer_data_1[1879:1872];
        layer3[42][31:24] = buffer_data_1[1887:1880];
        layer3[42][39:32] = buffer_data_1[1895:1888];
        layer4[42][7:0] = buffer_data_0[1863:1856];
        layer4[42][15:8] = buffer_data_0[1871:1864];
        layer4[42][23:16] = buffer_data_0[1879:1872];
        layer4[42][31:24] = buffer_data_0[1887:1880];
        layer4[42][39:32] = buffer_data_0[1895:1888];
        layer0[43][7:0] = buffer_data_4[1871:1864];
        layer0[43][15:8] = buffer_data_4[1879:1872];
        layer0[43][23:16] = buffer_data_4[1887:1880];
        layer0[43][31:24] = buffer_data_4[1895:1888];
        layer0[43][39:32] = buffer_data_4[1903:1896];
        layer1[43][7:0] = buffer_data_3[1871:1864];
        layer1[43][15:8] = buffer_data_3[1879:1872];
        layer1[43][23:16] = buffer_data_3[1887:1880];
        layer1[43][31:24] = buffer_data_3[1895:1888];
        layer1[43][39:32] = buffer_data_3[1903:1896];
        layer2[43][7:0] = buffer_data_2[1871:1864];
        layer2[43][15:8] = buffer_data_2[1879:1872];
        layer2[43][23:16] = buffer_data_2[1887:1880];
        layer2[43][31:24] = buffer_data_2[1895:1888];
        layer2[43][39:32] = buffer_data_2[1903:1896];
        layer3[43][7:0] = buffer_data_1[1871:1864];
        layer3[43][15:8] = buffer_data_1[1879:1872];
        layer3[43][23:16] = buffer_data_1[1887:1880];
        layer3[43][31:24] = buffer_data_1[1895:1888];
        layer3[43][39:32] = buffer_data_1[1903:1896];
        layer4[43][7:0] = buffer_data_0[1871:1864];
        layer4[43][15:8] = buffer_data_0[1879:1872];
        layer4[43][23:16] = buffer_data_0[1887:1880];
        layer4[43][31:24] = buffer_data_0[1895:1888];
        layer4[43][39:32] = buffer_data_0[1903:1896];
        layer0[44][7:0] = buffer_data_4[1879:1872];
        layer0[44][15:8] = buffer_data_4[1887:1880];
        layer0[44][23:16] = buffer_data_4[1895:1888];
        layer0[44][31:24] = buffer_data_4[1903:1896];
        layer0[44][39:32] = buffer_data_4[1911:1904];
        layer1[44][7:0] = buffer_data_3[1879:1872];
        layer1[44][15:8] = buffer_data_3[1887:1880];
        layer1[44][23:16] = buffer_data_3[1895:1888];
        layer1[44][31:24] = buffer_data_3[1903:1896];
        layer1[44][39:32] = buffer_data_3[1911:1904];
        layer2[44][7:0] = buffer_data_2[1879:1872];
        layer2[44][15:8] = buffer_data_2[1887:1880];
        layer2[44][23:16] = buffer_data_2[1895:1888];
        layer2[44][31:24] = buffer_data_2[1903:1896];
        layer2[44][39:32] = buffer_data_2[1911:1904];
        layer3[44][7:0] = buffer_data_1[1879:1872];
        layer3[44][15:8] = buffer_data_1[1887:1880];
        layer3[44][23:16] = buffer_data_1[1895:1888];
        layer3[44][31:24] = buffer_data_1[1903:1896];
        layer3[44][39:32] = buffer_data_1[1911:1904];
        layer4[44][7:0] = buffer_data_0[1879:1872];
        layer4[44][15:8] = buffer_data_0[1887:1880];
        layer4[44][23:16] = buffer_data_0[1895:1888];
        layer4[44][31:24] = buffer_data_0[1903:1896];
        layer4[44][39:32] = buffer_data_0[1911:1904];
        layer0[45][7:0] = buffer_data_4[1887:1880];
        layer0[45][15:8] = buffer_data_4[1895:1888];
        layer0[45][23:16] = buffer_data_4[1903:1896];
        layer0[45][31:24] = buffer_data_4[1911:1904];
        layer0[45][39:32] = buffer_data_4[1919:1912];
        layer1[45][7:0] = buffer_data_3[1887:1880];
        layer1[45][15:8] = buffer_data_3[1895:1888];
        layer1[45][23:16] = buffer_data_3[1903:1896];
        layer1[45][31:24] = buffer_data_3[1911:1904];
        layer1[45][39:32] = buffer_data_3[1919:1912];
        layer2[45][7:0] = buffer_data_2[1887:1880];
        layer2[45][15:8] = buffer_data_2[1895:1888];
        layer2[45][23:16] = buffer_data_2[1903:1896];
        layer2[45][31:24] = buffer_data_2[1911:1904];
        layer2[45][39:32] = buffer_data_2[1919:1912];
        layer3[45][7:0] = buffer_data_1[1887:1880];
        layer3[45][15:8] = buffer_data_1[1895:1888];
        layer3[45][23:16] = buffer_data_1[1903:1896];
        layer3[45][31:24] = buffer_data_1[1911:1904];
        layer3[45][39:32] = buffer_data_1[1919:1912];
        layer4[45][7:0] = buffer_data_0[1887:1880];
        layer4[45][15:8] = buffer_data_0[1895:1888];
        layer4[45][23:16] = buffer_data_0[1903:1896];
        layer4[45][31:24] = buffer_data_0[1911:1904];
        layer4[45][39:32] = buffer_data_0[1919:1912];
        layer0[46][7:0] = buffer_data_4[1895:1888];
        layer0[46][15:8] = buffer_data_4[1903:1896];
        layer0[46][23:16] = buffer_data_4[1911:1904];
        layer0[46][31:24] = buffer_data_4[1919:1912];
        layer0[46][39:32] = buffer_data_4[1927:1920];
        layer1[46][7:0] = buffer_data_3[1895:1888];
        layer1[46][15:8] = buffer_data_3[1903:1896];
        layer1[46][23:16] = buffer_data_3[1911:1904];
        layer1[46][31:24] = buffer_data_3[1919:1912];
        layer1[46][39:32] = buffer_data_3[1927:1920];
        layer2[46][7:0] = buffer_data_2[1895:1888];
        layer2[46][15:8] = buffer_data_2[1903:1896];
        layer2[46][23:16] = buffer_data_2[1911:1904];
        layer2[46][31:24] = buffer_data_2[1919:1912];
        layer2[46][39:32] = buffer_data_2[1927:1920];
        layer3[46][7:0] = buffer_data_1[1895:1888];
        layer3[46][15:8] = buffer_data_1[1903:1896];
        layer3[46][23:16] = buffer_data_1[1911:1904];
        layer3[46][31:24] = buffer_data_1[1919:1912];
        layer3[46][39:32] = buffer_data_1[1927:1920];
        layer4[46][7:0] = buffer_data_0[1895:1888];
        layer4[46][15:8] = buffer_data_0[1903:1896];
        layer4[46][23:16] = buffer_data_0[1911:1904];
        layer4[46][31:24] = buffer_data_0[1919:1912];
        layer4[46][39:32] = buffer_data_0[1927:1920];
        layer0[47][7:0] = buffer_data_4[1903:1896];
        layer0[47][15:8] = buffer_data_4[1911:1904];
        layer0[47][23:16] = buffer_data_4[1919:1912];
        layer0[47][31:24] = buffer_data_4[1927:1920];
        layer0[47][39:32] = buffer_data_4[1935:1928];
        layer1[47][7:0] = buffer_data_3[1903:1896];
        layer1[47][15:8] = buffer_data_3[1911:1904];
        layer1[47][23:16] = buffer_data_3[1919:1912];
        layer1[47][31:24] = buffer_data_3[1927:1920];
        layer1[47][39:32] = buffer_data_3[1935:1928];
        layer2[47][7:0] = buffer_data_2[1903:1896];
        layer2[47][15:8] = buffer_data_2[1911:1904];
        layer2[47][23:16] = buffer_data_2[1919:1912];
        layer2[47][31:24] = buffer_data_2[1927:1920];
        layer2[47][39:32] = buffer_data_2[1935:1928];
        layer3[47][7:0] = buffer_data_1[1903:1896];
        layer3[47][15:8] = buffer_data_1[1911:1904];
        layer3[47][23:16] = buffer_data_1[1919:1912];
        layer3[47][31:24] = buffer_data_1[1927:1920];
        layer3[47][39:32] = buffer_data_1[1935:1928];
        layer4[47][7:0] = buffer_data_0[1903:1896];
        layer4[47][15:8] = buffer_data_0[1911:1904];
        layer4[47][23:16] = buffer_data_0[1919:1912];
        layer4[47][31:24] = buffer_data_0[1927:1920];
        layer4[47][39:32] = buffer_data_0[1935:1928];
        layer0[48][7:0] = buffer_data_4[1911:1904];
        layer0[48][15:8] = buffer_data_4[1919:1912];
        layer0[48][23:16] = buffer_data_4[1927:1920];
        layer0[48][31:24] = buffer_data_4[1935:1928];
        layer0[48][39:32] = buffer_data_4[1943:1936];
        layer1[48][7:0] = buffer_data_3[1911:1904];
        layer1[48][15:8] = buffer_data_3[1919:1912];
        layer1[48][23:16] = buffer_data_3[1927:1920];
        layer1[48][31:24] = buffer_data_3[1935:1928];
        layer1[48][39:32] = buffer_data_3[1943:1936];
        layer2[48][7:0] = buffer_data_2[1911:1904];
        layer2[48][15:8] = buffer_data_2[1919:1912];
        layer2[48][23:16] = buffer_data_2[1927:1920];
        layer2[48][31:24] = buffer_data_2[1935:1928];
        layer2[48][39:32] = buffer_data_2[1943:1936];
        layer3[48][7:0] = buffer_data_1[1911:1904];
        layer3[48][15:8] = buffer_data_1[1919:1912];
        layer3[48][23:16] = buffer_data_1[1927:1920];
        layer3[48][31:24] = buffer_data_1[1935:1928];
        layer3[48][39:32] = buffer_data_1[1943:1936];
        layer4[48][7:0] = buffer_data_0[1911:1904];
        layer4[48][15:8] = buffer_data_0[1919:1912];
        layer4[48][23:16] = buffer_data_0[1927:1920];
        layer4[48][31:24] = buffer_data_0[1935:1928];
        layer4[48][39:32] = buffer_data_0[1943:1936];
        layer0[49][7:0] = buffer_data_4[1919:1912];
        layer0[49][15:8] = buffer_data_4[1927:1920];
        layer0[49][23:16] = buffer_data_4[1935:1928];
        layer0[49][31:24] = buffer_data_4[1943:1936];
        layer0[49][39:32] = buffer_data_4[1951:1944];
        layer1[49][7:0] = buffer_data_3[1919:1912];
        layer1[49][15:8] = buffer_data_3[1927:1920];
        layer1[49][23:16] = buffer_data_3[1935:1928];
        layer1[49][31:24] = buffer_data_3[1943:1936];
        layer1[49][39:32] = buffer_data_3[1951:1944];
        layer2[49][7:0] = buffer_data_2[1919:1912];
        layer2[49][15:8] = buffer_data_2[1927:1920];
        layer2[49][23:16] = buffer_data_2[1935:1928];
        layer2[49][31:24] = buffer_data_2[1943:1936];
        layer2[49][39:32] = buffer_data_2[1951:1944];
        layer3[49][7:0] = buffer_data_1[1919:1912];
        layer3[49][15:8] = buffer_data_1[1927:1920];
        layer3[49][23:16] = buffer_data_1[1935:1928];
        layer3[49][31:24] = buffer_data_1[1943:1936];
        layer3[49][39:32] = buffer_data_1[1951:1944];
        layer4[49][7:0] = buffer_data_0[1919:1912];
        layer4[49][15:8] = buffer_data_0[1927:1920];
        layer4[49][23:16] = buffer_data_0[1935:1928];
        layer4[49][31:24] = buffer_data_0[1943:1936];
        layer4[49][39:32] = buffer_data_0[1951:1944];
        layer0[50][7:0] = buffer_data_4[1927:1920];
        layer0[50][15:8] = buffer_data_4[1935:1928];
        layer0[50][23:16] = buffer_data_4[1943:1936];
        layer0[50][31:24] = buffer_data_4[1951:1944];
        layer0[50][39:32] = buffer_data_4[1959:1952];
        layer1[50][7:0] = buffer_data_3[1927:1920];
        layer1[50][15:8] = buffer_data_3[1935:1928];
        layer1[50][23:16] = buffer_data_3[1943:1936];
        layer1[50][31:24] = buffer_data_3[1951:1944];
        layer1[50][39:32] = buffer_data_3[1959:1952];
        layer2[50][7:0] = buffer_data_2[1927:1920];
        layer2[50][15:8] = buffer_data_2[1935:1928];
        layer2[50][23:16] = buffer_data_2[1943:1936];
        layer2[50][31:24] = buffer_data_2[1951:1944];
        layer2[50][39:32] = buffer_data_2[1959:1952];
        layer3[50][7:0] = buffer_data_1[1927:1920];
        layer3[50][15:8] = buffer_data_1[1935:1928];
        layer3[50][23:16] = buffer_data_1[1943:1936];
        layer3[50][31:24] = buffer_data_1[1951:1944];
        layer3[50][39:32] = buffer_data_1[1959:1952];
        layer4[50][7:0] = buffer_data_0[1927:1920];
        layer4[50][15:8] = buffer_data_0[1935:1928];
        layer4[50][23:16] = buffer_data_0[1943:1936];
        layer4[50][31:24] = buffer_data_0[1951:1944];
        layer4[50][39:32] = buffer_data_0[1959:1952];
        layer0[51][7:0] = buffer_data_4[1935:1928];
        layer0[51][15:8] = buffer_data_4[1943:1936];
        layer0[51][23:16] = buffer_data_4[1951:1944];
        layer0[51][31:24] = buffer_data_4[1959:1952];
        layer0[51][39:32] = buffer_data_4[1967:1960];
        layer1[51][7:0] = buffer_data_3[1935:1928];
        layer1[51][15:8] = buffer_data_3[1943:1936];
        layer1[51][23:16] = buffer_data_3[1951:1944];
        layer1[51][31:24] = buffer_data_3[1959:1952];
        layer1[51][39:32] = buffer_data_3[1967:1960];
        layer2[51][7:0] = buffer_data_2[1935:1928];
        layer2[51][15:8] = buffer_data_2[1943:1936];
        layer2[51][23:16] = buffer_data_2[1951:1944];
        layer2[51][31:24] = buffer_data_2[1959:1952];
        layer2[51][39:32] = buffer_data_2[1967:1960];
        layer3[51][7:0] = buffer_data_1[1935:1928];
        layer3[51][15:8] = buffer_data_1[1943:1936];
        layer3[51][23:16] = buffer_data_1[1951:1944];
        layer3[51][31:24] = buffer_data_1[1959:1952];
        layer3[51][39:32] = buffer_data_1[1967:1960];
        layer4[51][7:0] = buffer_data_0[1935:1928];
        layer4[51][15:8] = buffer_data_0[1943:1936];
        layer4[51][23:16] = buffer_data_0[1951:1944];
        layer4[51][31:24] = buffer_data_0[1959:1952];
        layer4[51][39:32] = buffer_data_0[1967:1960];
        layer0[52][7:0] = buffer_data_4[1943:1936];
        layer0[52][15:8] = buffer_data_4[1951:1944];
        layer0[52][23:16] = buffer_data_4[1959:1952];
        layer0[52][31:24] = buffer_data_4[1967:1960];
        layer0[52][39:32] = buffer_data_4[1975:1968];
        layer1[52][7:0] = buffer_data_3[1943:1936];
        layer1[52][15:8] = buffer_data_3[1951:1944];
        layer1[52][23:16] = buffer_data_3[1959:1952];
        layer1[52][31:24] = buffer_data_3[1967:1960];
        layer1[52][39:32] = buffer_data_3[1975:1968];
        layer2[52][7:0] = buffer_data_2[1943:1936];
        layer2[52][15:8] = buffer_data_2[1951:1944];
        layer2[52][23:16] = buffer_data_2[1959:1952];
        layer2[52][31:24] = buffer_data_2[1967:1960];
        layer2[52][39:32] = buffer_data_2[1975:1968];
        layer3[52][7:0] = buffer_data_1[1943:1936];
        layer3[52][15:8] = buffer_data_1[1951:1944];
        layer3[52][23:16] = buffer_data_1[1959:1952];
        layer3[52][31:24] = buffer_data_1[1967:1960];
        layer3[52][39:32] = buffer_data_1[1975:1968];
        layer4[52][7:0] = buffer_data_0[1943:1936];
        layer4[52][15:8] = buffer_data_0[1951:1944];
        layer4[52][23:16] = buffer_data_0[1959:1952];
        layer4[52][31:24] = buffer_data_0[1967:1960];
        layer4[52][39:32] = buffer_data_0[1975:1968];
        layer0[53][7:0] = buffer_data_4[1951:1944];
        layer0[53][15:8] = buffer_data_4[1959:1952];
        layer0[53][23:16] = buffer_data_4[1967:1960];
        layer0[53][31:24] = buffer_data_4[1975:1968];
        layer0[53][39:32] = buffer_data_4[1983:1976];
        layer1[53][7:0] = buffer_data_3[1951:1944];
        layer1[53][15:8] = buffer_data_3[1959:1952];
        layer1[53][23:16] = buffer_data_3[1967:1960];
        layer1[53][31:24] = buffer_data_3[1975:1968];
        layer1[53][39:32] = buffer_data_3[1983:1976];
        layer2[53][7:0] = buffer_data_2[1951:1944];
        layer2[53][15:8] = buffer_data_2[1959:1952];
        layer2[53][23:16] = buffer_data_2[1967:1960];
        layer2[53][31:24] = buffer_data_2[1975:1968];
        layer2[53][39:32] = buffer_data_2[1983:1976];
        layer3[53][7:0] = buffer_data_1[1951:1944];
        layer3[53][15:8] = buffer_data_1[1959:1952];
        layer3[53][23:16] = buffer_data_1[1967:1960];
        layer3[53][31:24] = buffer_data_1[1975:1968];
        layer3[53][39:32] = buffer_data_1[1983:1976];
        layer4[53][7:0] = buffer_data_0[1951:1944];
        layer4[53][15:8] = buffer_data_0[1959:1952];
        layer4[53][23:16] = buffer_data_0[1967:1960];
        layer4[53][31:24] = buffer_data_0[1975:1968];
        layer4[53][39:32] = buffer_data_0[1983:1976];
        layer0[54][7:0] = buffer_data_4[1959:1952];
        layer0[54][15:8] = buffer_data_4[1967:1960];
        layer0[54][23:16] = buffer_data_4[1975:1968];
        layer0[54][31:24] = buffer_data_4[1983:1976];
        layer0[54][39:32] = buffer_data_4[1991:1984];
        layer1[54][7:0] = buffer_data_3[1959:1952];
        layer1[54][15:8] = buffer_data_3[1967:1960];
        layer1[54][23:16] = buffer_data_3[1975:1968];
        layer1[54][31:24] = buffer_data_3[1983:1976];
        layer1[54][39:32] = buffer_data_3[1991:1984];
        layer2[54][7:0] = buffer_data_2[1959:1952];
        layer2[54][15:8] = buffer_data_2[1967:1960];
        layer2[54][23:16] = buffer_data_2[1975:1968];
        layer2[54][31:24] = buffer_data_2[1983:1976];
        layer2[54][39:32] = buffer_data_2[1991:1984];
        layer3[54][7:0] = buffer_data_1[1959:1952];
        layer3[54][15:8] = buffer_data_1[1967:1960];
        layer3[54][23:16] = buffer_data_1[1975:1968];
        layer3[54][31:24] = buffer_data_1[1983:1976];
        layer3[54][39:32] = buffer_data_1[1991:1984];
        layer4[54][7:0] = buffer_data_0[1959:1952];
        layer4[54][15:8] = buffer_data_0[1967:1960];
        layer4[54][23:16] = buffer_data_0[1975:1968];
        layer4[54][31:24] = buffer_data_0[1983:1976];
        layer4[54][39:32] = buffer_data_0[1991:1984];
        layer0[55][7:0] = buffer_data_4[1967:1960];
        layer0[55][15:8] = buffer_data_4[1975:1968];
        layer0[55][23:16] = buffer_data_4[1983:1976];
        layer0[55][31:24] = buffer_data_4[1991:1984];
        layer0[55][39:32] = buffer_data_4[1999:1992];
        layer1[55][7:0] = buffer_data_3[1967:1960];
        layer1[55][15:8] = buffer_data_3[1975:1968];
        layer1[55][23:16] = buffer_data_3[1983:1976];
        layer1[55][31:24] = buffer_data_3[1991:1984];
        layer1[55][39:32] = buffer_data_3[1999:1992];
        layer2[55][7:0] = buffer_data_2[1967:1960];
        layer2[55][15:8] = buffer_data_2[1975:1968];
        layer2[55][23:16] = buffer_data_2[1983:1976];
        layer2[55][31:24] = buffer_data_2[1991:1984];
        layer2[55][39:32] = buffer_data_2[1999:1992];
        layer3[55][7:0] = buffer_data_1[1967:1960];
        layer3[55][15:8] = buffer_data_1[1975:1968];
        layer3[55][23:16] = buffer_data_1[1983:1976];
        layer3[55][31:24] = buffer_data_1[1991:1984];
        layer3[55][39:32] = buffer_data_1[1999:1992];
        layer4[55][7:0] = buffer_data_0[1967:1960];
        layer4[55][15:8] = buffer_data_0[1975:1968];
        layer4[55][23:16] = buffer_data_0[1983:1976];
        layer4[55][31:24] = buffer_data_0[1991:1984];
        layer4[55][39:32] = buffer_data_0[1999:1992];
        layer0[56][7:0] = buffer_data_4[1975:1968];
        layer0[56][15:8] = buffer_data_4[1983:1976];
        layer0[56][23:16] = buffer_data_4[1991:1984];
        layer0[56][31:24] = buffer_data_4[1999:1992];
        layer0[56][39:32] = buffer_data_4[2007:2000];
        layer1[56][7:0] = buffer_data_3[1975:1968];
        layer1[56][15:8] = buffer_data_3[1983:1976];
        layer1[56][23:16] = buffer_data_3[1991:1984];
        layer1[56][31:24] = buffer_data_3[1999:1992];
        layer1[56][39:32] = buffer_data_3[2007:2000];
        layer2[56][7:0] = buffer_data_2[1975:1968];
        layer2[56][15:8] = buffer_data_2[1983:1976];
        layer2[56][23:16] = buffer_data_2[1991:1984];
        layer2[56][31:24] = buffer_data_2[1999:1992];
        layer2[56][39:32] = buffer_data_2[2007:2000];
        layer3[56][7:0] = buffer_data_1[1975:1968];
        layer3[56][15:8] = buffer_data_1[1983:1976];
        layer3[56][23:16] = buffer_data_1[1991:1984];
        layer3[56][31:24] = buffer_data_1[1999:1992];
        layer3[56][39:32] = buffer_data_1[2007:2000];
        layer4[56][7:0] = buffer_data_0[1975:1968];
        layer4[56][15:8] = buffer_data_0[1983:1976];
        layer4[56][23:16] = buffer_data_0[1991:1984];
        layer4[56][31:24] = buffer_data_0[1999:1992];
        layer4[56][39:32] = buffer_data_0[2007:2000];
        layer0[57][7:0] = buffer_data_4[1983:1976];
        layer0[57][15:8] = buffer_data_4[1991:1984];
        layer0[57][23:16] = buffer_data_4[1999:1992];
        layer0[57][31:24] = buffer_data_4[2007:2000];
        layer0[57][39:32] = buffer_data_4[2015:2008];
        layer1[57][7:0] = buffer_data_3[1983:1976];
        layer1[57][15:8] = buffer_data_3[1991:1984];
        layer1[57][23:16] = buffer_data_3[1999:1992];
        layer1[57][31:24] = buffer_data_3[2007:2000];
        layer1[57][39:32] = buffer_data_3[2015:2008];
        layer2[57][7:0] = buffer_data_2[1983:1976];
        layer2[57][15:8] = buffer_data_2[1991:1984];
        layer2[57][23:16] = buffer_data_2[1999:1992];
        layer2[57][31:24] = buffer_data_2[2007:2000];
        layer2[57][39:32] = buffer_data_2[2015:2008];
        layer3[57][7:0] = buffer_data_1[1983:1976];
        layer3[57][15:8] = buffer_data_1[1991:1984];
        layer3[57][23:16] = buffer_data_1[1999:1992];
        layer3[57][31:24] = buffer_data_1[2007:2000];
        layer3[57][39:32] = buffer_data_1[2015:2008];
        layer4[57][7:0] = buffer_data_0[1983:1976];
        layer4[57][15:8] = buffer_data_0[1991:1984];
        layer4[57][23:16] = buffer_data_0[1999:1992];
        layer4[57][31:24] = buffer_data_0[2007:2000];
        layer4[57][39:32] = buffer_data_0[2015:2008];
        layer0[58][7:0] = buffer_data_4[1991:1984];
        layer0[58][15:8] = buffer_data_4[1999:1992];
        layer0[58][23:16] = buffer_data_4[2007:2000];
        layer0[58][31:24] = buffer_data_4[2015:2008];
        layer0[58][39:32] = buffer_data_4[2023:2016];
        layer1[58][7:0] = buffer_data_3[1991:1984];
        layer1[58][15:8] = buffer_data_3[1999:1992];
        layer1[58][23:16] = buffer_data_3[2007:2000];
        layer1[58][31:24] = buffer_data_3[2015:2008];
        layer1[58][39:32] = buffer_data_3[2023:2016];
        layer2[58][7:0] = buffer_data_2[1991:1984];
        layer2[58][15:8] = buffer_data_2[1999:1992];
        layer2[58][23:16] = buffer_data_2[2007:2000];
        layer2[58][31:24] = buffer_data_2[2015:2008];
        layer2[58][39:32] = buffer_data_2[2023:2016];
        layer3[58][7:0] = buffer_data_1[1991:1984];
        layer3[58][15:8] = buffer_data_1[1999:1992];
        layer3[58][23:16] = buffer_data_1[2007:2000];
        layer3[58][31:24] = buffer_data_1[2015:2008];
        layer3[58][39:32] = buffer_data_1[2023:2016];
        layer4[58][7:0] = buffer_data_0[1991:1984];
        layer4[58][15:8] = buffer_data_0[1999:1992];
        layer4[58][23:16] = buffer_data_0[2007:2000];
        layer4[58][31:24] = buffer_data_0[2015:2008];
        layer4[58][39:32] = buffer_data_0[2023:2016];
        layer0[59][7:0] = buffer_data_4[1999:1992];
        layer0[59][15:8] = buffer_data_4[2007:2000];
        layer0[59][23:16] = buffer_data_4[2015:2008];
        layer0[59][31:24] = buffer_data_4[2023:2016];
        layer0[59][39:32] = buffer_data_4[2031:2024];
        layer1[59][7:0] = buffer_data_3[1999:1992];
        layer1[59][15:8] = buffer_data_3[2007:2000];
        layer1[59][23:16] = buffer_data_3[2015:2008];
        layer1[59][31:24] = buffer_data_3[2023:2016];
        layer1[59][39:32] = buffer_data_3[2031:2024];
        layer2[59][7:0] = buffer_data_2[1999:1992];
        layer2[59][15:8] = buffer_data_2[2007:2000];
        layer2[59][23:16] = buffer_data_2[2015:2008];
        layer2[59][31:24] = buffer_data_2[2023:2016];
        layer2[59][39:32] = buffer_data_2[2031:2024];
        layer3[59][7:0] = buffer_data_1[1999:1992];
        layer3[59][15:8] = buffer_data_1[2007:2000];
        layer3[59][23:16] = buffer_data_1[2015:2008];
        layer3[59][31:24] = buffer_data_1[2023:2016];
        layer3[59][39:32] = buffer_data_1[2031:2024];
        layer4[59][7:0] = buffer_data_0[1999:1992];
        layer4[59][15:8] = buffer_data_0[2007:2000];
        layer4[59][23:16] = buffer_data_0[2015:2008];
        layer4[59][31:24] = buffer_data_0[2023:2016];
        layer4[59][39:32] = buffer_data_0[2031:2024];
        layer0[60][7:0] = buffer_data_4[2007:2000];
        layer0[60][15:8] = buffer_data_4[2015:2008];
        layer0[60][23:16] = buffer_data_4[2023:2016];
        layer0[60][31:24] = buffer_data_4[2031:2024];
        layer0[60][39:32] = buffer_data_4[2039:2032];
        layer1[60][7:0] = buffer_data_3[2007:2000];
        layer1[60][15:8] = buffer_data_3[2015:2008];
        layer1[60][23:16] = buffer_data_3[2023:2016];
        layer1[60][31:24] = buffer_data_3[2031:2024];
        layer1[60][39:32] = buffer_data_3[2039:2032];
        layer2[60][7:0] = buffer_data_2[2007:2000];
        layer2[60][15:8] = buffer_data_2[2015:2008];
        layer2[60][23:16] = buffer_data_2[2023:2016];
        layer2[60][31:24] = buffer_data_2[2031:2024];
        layer2[60][39:32] = buffer_data_2[2039:2032];
        layer3[60][7:0] = buffer_data_1[2007:2000];
        layer3[60][15:8] = buffer_data_1[2015:2008];
        layer3[60][23:16] = buffer_data_1[2023:2016];
        layer3[60][31:24] = buffer_data_1[2031:2024];
        layer3[60][39:32] = buffer_data_1[2039:2032];
        layer4[60][7:0] = buffer_data_0[2007:2000];
        layer4[60][15:8] = buffer_data_0[2015:2008];
        layer4[60][23:16] = buffer_data_0[2023:2016];
        layer4[60][31:24] = buffer_data_0[2031:2024];
        layer4[60][39:32] = buffer_data_0[2039:2032];
        layer0[61][7:0] = buffer_data_4[2015:2008];
        layer0[61][15:8] = buffer_data_4[2023:2016];
        layer0[61][23:16] = buffer_data_4[2031:2024];
        layer0[61][31:24] = buffer_data_4[2039:2032];
        layer0[61][39:32] = buffer_data_4[2047:2040];
        layer1[61][7:0] = buffer_data_3[2015:2008];
        layer1[61][15:8] = buffer_data_3[2023:2016];
        layer1[61][23:16] = buffer_data_3[2031:2024];
        layer1[61][31:24] = buffer_data_3[2039:2032];
        layer1[61][39:32] = buffer_data_3[2047:2040];
        layer2[61][7:0] = buffer_data_2[2015:2008];
        layer2[61][15:8] = buffer_data_2[2023:2016];
        layer2[61][23:16] = buffer_data_2[2031:2024];
        layer2[61][31:24] = buffer_data_2[2039:2032];
        layer2[61][39:32] = buffer_data_2[2047:2040];
        layer3[61][7:0] = buffer_data_1[2015:2008];
        layer3[61][15:8] = buffer_data_1[2023:2016];
        layer3[61][23:16] = buffer_data_1[2031:2024];
        layer3[61][31:24] = buffer_data_1[2039:2032];
        layer3[61][39:32] = buffer_data_1[2047:2040];
        layer4[61][7:0] = buffer_data_0[2015:2008];
        layer4[61][15:8] = buffer_data_0[2023:2016];
        layer4[61][23:16] = buffer_data_0[2031:2024];
        layer4[61][31:24] = buffer_data_0[2039:2032];
        layer4[61][39:32] = buffer_data_0[2047:2040];
        layer0[62][7:0] = buffer_data_4[2023:2016];
        layer0[62][15:8] = buffer_data_4[2031:2024];
        layer0[62][23:16] = buffer_data_4[2039:2032];
        layer0[62][31:24] = buffer_data_4[2047:2040];
        layer0[62][39:32] = buffer_data_4[2055:2048];
        layer1[62][7:0] = buffer_data_3[2023:2016];
        layer1[62][15:8] = buffer_data_3[2031:2024];
        layer1[62][23:16] = buffer_data_3[2039:2032];
        layer1[62][31:24] = buffer_data_3[2047:2040];
        layer1[62][39:32] = buffer_data_3[2055:2048];
        layer2[62][7:0] = buffer_data_2[2023:2016];
        layer2[62][15:8] = buffer_data_2[2031:2024];
        layer2[62][23:16] = buffer_data_2[2039:2032];
        layer2[62][31:24] = buffer_data_2[2047:2040];
        layer2[62][39:32] = buffer_data_2[2055:2048];
        layer3[62][7:0] = buffer_data_1[2023:2016];
        layer3[62][15:8] = buffer_data_1[2031:2024];
        layer3[62][23:16] = buffer_data_1[2039:2032];
        layer3[62][31:24] = buffer_data_1[2047:2040];
        layer3[62][39:32] = buffer_data_1[2055:2048];
        layer4[62][7:0] = buffer_data_0[2023:2016];
        layer4[62][15:8] = buffer_data_0[2031:2024];
        layer4[62][23:16] = buffer_data_0[2039:2032];
        layer4[62][31:24] = buffer_data_0[2047:2040];
        layer4[62][39:32] = buffer_data_0[2055:2048];
        layer0[63][7:0] = buffer_data_4[2031:2024];
        layer0[63][15:8] = buffer_data_4[2039:2032];
        layer0[63][23:16] = buffer_data_4[2047:2040];
        layer0[63][31:24] = buffer_data_4[2055:2048];
        layer0[63][39:32] = buffer_data_4[2063:2056];
        layer1[63][7:0] = buffer_data_3[2031:2024];
        layer1[63][15:8] = buffer_data_3[2039:2032];
        layer1[63][23:16] = buffer_data_3[2047:2040];
        layer1[63][31:24] = buffer_data_3[2055:2048];
        layer1[63][39:32] = buffer_data_3[2063:2056];
        layer2[63][7:0] = buffer_data_2[2031:2024];
        layer2[63][15:8] = buffer_data_2[2039:2032];
        layer2[63][23:16] = buffer_data_2[2047:2040];
        layer2[63][31:24] = buffer_data_2[2055:2048];
        layer2[63][39:32] = buffer_data_2[2063:2056];
        layer3[63][7:0] = buffer_data_1[2031:2024];
        layer3[63][15:8] = buffer_data_1[2039:2032];
        layer3[63][23:16] = buffer_data_1[2047:2040];
        layer3[63][31:24] = buffer_data_1[2055:2048];
        layer3[63][39:32] = buffer_data_1[2063:2056];
        layer4[63][7:0] = buffer_data_0[2031:2024];
        layer4[63][15:8] = buffer_data_0[2039:2032];
        layer4[63][23:16] = buffer_data_0[2047:2040];
        layer4[63][31:24] = buffer_data_0[2055:2048];
        layer4[63][39:32] = buffer_data_0[2063:2056];
    end
    ST_GAUSSIAN_4: begin
        layer0[0][7:0] = buffer_data_4[2039:2032];
        layer0[0][15:8] = buffer_data_4[2047:2040];
        layer0[0][23:16] = buffer_data_4[2055:2048];
        layer0[0][31:24] = buffer_data_4[2063:2056];
        layer0[0][39:32] = buffer_data_4[2071:2064];
        layer1[0][7:0] = buffer_data_3[2039:2032];
        layer1[0][15:8] = buffer_data_3[2047:2040];
        layer1[0][23:16] = buffer_data_3[2055:2048];
        layer1[0][31:24] = buffer_data_3[2063:2056];
        layer1[0][39:32] = buffer_data_3[2071:2064];
        layer2[0][7:0] = buffer_data_2[2039:2032];
        layer2[0][15:8] = buffer_data_2[2047:2040];
        layer2[0][23:16] = buffer_data_2[2055:2048];
        layer2[0][31:24] = buffer_data_2[2063:2056];
        layer2[0][39:32] = buffer_data_2[2071:2064];
        layer3[0][7:0] = buffer_data_1[2039:2032];
        layer3[0][15:8] = buffer_data_1[2047:2040];
        layer3[0][23:16] = buffer_data_1[2055:2048];
        layer3[0][31:24] = buffer_data_1[2063:2056];
        layer3[0][39:32] = buffer_data_1[2071:2064];
        layer4[0][7:0] = buffer_data_0[2039:2032];
        layer4[0][15:8] = buffer_data_0[2047:2040];
        layer4[0][23:16] = buffer_data_0[2055:2048];
        layer4[0][31:24] = buffer_data_0[2063:2056];
        layer4[0][39:32] = buffer_data_0[2071:2064];
        layer0[1][7:0] = buffer_data_4[2047:2040];
        layer0[1][15:8] = buffer_data_4[2055:2048];
        layer0[1][23:16] = buffer_data_4[2063:2056];
        layer0[1][31:24] = buffer_data_4[2071:2064];
        layer0[1][39:32] = buffer_data_4[2079:2072];
        layer1[1][7:0] = buffer_data_3[2047:2040];
        layer1[1][15:8] = buffer_data_3[2055:2048];
        layer1[1][23:16] = buffer_data_3[2063:2056];
        layer1[1][31:24] = buffer_data_3[2071:2064];
        layer1[1][39:32] = buffer_data_3[2079:2072];
        layer2[1][7:0] = buffer_data_2[2047:2040];
        layer2[1][15:8] = buffer_data_2[2055:2048];
        layer2[1][23:16] = buffer_data_2[2063:2056];
        layer2[1][31:24] = buffer_data_2[2071:2064];
        layer2[1][39:32] = buffer_data_2[2079:2072];
        layer3[1][7:0] = buffer_data_1[2047:2040];
        layer3[1][15:8] = buffer_data_1[2055:2048];
        layer3[1][23:16] = buffer_data_1[2063:2056];
        layer3[1][31:24] = buffer_data_1[2071:2064];
        layer3[1][39:32] = buffer_data_1[2079:2072];
        layer4[1][7:0] = buffer_data_0[2047:2040];
        layer4[1][15:8] = buffer_data_0[2055:2048];
        layer4[1][23:16] = buffer_data_0[2063:2056];
        layer4[1][31:24] = buffer_data_0[2071:2064];
        layer4[1][39:32] = buffer_data_0[2079:2072];
        layer0[2][7:0] = buffer_data_4[2055:2048];
        layer0[2][15:8] = buffer_data_4[2063:2056];
        layer0[2][23:16] = buffer_data_4[2071:2064];
        layer0[2][31:24] = buffer_data_4[2079:2072];
        layer0[2][39:32] = buffer_data_4[2087:2080];
        layer1[2][7:0] = buffer_data_3[2055:2048];
        layer1[2][15:8] = buffer_data_3[2063:2056];
        layer1[2][23:16] = buffer_data_3[2071:2064];
        layer1[2][31:24] = buffer_data_3[2079:2072];
        layer1[2][39:32] = buffer_data_3[2087:2080];
        layer2[2][7:0] = buffer_data_2[2055:2048];
        layer2[2][15:8] = buffer_data_2[2063:2056];
        layer2[2][23:16] = buffer_data_2[2071:2064];
        layer2[2][31:24] = buffer_data_2[2079:2072];
        layer2[2][39:32] = buffer_data_2[2087:2080];
        layer3[2][7:0] = buffer_data_1[2055:2048];
        layer3[2][15:8] = buffer_data_1[2063:2056];
        layer3[2][23:16] = buffer_data_1[2071:2064];
        layer3[2][31:24] = buffer_data_1[2079:2072];
        layer3[2][39:32] = buffer_data_1[2087:2080];
        layer4[2][7:0] = buffer_data_0[2055:2048];
        layer4[2][15:8] = buffer_data_0[2063:2056];
        layer4[2][23:16] = buffer_data_0[2071:2064];
        layer4[2][31:24] = buffer_data_0[2079:2072];
        layer4[2][39:32] = buffer_data_0[2087:2080];
        layer0[3][7:0] = buffer_data_4[2063:2056];
        layer0[3][15:8] = buffer_data_4[2071:2064];
        layer0[3][23:16] = buffer_data_4[2079:2072];
        layer0[3][31:24] = buffer_data_4[2087:2080];
        layer0[3][39:32] = buffer_data_4[2095:2088];
        layer1[3][7:0] = buffer_data_3[2063:2056];
        layer1[3][15:8] = buffer_data_3[2071:2064];
        layer1[3][23:16] = buffer_data_3[2079:2072];
        layer1[3][31:24] = buffer_data_3[2087:2080];
        layer1[3][39:32] = buffer_data_3[2095:2088];
        layer2[3][7:0] = buffer_data_2[2063:2056];
        layer2[3][15:8] = buffer_data_2[2071:2064];
        layer2[3][23:16] = buffer_data_2[2079:2072];
        layer2[3][31:24] = buffer_data_2[2087:2080];
        layer2[3][39:32] = buffer_data_2[2095:2088];
        layer3[3][7:0] = buffer_data_1[2063:2056];
        layer3[3][15:8] = buffer_data_1[2071:2064];
        layer3[3][23:16] = buffer_data_1[2079:2072];
        layer3[3][31:24] = buffer_data_1[2087:2080];
        layer3[3][39:32] = buffer_data_1[2095:2088];
        layer4[3][7:0] = buffer_data_0[2063:2056];
        layer4[3][15:8] = buffer_data_0[2071:2064];
        layer4[3][23:16] = buffer_data_0[2079:2072];
        layer4[3][31:24] = buffer_data_0[2087:2080];
        layer4[3][39:32] = buffer_data_0[2095:2088];
        layer0[4][7:0] = buffer_data_4[2071:2064];
        layer0[4][15:8] = buffer_data_4[2079:2072];
        layer0[4][23:16] = buffer_data_4[2087:2080];
        layer0[4][31:24] = buffer_data_4[2095:2088];
        layer0[4][39:32] = buffer_data_4[2103:2096];
        layer1[4][7:0] = buffer_data_3[2071:2064];
        layer1[4][15:8] = buffer_data_3[2079:2072];
        layer1[4][23:16] = buffer_data_3[2087:2080];
        layer1[4][31:24] = buffer_data_3[2095:2088];
        layer1[4][39:32] = buffer_data_3[2103:2096];
        layer2[4][7:0] = buffer_data_2[2071:2064];
        layer2[4][15:8] = buffer_data_2[2079:2072];
        layer2[4][23:16] = buffer_data_2[2087:2080];
        layer2[4][31:24] = buffer_data_2[2095:2088];
        layer2[4][39:32] = buffer_data_2[2103:2096];
        layer3[4][7:0] = buffer_data_1[2071:2064];
        layer3[4][15:8] = buffer_data_1[2079:2072];
        layer3[4][23:16] = buffer_data_1[2087:2080];
        layer3[4][31:24] = buffer_data_1[2095:2088];
        layer3[4][39:32] = buffer_data_1[2103:2096];
        layer4[4][7:0] = buffer_data_0[2071:2064];
        layer4[4][15:8] = buffer_data_0[2079:2072];
        layer4[4][23:16] = buffer_data_0[2087:2080];
        layer4[4][31:24] = buffer_data_0[2095:2088];
        layer4[4][39:32] = buffer_data_0[2103:2096];
        layer0[5][7:0] = buffer_data_4[2079:2072];
        layer0[5][15:8] = buffer_data_4[2087:2080];
        layer0[5][23:16] = buffer_data_4[2095:2088];
        layer0[5][31:24] = buffer_data_4[2103:2096];
        layer0[5][39:32] = buffer_data_4[2111:2104];
        layer1[5][7:0] = buffer_data_3[2079:2072];
        layer1[5][15:8] = buffer_data_3[2087:2080];
        layer1[5][23:16] = buffer_data_3[2095:2088];
        layer1[5][31:24] = buffer_data_3[2103:2096];
        layer1[5][39:32] = buffer_data_3[2111:2104];
        layer2[5][7:0] = buffer_data_2[2079:2072];
        layer2[5][15:8] = buffer_data_2[2087:2080];
        layer2[5][23:16] = buffer_data_2[2095:2088];
        layer2[5][31:24] = buffer_data_2[2103:2096];
        layer2[5][39:32] = buffer_data_2[2111:2104];
        layer3[5][7:0] = buffer_data_1[2079:2072];
        layer3[5][15:8] = buffer_data_1[2087:2080];
        layer3[5][23:16] = buffer_data_1[2095:2088];
        layer3[5][31:24] = buffer_data_1[2103:2096];
        layer3[5][39:32] = buffer_data_1[2111:2104];
        layer4[5][7:0] = buffer_data_0[2079:2072];
        layer4[5][15:8] = buffer_data_0[2087:2080];
        layer4[5][23:16] = buffer_data_0[2095:2088];
        layer4[5][31:24] = buffer_data_0[2103:2096];
        layer4[5][39:32] = buffer_data_0[2111:2104];
        layer0[6][7:0] = buffer_data_4[2087:2080];
        layer0[6][15:8] = buffer_data_4[2095:2088];
        layer0[6][23:16] = buffer_data_4[2103:2096];
        layer0[6][31:24] = buffer_data_4[2111:2104];
        layer0[6][39:32] = buffer_data_4[2119:2112];
        layer1[6][7:0] = buffer_data_3[2087:2080];
        layer1[6][15:8] = buffer_data_3[2095:2088];
        layer1[6][23:16] = buffer_data_3[2103:2096];
        layer1[6][31:24] = buffer_data_3[2111:2104];
        layer1[6][39:32] = buffer_data_3[2119:2112];
        layer2[6][7:0] = buffer_data_2[2087:2080];
        layer2[6][15:8] = buffer_data_2[2095:2088];
        layer2[6][23:16] = buffer_data_2[2103:2096];
        layer2[6][31:24] = buffer_data_2[2111:2104];
        layer2[6][39:32] = buffer_data_2[2119:2112];
        layer3[6][7:0] = buffer_data_1[2087:2080];
        layer3[6][15:8] = buffer_data_1[2095:2088];
        layer3[6][23:16] = buffer_data_1[2103:2096];
        layer3[6][31:24] = buffer_data_1[2111:2104];
        layer3[6][39:32] = buffer_data_1[2119:2112];
        layer4[6][7:0] = buffer_data_0[2087:2080];
        layer4[6][15:8] = buffer_data_0[2095:2088];
        layer4[6][23:16] = buffer_data_0[2103:2096];
        layer4[6][31:24] = buffer_data_0[2111:2104];
        layer4[6][39:32] = buffer_data_0[2119:2112];
        layer0[7][7:0] = buffer_data_4[2095:2088];
        layer0[7][15:8] = buffer_data_4[2103:2096];
        layer0[7][23:16] = buffer_data_4[2111:2104];
        layer0[7][31:24] = buffer_data_4[2119:2112];
        layer0[7][39:32] = buffer_data_4[2127:2120];
        layer1[7][7:0] = buffer_data_3[2095:2088];
        layer1[7][15:8] = buffer_data_3[2103:2096];
        layer1[7][23:16] = buffer_data_3[2111:2104];
        layer1[7][31:24] = buffer_data_3[2119:2112];
        layer1[7][39:32] = buffer_data_3[2127:2120];
        layer2[7][7:0] = buffer_data_2[2095:2088];
        layer2[7][15:8] = buffer_data_2[2103:2096];
        layer2[7][23:16] = buffer_data_2[2111:2104];
        layer2[7][31:24] = buffer_data_2[2119:2112];
        layer2[7][39:32] = buffer_data_2[2127:2120];
        layer3[7][7:0] = buffer_data_1[2095:2088];
        layer3[7][15:8] = buffer_data_1[2103:2096];
        layer3[7][23:16] = buffer_data_1[2111:2104];
        layer3[7][31:24] = buffer_data_1[2119:2112];
        layer3[7][39:32] = buffer_data_1[2127:2120];
        layer4[7][7:0] = buffer_data_0[2095:2088];
        layer4[7][15:8] = buffer_data_0[2103:2096];
        layer4[7][23:16] = buffer_data_0[2111:2104];
        layer4[7][31:24] = buffer_data_0[2119:2112];
        layer4[7][39:32] = buffer_data_0[2127:2120];
        layer0[8][7:0] = buffer_data_4[2103:2096];
        layer0[8][15:8] = buffer_data_4[2111:2104];
        layer0[8][23:16] = buffer_data_4[2119:2112];
        layer0[8][31:24] = buffer_data_4[2127:2120];
        layer0[8][39:32] = buffer_data_4[2135:2128];
        layer1[8][7:0] = buffer_data_3[2103:2096];
        layer1[8][15:8] = buffer_data_3[2111:2104];
        layer1[8][23:16] = buffer_data_3[2119:2112];
        layer1[8][31:24] = buffer_data_3[2127:2120];
        layer1[8][39:32] = buffer_data_3[2135:2128];
        layer2[8][7:0] = buffer_data_2[2103:2096];
        layer2[8][15:8] = buffer_data_2[2111:2104];
        layer2[8][23:16] = buffer_data_2[2119:2112];
        layer2[8][31:24] = buffer_data_2[2127:2120];
        layer2[8][39:32] = buffer_data_2[2135:2128];
        layer3[8][7:0] = buffer_data_1[2103:2096];
        layer3[8][15:8] = buffer_data_1[2111:2104];
        layer3[8][23:16] = buffer_data_1[2119:2112];
        layer3[8][31:24] = buffer_data_1[2127:2120];
        layer3[8][39:32] = buffer_data_1[2135:2128];
        layer4[8][7:0] = buffer_data_0[2103:2096];
        layer4[8][15:8] = buffer_data_0[2111:2104];
        layer4[8][23:16] = buffer_data_0[2119:2112];
        layer4[8][31:24] = buffer_data_0[2127:2120];
        layer4[8][39:32] = buffer_data_0[2135:2128];
        layer0[9][7:0] = buffer_data_4[2111:2104];
        layer0[9][15:8] = buffer_data_4[2119:2112];
        layer0[9][23:16] = buffer_data_4[2127:2120];
        layer0[9][31:24] = buffer_data_4[2135:2128];
        layer0[9][39:32] = buffer_data_4[2143:2136];
        layer1[9][7:0] = buffer_data_3[2111:2104];
        layer1[9][15:8] = buffer_data_3[2119:2112];
        layer1[9][23:16] = buffer_data_3[2127:2120];
        layer1[9][31:24] = buffer_data_3[2135:2128];
        layer1[9][39:32] = buffer_data_3[2143:2136];
        layer2[9][7:0] = buffer_data_2[2111:2104];
        layer2[9][15:8] = buffer_data_2[2119:2112];
        layer2[9][23:16] = buffer_data_2[2127:2120];
        layer2[9][31:24] = buffer_data_2[2135:2128];
        layer2[9][39:32] = buffer_data_2[2143:2136];
        layer3[9][7:0] = buffer_data_1[2111:2104];
        layer3[9][15:8] = buffer_data_1[2119:2112];
        layer3[9][23:16] = buffer_data_1[2127:2120];
        layer3[9][31:24] = buffer_data_1[2135:2128];
        layer3[9][39:32] = buffer_data_1[2143:2136];
        layer4[9][7:0] = buffer_data_0[2111:2104];
        layer4[9][15:8] = buffer_data_0[2119:2112];
        layer4[9][23:16] = buffer_data_0[2127:2120];
        layer4[9][31:24] = buffer_data_0[2135:2128];
        layer4[9][39:32] = buffer_data_0[2143:2136];
        layer0[10][7:0] = buffer_data_4[2119:2112];
        layer0[10][15:8] = buffer_data_4[2127:2120];
        layer0[10][23:16] = buffer_data_4[2135:2128];
        layer0[10][31:24] = buffer_data_4[2143:2136];
        layer0[10][39:32] = buffer_data_4[2151:2144];
        layer1[10][7:0] = buffer_data_3[2119:2112];
        layer1[10][15:8] = buffer_data_3[2127:2120];
        layer1[10][23:16] = buffer_data_3[2135:2128];
        layer1[10][31:24] = buffer_data_3[2143:2136];
        layer1[10][39:32] = buffer_data_3[2151:2144];
        layer2[10][7:0] = buffer_data_2[2119:2112];
        layer2[10][15:8] = buffer_data_2[2127:2120];
        layer2[10][23:16] = buffer_data_2[2135:2128];
        layer2[10][31:24] = buffer_data_2[2143:2136];
        layer2[10][39:32] = buffer_data_2[2151:2144];
        layer3[10][7:0] = buffer_data_1[2119:2112];
        layer3[10][15:8] = buffer_data_1[2127:2120];
        layer3[10][23:16] = buffer_data_1[2135:2128];
        layer3[10][31:24] = buffer_data_1[2143:2136];
        layer3[10][39:32] = buffer_data_1[2151:2144];
        layer4[10][7:0] = buffer_data_0[2119:2112];
        layer4[10][15:8] = buffer_data_0[2127:2120];
        layer4[10][23:16] = buffer_data_0[2135:2128];
        layer4[10][31:24] = buffer_data_0[2143:2136];
        layer4[10][39:32] = buffer_data_0[2151:2144];
        layer0[11][7:0] = buffer_data_4[2127:2120];
        layer0[11][15:8] = buffer_data_4[2135:2128];
        layer0[11][23:16] = buffer_data_4[2143:2136];
        layer0[11][31:24] = buffer_data_4[2151:2144];
        layer0[11][39:32] = buffer_data_4[2159:2152];
        layer1[11][7:0] = buffer_data_3[2127:2120];
        layer1[11][15:8] = buffer_data_3[2135:2128];
        layer1[11][23:16] = buffer_data_3[2143:2136];
        layer1[11][31:24] = buffer_data_3[2151:2144];
        layer1[11][39:32] = buffer_data_3[2159:2152];
        layer2[11][7:0] = buffer_data_2[2127:2120];
        layer2[11][15:8] = buffer_data_2[2135:2128];
        layer2[11][23:16] = buffer_data_2[2143:2136];
        layer2[11][31:24] = buffer_data_2[2151:2144];
        layer2[11][39:32] = buffer_data_2[2159:2152];
        layer3[11][7:0] = buffer_data_1[2127:2120];
        layer3[11][15:8] = buffer_data_1[2135:2128];
        layer3[11][23:16] = buffer_data_1[2143:2136];
        layer3[11][31:24] = buffer_data_1[2151:2144];
        layer3[11][39:32] = buffer_data_1[2159:2152];
        layer4[11][7:0] = buffer_data_0[2127:2120];
        layer4[11][15:8] = buffer_data_0[2135:2128];
        layer4[11][23:16] = buffer_data_0[2143:2136];
        layer4[11][31:24] = buffer_data_0[2151:2144];
        layer4[11][39:32] = buffer_data_0[2159:2152];
        layer0[12][7:0] = buffer_data_4[2135:2128];
        layer0[12][15:8] = buffer_data_4[2143:2136];
        layer0[12][23:16] = buffer_data_4[2151:2144];
        layer0[12][31:24] = buffer_data_4[2159:2152];
        layer0[12][39:32] = buffer_data_4[2167:2160];
        layer1[12][7:0] = buffer_data_3[2135:2128];
        layer1[12][15:8] = buffer_data_3[2143:2136];
        layer1[12][23:16] = buffer_data_3[2151:2144];
        layer1[12][31:24] = buffer_data_3[2159:2152];
        layer1[12][39:32] = buffer_data_3[2167:2160];
        layer2[12][7:0] = buffer_data_2[2135:2128];
        layer2[12][15:8] = buffer_data_2[2143:2136];
        layer2[12][23:16] = buffer_data_2[2151:2144];
        layer2[12][31:24] = buffer_data_2[2159:2152];
        layer2[12][39:32] = buffer_data_2[2167:2160];
        layer3[12][7:0] = buffer_data_1[2135:2128];
        layer3[12][15:8] = buffer_data_1[2143:2136];
        layer3[12][23:16] = buffer_data_1[2151:2144];
        layer3[12][31:24] = buffer_data_1[2159:2152];
        layer3[12][39:32] = buffer_data_1[2167:2160];
        layer4[12][7:0] = buffer_data_0[2135:2128];
        layer4[12][15:8] = buffer_data_0[2143:2136];
        layer4[12][23:16] = buffer_data_0[2151:2144];
        layer4[12][31:24] = buffer_data_0[2159:2152];
        layer4[12][39:32] = buffer_data_0[2167:2160];
        layer0[13][7:0] = buffer_data_4[2143:2136];
        layer0[13][15:8] = buffer_data_4[2151:2144];
        layer0[13][23:16] = buffer_data_4[2159:2152];
        layer0[13][31:24] = buffer_data_4[2167:2160];
        layer0[13][39:32] = buffer_data_4[2175:2168];
        layer1[13][7:0] = buffer_data_3[2143:2136];
        layer1[13][15:8] = buffer_data_3[2151:2144];
        layer1[13][23:16] = buffer_data_3[2159:2152];
        layer1[13][31:24] = buffer_data_3[2167:2160];
        layer1[13][39:32] = buffer_data_3[2175:2168];
        layer2[13][7:0] = buffer_data_2[2143:2136];
        layer2[13][15:8] = buffer_data_2[2151:2144];
        layer2[13][23:16] = buffer_data_2[2159:2152];
        layer2[13][31:24] = buffer_data_2[2167:2160];
        layer2[13][39:32] = buffer_data_2[2175:2168];
        layer3[13][7:0] = buffer_data_1[2143:2136];
        layer3[13][15:8] = buffer_data_1[2151:2144];
        layer3[13][23:16] = buffer_data_1[2159:2152];
        layer3[13][31:24] = buffer_data_1[2167:2160];
        layer3[13][39:32] = buffer_data_1[2175:2168];
        layer4[13][7:0] = buffer_data_0[2143:2136];
        layer4[13][15:8] = buffer_data_0[2151:2144];
        layer4[13][23:16] = buffer_data_0[2159:2152];
        layer4[13][31:24] = buffer_data_0[2167:2160];
        layer4[13][39:32] = buffer_data_0[2175:2168];
        layer0[14][7:0] = buffer_data_4[2151:2144];
        layer0[14][15:8] = buffer_data_4[2159:2152];
        layer0[14][23:16] = buffer_data_4[2167:2160];
        layer0[14][31:24] = buffer_data_4[2175:2168];
        layer0[14][39:32] = buffer_data_4[2183:2176];
        layer1[14][7:0] = buffer_data_3[2151:2144];
        layer1[14][15:8] = buffer_data_3[2159:2152];
        layer1[14][23:16] = buffer_data_3[2167:2160];
        layer1[14][31:24] = buffer_data_3[2175:2168];
        layer1[14][39:32] = buffer_data_3[2183:2176];
        layer2[14][7:0] = buffer_data_2[2151:2144];
        layer2[14][15:8] = buffer_data_2[2159:2152];
        layer2[14][23:16] = buffer_data_2[2167:2160];
        layer2[14][31:24] = buffer_data_2[2175:2168];
        layer2[14][39:32] = buffer_data_2[2183:2176];
        layer3[14][7:0] = buffer_data_1[2151:2144];
        layer3[14][15:8] = buffer_data_1[2159:2152];
        layer3[14][23:16] = buffer_data_1[2167:2160];
        layer3[14][31:24] = buffer_data_1[2175:2168];
        layer3[14][39:32] = buffer_data_1[2183:2176];
        layer4[14][7:0] = buffer_data_0[2151:2144];
        layer4[14][15:8] = buffer_data_0[2159:2152];
        layer4[14][23:16] = buffer_data_0[2167:2160];
        layer4[14][31:24] = buffer_data_0[2175:2168];
        layer4[14][39:32] = buffer_data_0[2183:2176];
        layer0[15][7:0] = buffer_data_4[2159:2152];
        layer0[15][15:8] = buffer_data_4[2167:2160];
        layer0[15][23:16] = buffer_data_4[2175:2168];
        layer0[15][31:24] = buffer_data_4[2183:2176];
        layer0[15][39:32] = buffer_data_4[2191:2184];
        layer1[15][7:0] = buffer_data_3[2159:2152];
        layer1[15][15:8] = buffer_data_3[2167:2160];
        layer1[15][23:16] = buffer_data_3[2175:2168];
        layer1[15][31:24] = buffer_data_3[2183:2176];
        layer1[15][39:32] = buffer_data_3[2191:2184];
        layer2[15][7:0] = buffer_data_2[2159:2152];
        layer2[15][15:8] = buffer_data_2[2167:2160];
        layer2[15][23:16] = buffer_data_2[2175:2168];
        layer2[15][31:24] = buffer_data_2[2183:2176];
        layer2[15][39:32] = buffer_data_2[2191:2184];
        layer3[15][7:0] = buffer_data_1[2159:2152];
        layer3[15][15:8] = buffer_data_1[2167:2160];
        layer3[15][23:16] = buffer_data_1[2175:2168];
        layer3[15][31:24] = buffer_data_1[2183:2176];
        layer3[15][39:32] = buffer_data_1[2191:2184];
        layer4[15][7:0] = buffer_data_0[2159:2152];
        layer4[15][15:8] = buffer_data_0[2167:2160];
        layer4[15][23:16] = buffer_data_0[2175:2168];
        layer4[15][31:24] = buffer_data_0[2183:2176];
        layer4[15][39:32] = buffer_data_0[2191:2184];
        layer0[16][7:0] = buffer_data_4[2167:2160];
        layer0[16][15:8] = buffer_data_4[2175:2168];
        layer0[16][23:16] = buffer_data_4[2183:2176];
        layer0[16][31:24] = buffer_data_4[2191:2184];
        layer0[16][39:32] = buffer_data_4[2199:2192];
        layer1[16][7:0] = buffer_data_3[2167:2160];
        layer1[16][15:8] = buffer_data_3[2175:2168];
        layer1[16][23:16] = buffer_data_3[2183:2176];
        layer1[16][31:24] = buffer_data_3[2191:2184];
        layer1[16][39:32] = buffer_data_3[2199:2192];
        layer2[16][7:0] = buffer_data_2[2167:2160];
        layer2[16][15:8] = buffer_data_2[2175:2168];
        layer2[16][23:16] = buffer_data_2[2183:2176];
        layer2[16][31:24] = buffer_data_2[2191:2184];
        layer2[16][39:32] = buffer_data_2[2199:2192];
        layer3[16][7:0] = buffer_data_1[2167:2160];
        layer3[16][15:8] = buffer_data_1[2175:2168];
        layer3[16][23:16] = buffer_data_1[2183:2176];
        layer3[16][31:24] = buffer_data_1[2191:2184];
        layer3[16][39:32] = buffer_data_1[2199:2192];
        layer4[16][7:0] = buffer_data_0[2167:2160];
        layer4[16][15:8] = buffer_data_0[2175:2168];
        layer4[16][23:16] = buffer_data_0[2183:2176];
        layer4[16][31:24] = buffer_data_0[2191:2184];
        layer4[16][39:32] = buffer_data_0[2199:2192];
        layer0[17][7:0] = buffer_data_4[2175:2168];
        layer0[17][15:8] = buffer_data_4[2183:2176];
        layer0[17][23:16] = buffer_data_4[2191:2184];
        layer0[17][31:24] = buffer_data_4[2199:2192];
        layer0[17][39:32] = buffer_data_4[2207:2200];
        layer1[17][7:0] = buffer_data_3[2175:2168];
        layer1[17][15:8] = buffer_data_3[2183:2176];
        layer1[17][23:16] = buffer_data_3[2191:2184];
        layer1[17][31:24] = buffer_data_3[2199:2192];
        layer1[17][39:32] = buffer_data_3[2207:2200];
        layer2[17][7:0] = buffer_data_2[2175:2168];
        layer2[17][15:8] = buffer_data_2[2183:2176];
        layer2[17][23:16] = buffer_data_2[2191:2184];
        layer2[17][31:24] = buffer_data_2[2199:2192];
        layer2[17][39:32] = buffer_data_2[2207:2200];
        layer3[17][7:0] = buffer_data_1[2175:2168];
        layer3[17][15:8] = buffer_data_1[2183:2176];
        layer3[17][23:16] = buffer_data_1[2191:2184];
        layer3[17][31:24] = buffer_data_1[2199:2192];
        layer3[17][39:32] = buffer_data_1[2207:2200];
        layer4[17][7:0] = buffer_data_0[2175:2168];
        layer4[17][15:8] = buffer_data_0[2183:2176];
        layer4[17][23:16] = buffer_data_0[2191:2184];
        layer4[17][31:24] = buffer_data_0[2199:2192];
        layer4[17][39:32] = buffer_data_0[2207:2200];
        layer0[18][7:0] = buffer_data_4[2183:2176];
        layer0[18][15:8] = buffer_data_4[2191:2184];
        layer0[18][23:16] = buffer_data_4[2199:2192];
        layer0[18][31:24] = buffer_data_4[2207:2200];
        layer0[18][39:32] = buffer_data_4[2215:2208];
        layer1[18][7:0] = buffer_data_3[2183:2176];
        layer1[18][15:8] = buffer_data_3[2191:2184];
        layer1[18][23:16] = buffer_data_3[2199:2192];
        layer1[18][31:24] = buffer_data_3[2207:2200];
        layer1[18][39:32] = buffer_data_3[2215:2208];
        layer2[18][7:0] = buffer_data_2[2183:2176];
        layer2[18][15:8] = buffer_data_2[2191:2184];
        layer2[18][23:16] = buffer_data_2[2199:2192];
        layer2[18][31:24] = buffer_data_2[2207:2200];
        layer2[18][39:32] = buffer_data_2[2215:2208];
        layer3[18][7:0] = buffer_data_1[2183:2176];
        layer3[18][15:8] = buffer_data_1[2191:2184];
        layer3[18][23:16] = buffer_data_1[2199:2192];
        layer3[18][31:24] = buffer_data_1[2207:2200];
        layer3[18][39:32] = buffer_data_1[2215:2208];
        layer4[18][7:0] = buffer_data_0[2183:2176];
        layer4[18][15:8] = buffer_data_0[2191:2184];
        layer4[18][23:16] = buffer_data_0[2199:2192];
        layer4[18][31:24] = buffer_data_0[2207:2200];
        layer4[18][39:32] = buffer_data_0[2215:2208];
        layer0[19][7:0] = buffer_data_4[2191:2184];
        layer0[19][15:8] = buffer_data_4[2199:2192];
        layer0[19][23:16] = buffer_data_4[2207:2200];
        layer0[19][31:24] = buffer_data_4[2215:2208];
        layer0[19][39:32] = buffer_data_4[2223:2216];
        layer1[19][7:0] = buffer_data_3[2191:2184];
        layer1[19][15:8] = buffer_data_3[2199:2192];
        layer1[19][23:16] = buffer_data_3[2207:2200];
        layer1[19][31:24] = buffer_data_3[2215:2208];
        layer1[19][39:32] = buffer_data_3[2223:2216];
        layer2[19][7:0] = buffer_data_2[2191:2184];
        layer2[19][15:8] = buffer_data_2[2199:2192];
        layer2[19][23:16] = buffer_data_2[2207:2200];
        layer2[19][31:24] = buffer_data_2[2215:2208];
        layer2[19][39:32] = buffer_data_2[2223:2216];
        layer3[19][7:0] = buffer_data_1[2191:2184];
        layer3[19][15:8] = buffer_data_1[2199:2192];
        layer3[19][23:16] = buffer_data_1[2207:2200];
        layer3[19][31:24] = buffer_data_1[2215:2208];
        layer3[19][39:32] = buffer_data_1[2223:2216];
        layer4[19][7:0] = buffer_data_0[2191:2184];
        layer4[19][15:8] = buffer_data_0[2199:2192];
        layer4[19][23:16] = buffer_data_0[2207:2200];
        layer4[19][31:24] = buffer_data_0[2215:2208];
        layer4[19][39:32] = buffer_data_0[2223:2216];
        layer0[20][7:0] = buffer_data_4[2199:2192];
        layer0[20][15:8] = buffer_data_4[2207:2200];
        layer0[20][23:16] = buffer_data_4[2215:2208];
        layer0[20][31:24] = buffer_data_4[2223:2216];
        layer0[20][39:32] = buffer_data_4[2231:2224];
        layer1[20][7:0] = buffer_data_3[2199:2192];
        layer1[20][15:8] = buffer_data_3[2207:2200];
        layer1[20][23:16] = buffer_data_3[2215:2208];
        layer1[20][31:24] = buffer_data_3[2223:2216];
        layer1[20][39:32] = buffer_data_3[2231:2224];
        layer2[20][7:0] = buffer_data_2[2199:2192];
        layer2[20][15:8] = buffer_data_2[2207:2200];
        layer2[20][23:16] = buffer_data_2[2215:2208];
        layer2[20][31:24] = buffer_data_2[2223:2216];
        layer2[20][39:32] = buffer_data_2[2231:2224];
        layer3[20][7:0] = buffer_data_1[2199:2192];
        layer3[20][15:8] = buffer_data_1[2207:2200];
        layer3[20][23:16] = buffer_data_1[2215:2208];
        layer3[20][31:24] = buffer_data_1[2223:2216];
        layer3[20][39:32] = buffer_data_1[2231:2224];
        layer4[20][7:0] = buffer_data_0[2199:2192];
        layer4[20][15:8] = buffer_data_0[2207:2200];
        layer4[20][23:16] = buffer_data_0[2215:2208];
        layer4[20][31:24] = buffer_data_0[2223:2216];
        layer4[20][39:32] = buffer_data_0[2231:2224];
        layer0[21][7:0] = buffer_data_4[2207:2200];
        layer0[21][15:8] = buffer_data_4[2215:2208];
        layer0[21][23:16] = buffer_data_4[2223:2216];
        layer0[21][31:24] = buffer_data_4[2231:2224];
        layer0[21][39:32] = buffer_data_4[2239:2232];
        layer1[21][7:0] = buffer_data_3[2207:2200];
        layer1[21][15:8] = buffer_data_3[2215:2208];
        layer1[21][23:16] = buffer_data_3[2223:2216];
        layer1[21][31:24] = buffer_data_3[2231:2224];
        layer1[21][39:32] = buffer_data_3[2239:2232];
        layer2[21][7:0] = buffer_data_2[2207:2200];
        layer2[21][15:8] = buffer_data_2[2215:2208];
        layer2[21][23:16] = buffer_data_2[2223:2216];
        layer2[21][31:24] = buffer_data_2[2231:2224];
        layer2[21][39:32] = buffer_data_2[2239:2232];
        layer3[21][7:0] = buffer_data_1[2207:2200];
        layer3[21][15:8] = buffer_data_1[2215:2208];
        layer3[21][23:16] = buffer_data_1[2223:2216];
        layer3[21][31:24] = buffer_data_1[2231:2224];
        layer3[21][39:32] = buffer_data_1[2239:2232];
        layer4[21][7:0] = buffer_data_0[2207:2200];
        layer4[21][15:8] = buffer_data_0[2215:2208];
        layer4[21][23:16] = buffer_data_0[2223:2216];
        layer4[21][31:24] = buffer_data_0[2231:2224];
        layer4[21][39:32] = buffer_data_0[2239:2232];
        layer0[22][7:0] = buffer_data_4[2215:2208];
        layer0[22][15:8] = buffer_data_4[2223:2216];
        layer0[22][23:16] = buffer_data_4[2231:2224];
        layer0[22][31:24] = buffer_data_4[2239:2232];
        layer0[22][39:32] = buffer_data_4[2247:2240];
        layer1[22][7:0] = buffer_data_3[2215:2208];
        layer1[22][15:8] = buffer_data_3[2223:2216];
        layer1[22][23:16] = buffer_data_3[2231:2224];
        layer1[22][31:24] = buffer_data_3[2239:2232];
        layer1[22][39:32] = buffer_data_3[2247:2240];
        layer2[22][7:0] = buffer_data_2[2215:2208];
        layer2[22][15:8] = buffer_data_2[2223:2216];
        layer2[22][23:16] = buffer_data_2[2231:2224];
        layer2[22][31:24] = buffer_data_2[2239:2232];
        layer2[22][39:32] = buffer_data_2[2247:2240];
        layer3[22][7:0] = buffer_data_1[2215:2208];
        layer3[22][15:8] = buffer_data_1[2223:2216];
        layer3[22][23:16] = buffer_data_1[2231:2224];
        layer3[22][31:24] = buffer_data_1[2239:2232];
        layer3[22][39:32] = buffer_data_1[2247:2240];
        layer4[22][7:0] = buffer_data_0[2215:2208];
        layer4[22][15:8] = buffer_data_0[2223:2216];
        layer4[22][23:16] = buffer_data_0[2231:2224];
        layer4[22][31:24] = buffer_data_0[2239:2232];
        layer4[22][39:32] = buffer_data_0[2247:2240];
        layer0[23][7:0] = buffer_data_4[2223:2216];
        layer0[23][15:8] = buffer_data_4[2231:2224];
        layer0[23][23:16] = buffer_data_4[2239:2232];
        layer0[23][31:24] = buffer_data_4[2247:2240];
        layer0[23][39:32] = buffer_data_4[2255:2248];
        layer1[23][7:0] = buffer_data_3[2223:2216];
        layer1[23][15:8] = buffer_data_3[2231:2224];
        layer1[23][23:16] = buffer_data_3[2239:2232];
        layer1[23][31:24] = buffer_data_3[2247:2240];
        layer1[23][39:32] = buffer_data_3[2255:2248];
        layer2[23][7:0] = buffer_data_2[2223:2216];
        layer2[23][15:8] = buffer_data_2[2231:2224];
        layer2[23][23:16] = buffer_data_2[2239:2232];
        layer2[23][31:24] = buffer_data_2[2247:2240];
        layer2[23][39:32] = buffer_data_2[2255:2248];
        layer3[23][7:0] = buffer_data_1[2223:2216];
        layer3[23][15:8] = buffer_data_1[2231:2224];
        layer3[23][23:16] = buffer_data_1[2239:2232];
        layer3[23][31:24] = buffer_data_1[2247:2240];
        layer3[23][39:32] = buffer_data_1[2255:2248];
        layer4[23][7:0] = buffer_data_0[2223:2216];
        layer4[23][15:8] = buffer_data_0[2231:2224];
        layer4[23][23:16] = buffer_data_0[2239:2232];
        layer4[23][31:24] = buffer_data_0[2247:2240];
        layer4[23][39:32] = buffer_data_0[2255:2248];
        layer0[24][7:0] = buffer_data_4[2231:2224];
        layer0[24][15:8] = buffer_data_4[2239:2232];
        layer0[24][23:16] = buffer_data_4[2247:2240];
        layer0[24][31:24] = buffer_data_4[2255:2248];
        layer0[24][39:32] = buffer_data_4[2263:2256];
        layer1[24][7:0] = buffer_data_3[2231:2224];
        layer1[24][15:8] = buffer_data_3[2239:2232];
        layer1[24][23:16] = buffer_data_3[2247:2240];
        layer1[24][31:24] = buffer_data_3[2255:2248];
        layer1[24][39:32] = buffer_data_3[2263:2256];
        layer2[24][7:0] = buffer_data_2[2231:2224];
        layer2[24][15:8] = buffer_data_2[2239:2232];
        layer2[24][23:16] = buffer_data_2[2247:2240];
        layer2[24][31:24] = buffer_data_2[2255:2248];
        layer2[24][39:32] = buffer_data_2[2263:2256];
        layer3[24][7:0] = buffer_data_1[2231:2224];
        layer3[24][15:8] = buffer_data_1[2239:2232];
        layer3[24][23:16] = buffer_data_1[2247:2240];
        layer3[24][31:24] = buffer_data_1[2255:2248];
        layer3[24][39:32] = buffer_data_1[2263:2256];
        layer4[24][7:0] = buffer_data_0[2231:2224];
        layer4[24][15:8] = buffer_data_0[2239:2232];
        layer4[24][23:16] = buffer_data_0[2247:2240];
        layer4[24][31:24] = buffer_data_0[2255:2248];
        layer4[24][39:32] = buffer_data_0[2263:2256];
        layer0[25][7:0] = buffer_data_4[2239:2232];
        layer0[25][15:8] = buffer_data_4[2247:2240];
        layer0[25][23:16] = buffer_data_4[2255:2248];
        layer0[25][31:24] = buffer_data_4[2263:2256];
        layer0[25][39:32] = buffer_data_4[2271:2264];
        layer1[25][7:0] = buffer_data_3[2239:2232];
        layer1[25][15:8] = buffer_data_3[2247:2240];
        layer1[25][23:16] = buffer_data_3[2255:2248];
        layer1[25][31:24] = buffer_data_3[2263:2256];
        layer1[25][39:32] = buffer_data_3[2271:2264];
        layer2[25][7:0] = buffer_data_2[2239:2232];
        layer2[25][15:8] = buffer_data_2[2247:2240];
        layer2[25][23:16] = buffer_data_2[2255:2248];
        layer2[25][31:24] = buffer_data_2[2263:2256];
        layer2[25][39:32] = buffer_data_2[2271:2264];
        layer3[25][7:0] = buffer_data_1[2239:2232];
        layer3[25][15:8] = buffer_data_1[2247:2240];
        layer3[25][23:16] = buffer_data_1[2255:2248];
        layer3[25][31:24] = buffer_data_1[2263:2256];
        layer3[25][39:32] = buffer_data_1[2271:2264];
        layer4[25][7:0] = buffer_data_0[2239:2232];
        layer4[25][15:8] = buffer_data_0[2247:2240];
        layer4[25][23:16] = buffer_data_0[2255:2248];
        layer4[25][31:24] = buffer_data_0[2263:2256];
        layer4[25][39:32] = buffer_data_0[2271:2264];
        layer0[26][7:0] = buffer_data_4[2247:2240];
        layer0[26][15:8] = buffer_data_4[2255:2248];
        layer0[26][23:16] = buffer_data_4[2263:2256];
        layer0[26][31:24] = buffer_data_4[2271:2264];
        layer0[26][39:32] = buffer_data_4[2279:2272];
        layer1[26][7:0] = buffer_data_3[2247:2240];
        layer1[26][15:8] = buffer_data_3[2255:2248];
        layer1[26][23:16] = buffer_data_3[2263:2256];
        layer1[26][31:24] = buffer_data_3[2271:2264];
        layer1[26][39:32] = buffer_data_3[2279:2272];
        layer2[26][7:0] = buffer_data_2[2247:2240];
        layer2[26][15:8] = buffer_data_2[2255:2248];
        layer2[26][23:16] = buffer_data_2[2263:2256];
        layer2[26][31:24] = buffer_data_2[2271:2264];
        layer2[26][39:32] = buffer_data_2[2279:2272];
        layer3[26][7:0] = buffer_data_1[2247:2240];
        layer3[26][15:8] = buffer_data_1[2255:2248];
        layer3[26][23:16] = buffer_data_1[2263:2256];
        layer3[26][31:24] = buffer_data_1[2271:2264];
        layer3[26][39:32] = buffer_data_1[2279:2272];
        layer4[26][7:0] = buffer_data_0[2247:2240];
        layer4[26][15:8] = buffer_data_0[2255:2248];
        layer4[26][23:16] = buffer_data_0[2263:2256];
        layer4[26][31:24] = buffer_data_0[2271:2264];
        layer4[26][39:32] = buffer_data_0[2279:2272];
        layer0[27][7:0] = buffer_data_4[2255:2248];
        layer0[27][15:8] = buffer_data_4[2263:2256];
        layer0[27][23:16] = buffer_data_4[2271:2264];
        layer0[27][31:24] = buffer_data_4[2279:2272];
        layer0[27][39:32] = buffer_data_4[2287:2280];
        layer1[27][7:0] = buffer_data_3[2255:2248];
        layer1[27][15:8] = buffer_data_3[2263:2256];
        layer1[27][23:16] = buffer_data_3[2271:2264];
        layer1[27][31:24] = buffer_data_3[2279:2272];
        layer1[27][39:32] = buffer_data_3[2287:2280];
        layer2[27][7:0] = buffer_data_2[2255:2248];
        layer2[27][15:8] = buffer_data_2[2263:2256];
        layer2[27][23:16] = buffer_data_2[2271:2264];
        layer2[27][31:24] = buffer_data_2[2279:2272];
        layer2[27][39:32] = buffer_data_2[2287:2280];
        layer3[27][7:0] = buffer_data_1[2255:2248];
        layer3[27][15:8] = buffer_data_1[2263:2256];
        layer3[27][23:16] = buffer_data_1[2271:2264];
        layer3[27][31:24] = buffer_data_1[2279:2272];
        layer3[27][39:32] = buffer_data_1[2287:2280];
        layer4[27][7:0] = buffer_data_0[2255:2248];
        layer4[27][15:8] = buffer_data_0[2263:2256];
        layer4[27][23:16] = buffer_data_0[2271:2264];
        layer4[27][31:24] = buffer_data_0[2279:2272];
        layer4[27][39:32] = buffer_data_0[2287:2280];
        layer0[28][7:0] = buffer_data_4[2263:2256];
        layer0[28][15:8] = buffer_data_4[2271:2264];
        layer0[28][23:16] = buffer_data_4[2279:2272];
        layer0[28][31:24] = buffer_data_4[2287:2280];
        layer0[28][39:32] = buffer_data_4[2295:2288];
        layer1[28][7:0] = buffer_data_3[2263:2256];
        layer1[28][15:8] = buffer_data_3[2271:2264];
        layer1[28][23:16] = buffer_data_3[2279:2272];
        layer1[28][31:24] = buffer_data_3[2287:2280];
        layer1[28][39:32] = buffer_data_3[2295:2288];
        layer2[28][7:0] = buffer_data_2[2263:2256];
        layer2[28][15:8] = buffer_data_2[2271:2264];
        layer2[28][23:16] = buffer_data_2[2279:2272];
        layer2[28][31:24] = buffer_data_2[2287:2280];
        layer2[28][39:32] = buffer_data_2[2295:2288];
        layer3[28][7:0] = buffer_data_1[2263:2256];
        layer3[28][15:8] = buffer_data_1[2271:2264];
        layer3[28][23:16] = buffer_data_1[2279:2272];
        layer3[28][31:24] = buffer_data_1[2287:2280];
        layer3[28][39:32] = buffer_data_1[2295:2288];
        layer4[28][7:0] = buffer_data_0[2263:2256];
        layer4[28][15:8] = buffer_data_0[2271:2264];
        layer4[28][23:16] = buffer_data_0[2279:2272];
        layer4[28][31:24] = buffer_data_0[2287:2280];
        layer4[28][39:32] = buffer_data_0[2295:2288];
        layer0[29][7:0] = buffer_data_4[2271:2264];
        layer0[29][15:8] = buffer_data_4[2279:2272];
        layer0[29][23:16] = buffer_data_4[2287:2280];
        layer0[29][31:24] = buffer_data_4[2295:2288];
        layer0[29][39:32] = buffer_data_4[2303:2296];
        layer1[29][7:0] = buffer_data_3[2271:2264];
        layer1[29][15:8] = buffer_data_3[2279:2272];
        layer1[29][23:16] = buffer_data_3[2287:2280];
        layer1[29][31:24] = buffer_data_3[2295:2288];
        layer1[29][39:32] = buffer_data_3[2303:2296];
        layer2[29][7:0] = buffer_data_2[2271:2264];
        layer2[29][15:8] = buffer_data_2[2279:2272];
        layer2[29][23:16] = buffer_data_2[2287:2280];
        layer2[29][31:24] = buffer_data_2[2295:2288];
        layer2[29][39:32] = buffer_data_2[2303:2296];
        layer3[29][7:0] = buffer_data_1[2271:2264];
        layer3[29][15:8] = buffer_data_1[2279:2272];
        layer3[29][23:16] = buffer_data_1[2287:2280];
        layer3[29][31:24] = buffer_data_1[2295:2288];
        layer3[29][39:32] = buffer_data_1[2303:2296];
        layer4[29][7:0] = buffer_data_0[2271:2264];
        layer4[29][15:8] = buffer_data_0[2279:2272];
        layer4[29][23:16] = buffer_data_0[2287:2280];
        layer4[29][31:24] = buffer_data_0[2295:2288];
        layer4[29][39:32] = buffer_data_0[2303:2296];
        layer0[30][7:0] = buffer_data_4[2279:2272];
        layer0[30][15:8] = buffer_data_4[2287:2280];
        layer0[30][23:16] = buffer_data_4[2295:2288];
        layer0[30][31:24] = buffer_data_4[2303:2296];
        layer0[30][39:32] = buffer_data_4[2311:2304];
        layer1[30][7:0] = buffer_data_3[2279:2272];
        layer1[30][15:8] = buffer_data_3[2287:2280];
        layer1[30][23:16] = buffer_data_3[2295:2288];
        layer1[30][31:24] = buffer_data_3[2303:2296];
        layer1[30][39:32] = buffer_data_3[2311:2304];
        layer2[30][7:0] = buffer_data_2[2279:2272];
        layer2[30][15:8] = buffer_data_2[2287:2280];
        layer2[30][23:16] = buffer_data_2[2295:2288];
        layer2[30][31:24] = buffer_data_2[2303:2296];
        layer2[30][39:32] = buffer_data_2[2311:2304];
        layer3[30][7:0] = buffer_data_1[2279:2272];
        layer3[30][15:8] = buffer_data_1[2287:2280];
        layer3[30][23:16] = buffer_data_1[2295:2288];
        layer3[30][31:24] = buffer_data_1[2303:2296];
        layer3[30][39:32] = buffer_data_1[2311:2304];
        layer4[30][7:0] = buffer_data_0[2279:2272];
        layer4[30][15:8] = buffer_data_0[2287:2280];
        layer4[30][23:16] = buffer_data_0[2295:2288];
        layer4[30][31:24] = buffer_data_0[2303:2296];
        layer4[30][39:32] = buffer_data_0[2311:2304];
        layer0[31][7:0] = buffer_data_4[2287:2280];
        layer0[31][15:8] = buffer_data_4[2295:2288];
        layer0[31][23:16] = buffer_data_4[2303:2296];
        layer0[31][31:24] = buffer_data_4[2311:2304];
        layer0[31][39:32] = buffer_data_4[2319:2312];
        layer1[31][7:0] = buffer_data_3[2287:2280];
        layer1[31][15:8] = buffer_data_3[2295:2288];
        layer1[31][23:16] = buffer_data_3[2303:2296];
        layer1[31][31:24] = buffer_data_3[2311:2304];
        layer1[31][39:32] = buffer_data_3[2319:2312];
        layer2[31][7:0] = buffer_data_2[2287:2280];
        layer2[31][15:8] = buffer_data_2[2295:2288];
        layer2[31][23:16] = buffer_data_2[2303:2296];
        layer2[31][31:24] = buffer_data_2[2311:2304];
        layer2[31][39:32] = buffer_data_2[2319:2312];
        layer3[31][7:0] = buffer_data_1[2287:2280];
        layer3[31][15:8] = buffer_data_1[2295:2288];
        layer3[31][23:16] = buffer_data_1[2303:2296];
        layer3[31][31:24] = buffer_data_1[2311:2304];
        layer3[31][39:32] = buffer_data_1[2319:2312];
        layer4[31][7:0] = buffer_data_0[2287:2280];
        layer4[31][15:8] = buffer_data_0[2295:2288];
        layer4[31][23:16] = buffer_data_0[2303:2296];
        layer4[31][31:24] = buffer_data_0[2311:2304];
        layer4[31][39:32] = buffer_data_0[2319:2312];
        layer0[32][7:0] = buffer_data_4[2295:2288];
        layer0[32][15:8] = buffer_data_4[2303:2296];
        layer0[32][23:16] = buffer_data_4[2311:2304];
        layer0[32][31:24] = buffer_data_4[2319:2312];
        layer0[32][39:32] = buffer_data_4[2327:2320];
        layer1[32][7:0] = buffer_data_3[2295:2288];
        layer1[32][15:8] = buffer_data_3[2303:2296];
        layer1[32][23:16] = buffer_data_3[2311:2304];
        layer1[32][31:24] = buffer_data_3[2319:2312];
        layer1[32][39:32] = buffer_data_3[2327:2320];
        layer2[32][7:0] = buffer_data_2[2295:2288];
        layer2[32][15:8] = buffer_data_2[2303:2296];
        layer2[32][23:16] = buffer_data_2[2311:2304];
        layer2[32][31:24] = buffer_data_2[2319:2312];
        layer2[32][39:32] = buffer_data_2[2327:2320];
        layer3[32][7:0] = buffer_data_1[2295:2288];
        layer3[32][15:8] = buffer_data_1[2303:2296];
        layer3[32][23:16] = buffer_data_1[2311:2304];
        layer3[32][31:24] = buffer_data_1[2319:2312];
        layer3[32][39:32] = buffer_data_1[2327:2320];
        layer4[32][7:0] = buffer_data_0[2295:2288];
        layer4[32][15:8] = buffer_data_0[2303:2296];
        layer4[32][23:16] = buffer_data_0[2311:2304];
        layer4[32][31:24] = buffer_data_0[2319:2312];
        layer4[32][39:32] = buffer_data_0[2327:2320];
        layer0[33][7:0] = buffer_data_4[2303:2296];
        layer0[33][15:8] = buffer_data_4[2311:2304];
        layer0[33][23:16] = buffer_data_4[2319:2312];
        layer0[33][31:24] = buffer_data_4[2327:2320];
        layer0[33][39:32] = buffer_data_4[2335:2328];
        layer1[33][7:0] = buffer_data_3[2303:2296];
        layer1[33][15:8] = buffer_data_3[2311:2304];
        layer1[33][23:16] = buffer_data_3[2319:2312];
        layer1[33][31:24] = buffer_data_3[2327:2320];
        layer1[33][39:32] = buffer_data_3[2335:2328];
        layer2[33][7:0] = buffer_data_2[2303:2296];
        layer2[33][15:8] = buffer_data_2[2311:2304];
        layer2[33][23:16] = buffer_data_2[2319:2312];
        layer2[33][31:24] = buffer_data_2[2327:2320];
        layer2[33][39:32] = buffer_data_2[2335:2328];
        layer3[33][7:0] = buffer_data_1[2303:2296];
        layer3[33][15:8] = buffer_data_1[2311:2304];
        layer3[33][23:16] = buffer_data_1[2319:2312];
        layer3[33][31:24] = buffer_data_1[2327:2320];
        layer3[33][39:32] = buffer_data_1[2335:2328];
        layer4[33][7:0] = buffer_data_0[2303:2296];
        layer4[33][15:8] = buffer_data_0[2311:2304];
        layer4[33][23:16] = buffer_data_0[2319:2312];
        layer4[33][31:24] = buffer_data_0[2327:2320];
        layer4[33][39:32] = buffer_data_0[2335:2328];
        layer0[34][7:0] = buffer_data_4[2311:2304];
        layer0[34][15:8] = buffer_data_4[2319:2312];
        layer0[34][23:16] = buffer_data_4[2327:2320];
        layer0[34][31:24] = buffer_data_4[2335:2328];
        layer0[34][39:32] = buffer_data_4[2343:2336];
        layer1[34][7:0] = buffer_data_3[2311:2304];
        layer1[34][15:8] = buffer_data_3[2319:2312];
        layer1[34][23:16] = buffer_data_3[2327:2320];
        layer1[34][31:24] = buffer_data_3[2335:2328];
        layer1[34][39:32] = buffer_data_3[2343:2336];
        layer2[34][7:0] = buffer_data_2[2311:2304];
        layer2[34][15:8] = buffer_data_2[2319:2312];
        layer2[34][23:16] = buffer_data_2[2327:2320];
        layer2[34][31:24] = buffer_data_2[2335:2328];
        layer2[34][39:32] = buffer_data_2[2343:2336];
        layer3[34][7:0] = buffer_data_1[2311:2304];
        layer3[34][15:8] = buffer_data_1[2319:2312];
        layer3[34][23:16] = buffer_data_1[2327:2320];
        layer3[34][31:24] = buffer_data_1[2335:2328];
        layer3[34][39:32] = buffer_data_1[2343:2336];
        layer4[34][7:0] = buffer_data_0[2311:2304];
        layer4[34][15:8] = buffer_data_0[2319:2312];
        layer4[34][23:16] = buffer_data_0[2327:2320];
        layer4[34][31:24] = buffer_data_0[2335:2328];
        layer4[34][39:32] = buffer_data_0[2343:2336];
        layer0[35][7:0] = buffer_data_4[2319:2312];
        layer0[35][15:8] = buffer_data_4[2327:2320];
        layer0[35][23:16] = buffer_data_4[2335:2328];
        layer0[35][31:24] = buffer_data_4[2343:2336];
        layer0[35][39:32] = buffer_data_4[2351:2344];
        layer1[35][7:0] = buffer_data_3[2319:2312];
        layer1[35][15:8] = buffer_data_3[2327:2320];
        layer1[35][23:16] = buffer_data_3[2335:2328];
        layer1[35][31:24] = buffer_data_3[2343:2336];
        layer1[35][39:32] = buffer_data_3[2351:2344];
        layer2[35][7:0] = buffer_data_2[2319:2312];
        layer2[35][15:8] = buffer_data_2[2327:2320];
        layer2[35][23:16] = buffer_data_2[2335:2328];
        layer2[35][31:24] = buffer_data_2[2343:2336];
        layer2[35][39:32] = buffer_data_2[2351:2344];
        layer3[35][7:0] = buffer_data_1[2319:2312];
        layer3[35][15:8] = buffer_data_1[2327:2320];
        layer3[35][23:16] = buffer_data_1[2335:2328];
        layer3[35][31:24] = buffer_data_1[2343:2336];
        layer3[35][39:32] = buffer_data_1[2351:2344];
        layer4[35][7:0] = buffer_data_0[2319:2312];
        layer4[35][15:8] = buffer_data_0[2327:2320];
        layer4[35][23:16] = buffer_data_0[2335:2328];
        layer4[35][31:24] = buffer_data_0[2343:2336];
        layer4[35][39:32] = buffer_data_0[2351:2344];
        layer0[36][7:0] = buffer_data_4[2327:2320];
        layer0[36][15:8] = buffer_data_4[2335:2328];
        layer0[36][23:16] = buffer_data_4[2343:2336];
        layer0[36][31:24] = buffer_data_4[2351:2344];
        layer0[36][39:32] = buffer_data_4[2359:2352];
        layer1[36][7:0] = buffer_data_3[2327:2320];
        layer1[36][15:8] = buffer_data_3[2335:2328];
        layer1[36][23:16] = buffer_data_3[2343:2336];
        layer1[36][31:24] = buffer_data_3[2351:2344];
        layer1[36][39:32] = buffer_data_3[2359:2352];
        layer2[36][7:0] = buffer_data_2[2327:2320];
        layer2[36][15:8] = buffer_data_2[2335:2328];
        layer2[36][23:16] = buffer_data_2[2343:2336];
        layer2[36][31:24] = buffer_data_2[2351:2344];
        layer2[36][39:32] = buffer_data_2[2359:2352];
        layer3[36][7:0] = buffer_data_1[2327:2320];
        layer3[36][15:8] = buffer_data_1[2335:2328];
        layer3[36][23:16] = buffer_data_1[2343:2336];
        layer3[36][31:24] = buffer_data_1[2351:2344];
        layer3[36][39:32] = buffer_data_1[2359:2352];
        layer4[36][7:0] = buffer_data_0[2327:2320];
        layer4[36][15:8] = buffer_data_0[2335:2328];
        layer4[36][23:16] = buffer_data_0[2343:2336];
        layer4[36][31:24] = buffer_data_0[2351:2344];
        layer4[36][39:32] = buffer_data_0[2359:2352];
        layer0[37][7:0] = buffer_data_4[2335:2328];
        layer0[37][15:8] = buffer_data_4[2343:2336];
        layer0[37][23:16] = buffer_data_4[2351:2344];
        layer0[37][31:24] = buffer_data_4[2359:2352];
        layer0[37][39:32] = buffer_data_4[2367:2360];
        layer1[37][7:0] = buffer_data_3[2335:2328];
        layer1[37][15:8] = buffer_data_3[2343:2336];
        layer1[37][23:16] = buffer_data_3[2351:2344];
        layer1[37][31:24] = buffer_data_3[2359:2352];
        layer1[37][39:32] = buffer_data_3[2367:2360];
        layer2[37][7:0] = buffer_data_2[2335:2328];
        layer2[37][15:8] = buffer_data_2[2343:2336];
        layer2[37][23:16] = buffer_data_2[2351:2344];
        layer2[37][31:24] = buffer_data_2[2359:2352];
        layer2[37][39:32] = buffer_data_2[2367:2360];
        layer3[37][7:0] = buffer_data_1[2335:2328];
        layer3[37][15:8] = buffer_data_1[2343:2336];
        layer3[37][23:16] = buffer_data_1[2351:2344];
        layer3[37][31:24] = buffer_data_1[2359:2352];
        layer3[37][39:32] = buffer_data_1[2367:2360];
        layer4[37][7:0] = buffer_data_0[2335:2328];
        layer4[37][15:8] = buffer_data_0[2343:2336];
        layer4[37][23:16] = buffer_data_0[2351:2344];
        layer4[37][31:24] = buffer_data_0[2359:2352];
        layer4[37][39:32] = buffer_data_0[2367:2360];
        layer0[38][7:0] = buffer_data_4[2343:2336];
        layer0[38][15:8] = buffer_data_4[2351:2344];
        layer0[38][23:16] = buffer_data_4[2359:2352];
        layer0[38][31:24] = buffer_data_4[2367:2360];
        layer0[38][39:32] = buffer_data_4[2375:2368];
        layer1[38][7:0] = buffer_data_3[2343:2336];
        layer1[38][15:8] = buffer_data_3[2351:2344];
        layer1[38][23:16] = buffer_data_3[2359:2352];
        layer1[38][31:24] = buffer_data_3[2367:2360];
        layer1[38][39:32] = buffer_data_3[2375:2368];
        layer2[38][7:0] = buffer_data_2[2343:2336];
        layer2[38][15:8] = buffer_data_2[2351:2344];
        layer2[38][23:16] = buffer_data_2[2359:2352];
        layer2[38][31:24] = buffer_data_2[2367:2360];
        layer2[38][39:32] = buffer_data_2[2375:2368];
        layer3[38][7:0] = buffer_data_1[2343:2336];
        layer3[38][15:8] = buffer_data_1[2351:2344];
        layer3[38][23:16] = buffer_data_1[2359:2352];
        layer3[38][31:24] = buffer_data_1[2367:2360];
        layer3[38][39:32] = buffer_data_1[2375:2368];
        layer4[38][7:0] = buffer_data_0[2343:2336];
        layer4[38][15:8] = buffer_data_0[2351:2344];
        layer4[38][23:16] = buffer_data_0[2359:2352];
        layer4[38][31:24] = buffer_data_0[2367:2360];
        layer4[38][39:32] = buffer_data_0[2375:2368];
        layer0[39][7:0] = buffer_data_4[2351:2344];
        layer0[39][15:8] = buffer_data_4[2359:2352];
        layer0[39][23:16] = buffer_data_4[2367:2360];
        layer0[39][31:24] = buffer_data_4[2375:2368];
        layer0[39][39:32] = buffer_data_4[2383:2376];
        layer1[39][7:0] = buffer_data_3[2351:2344];
        layer1[39][15:8] = buffer_data_3[2359:2352];
        layer1[39][23:16] = buffer_data_3[2367:2360];
        layer1[39][31:24] = buffer_data_3[2375:2368];
        layer1[39][39:32] = buffer_data_3[2383:2376];
        layer2[39][7:0] = buffer_data_2[2351:2344];
        layer2[39][15:8] = buffer_data_2[2359:2352];
        layer2[39][23:16] = buffer_data_2[2367:2360];
        layer2[39][31:24] = buffer_data_2[2375:2368];
        layer2[39][39:32] = buffer_data_2[2383:2376];
        layer3[39][7:0] = buffer_data_1[2351:2344];
        layer3[39][15:8] = buffer_data_1[2359:2352];
        layer3[39][23:16] = buffer_data_1[2367:2360];
        layer3[39][31:24] = buffer_data_1[2375:2368];
        layer3[39][39:32] = buffer_data_1[2383:2376];
        layer4[39][7:0] = buffer_data_0[2351:2344];
        layer4[39][15:8] = buffer_data_0[2359:2352];
        layer4[39][23:16] = buffer_data_0[2367:2360];
        layer4[39][31:24] = buffer_data_0[2375:2368];
        layer4[39][39:32] = buffer_data_0[2383:2376];
        layer0[40][7:0] = buffer_data_4[2359:2352];
        layer0[40][15:8] = buffer_data_4[2367:2360];
        layer0[40][23:16] = buffer_data_4[2375:2368];
        layer0[40][31:24] = buffer_data_4[2383:2376];
        layer0[40][39:32] = buffer_data_4[2391:2384];
        layer1[40][7:0] = buffer_data_3[2359:2352];
        layer1[40][15:8] = buffer_data_3[2367:2360];
        layer1[40][23:16] = buffer_data_3[2375:2368];
        layer1[40][31:24] = buffer_data_3[2383:2376];
        layer1[40][39:32] = buffer_data_3[2391:2384];
        layer2[40][7:0] = buffer_data_2[2359:2352];
        layer2[40][15:8] = buffer_data_2[2367:2360];
        layer2[40][23:16] = buffer_data_2[2375:2368];
        layer2[40][31:24] = buffer_data_2[2383:2376];
        layer2[40][39:32] = buffer_data_2[2391:2384];
        layer3[40][7:0] = buffer_data_1[2359:2352];
        layer3[40][15:8] = buffer_data_1[2367:2360];
        layer3[40][23:16] = buffer_data_1[2375:2368];
        layer3[40][31:24] = buffer_data_1[2383:2376];
        layer3[40][39:32] = buffer_data_1[2391:2384];
        layer4[40][7:0] = buffer_data_0[2359:2352];
        layer4[40][15:8] = buffer_data_0[2367:2360];
        layer4[40][23:16] = buffer_data_0[2375:2368];
        layer4[40][31:24] = buffer_data_0[2383:2376];
        layer4[40][39:32] = buffer_data_0[2391:2384];
        layer0[41][7:0] = buffer_data_4[2367:2360];
        layer0[41][15:8] = buffer_data_4[2375:2368];
        layer0[41][23:16] = buffer_data_4[2383:2376];
        layer0[41][31:24] = buffer_data_4[2391:2384];
        layer0[41][39:32] = buffer_data_4[2399:2392];
        layer1[41][7:0] = buffer_data_3[2367:2360];
        layer1[41][15:8] = buffer_data_3[2375:2368];
        layer1[41][23:16] = buffer_data_3[2383:2376];
        layer1[41][31:24] = buffer_data_3[2391:2384];
        layer1[41][39:32] = buffer_data_3[2399:2392];
        layer2[41][7:0] = buffer_data_2[2367:2360];
        layer2[41][15:8] = buffer_data_2[2375:2368];
        layer2[41][23:16] = buffer_data_2[2383:2376];
        layer2[41][31:24] = buffer_data_2[2391:2384];
        layer2[41][39:32] = buffer_data_2[2399:2392];
        layer3[41][7:0] = buffer_data_1[2367:2360];
        layer3[41][15:8] = buffer_data_1[2375:2368];
        layer3[41][23:16] = buffer_data_1[2383:2376];
        layer3[41][31:24] = buffer_data_1[2391:2384];
        layer3[41][39:32] = buffer_data_1[2399:2392];
        layer4[41][7:0] = buffer_data_0[2367:2360];
        layer4[41][15:8] = buffer_data_0[2375:2368];
        layer4[41][23:16] = buffer_data_0[2383:2376];
        layer4[41][31:24] = buffer_data_0[2391:2384];
        layer4[41][39:32] = buffer_data_0[2399:2392];
        layer0[42][7:0] = buffer_data_4[2375:2368];
        layer0[42][15:8] = buffer_data_4[2383:2376];
        layer0[42][23:16] = buffer_data_4[2391:2384];
        layer0[42][31:24] = buffer_data_4[2399:2392];
        layer0[42][39:32] = buffer_data_4[2407:2400];
        layer1[42][7:0] = buffer_data_3[2375:2368];
        layer1[42][15:8] = buffer_data_3[2383:2376];
        layer1[42][23:16] = buffer_data_3[2391:2384];
        layer1[42][31:24] = buffer_data_3[2399:2392];
        layer1[42][39:32] = buffer_data_3[2407:2400];
        layer2[42][7:0] = buffer_data_2[2375:2368];
        layer2[42][15:8] = buffer_data_2[2383:2376];
        layer2[42][23:16] = buffer_data_2[2391:2384];
        layer2[42][31:24] = buffer_data_2[2399:2392];
        layer2[42][39:32] = buffer_data_2[2407:2400];
        layer3[42][7:0] = buffer_data_1[2375:2368];
        layer3[42][15:8] = buffer_data_1[2383:2376];
        layer3[42][23:16] = buffer_data_1[2391:2384];
        layer3[42][31:24] = buffer_data_1[2399:2392];
        layer3[42][39:32] = buffer_data_1[2407:2400];
        layer4[42][7:0] = buffer_data_0[2375:2368];
        layer4[42][15:8] = buffer_data_0[2383:2376];
        layer4[42][23:16] = buffer_data_0[2391:2384];
        layer4[42][31:24] = buffer_data_0[2399:2392];
        layer4[42][39:32] = buffer_data_0[2407:2400];
        layer0[43][7:0] = buffer_data_4[2383:2376];
        layer0[43][15:8] = buffer_data_4[2391:2384];
        layer0[43][23:16] = buffer_data_4[2399:2392];
        layer0[43][31:24] = buffer_data_4[2407:2400];
        layer0[43][39:32] = buffer_data_4[2415:2408];
        layer1[43][7:0] = buffer_data_3[2383:2376];
        layer1[43][15:8] = buffer_data_3[2391:2384];
        layer1[43][23:16] = buffer_data_3[2399:2392];
        layer1[43][31:24] = buffer_data_3[2407:2400];
        layer1[43][39:32] = buffer_data_3[2415:2408];
        layer2[43][7:0] = buffer_data_2[2383:2376];
        layer2[43][15:8] = buffer_data_2[2391:2384];
        layer2[43][23:16] = buffer_data_2[2399:2392];
        layer2[43][31:24] = buffer_data_2[2407:2400];
        layer2[43][39:32] = buffer_data_2[2415:2408];
        layer3[43][7:0] = buffer_data_1[2383:2376];
        layer3[43][15:8] = buffer_data_1[2391:2384];
        layer3[43][23:16] = buffer_data_1[2399:2392];
        layer3[43][31:24] = buffer_data_1[2407:2400];
        layer3[43][39:32] = buffer_data_1[2415:2408];
        layer4[43][7:0] = buffer_data_0[2383:2376];
        layer4[43][15:8] = buffer_data_0[2391:2384];
        layer4[43][23:16] = buffer_data_0[2399:2392];
        layer4[43][31:24] = buffer_data_0[2407:2400];
        layer4[43][39:32] = buffer_data_0[2415:2408];
        layer0[44][7:0] = buffer_data_4[2391:2384];
        layer0[44][15:8] = buffer_data_4[2399:2392];
        layer0[44][23:16] = buffer_data_4[2407:2400];
        layer0[44][31:24] = buffer_data_4[2415:2408];
        layer0[44][39:32] = buffer_data_4[2423:2416];
        layer1[44][7:0] = buffer_data_3[2391:2384];
        layer1[44][15:8] = buffer_data_3[2399:2392];
        layer1[44][23:16] = buffer_data_3[2407:2400];
        layer1[44][31:24] = buffer_data_3[2415:2408];
        layer1[44][39:32] = buffer_data_3[2423:2416];
        layer2[44][7:0] = buffer_data_2[2391:2384];
        layer2[44][15:8] = buffer_data_2[2399:2392];
        layer2[44][23:16] = buffer_data_2[2407:2400];
        layer2[44][31:24] = buffer_data_2[2415:2408];
        layer2[44][39:32] = buffer_data_2[2423:2416];
        layer3[44][7:0] = buffer_data_1[2391:2384];
        layer3[44][15:8] = buffer_data_1[2399:2392];
        layer3[44][23:16] = buffer_data_1[2407:2400];
        layer3[44][31:24] = buffer_data_1[2415:2408];
        layer3[44][39:32] = buffer_data_1[2423:2416];
        layer4[44][7:0] = buffer_data_0[2391:2384];
        layer4[44][15:8] = buffer_data_0[2399:2392];
        layer4[44][23:16] = buffer_data_0[2407:2400];
        layer4[44][31:24] = buffer_data_0[2415:2408];
        layer4[44][39:32] = buffer_data_0[2423:2416];
        layer0[45][7:0] = buffer_data_4[2399:2392];
        layer0[45][15:8] = buffer_data_4[2407:2400];
        layer0[45][23:16] = buffer_data_4[2415:2408];
        layer0[45][31:24] = buffer_data_4[2423:2416];
        layer0[45][39:32] = buffer_data_4[2431:2424];
        layer1[45][7:0] = buffer_data_3[2399:2392];
        layer1[45][15:8] = buffer_data_3[2407:2400];
        layer1[45][23:16] = buffer_data_3[2415:2408];
        layer1[45][31:24] = buffer_data_3[2423:2416];
        layer1[45][39:32] = buffer_data_3[2431:2424];
        layer2[45][7:0] = buffer_data_2[2399:2392];
        layer2[45][15:8] = buffer_data_2[2407:2400];
        layer2[45][23:16] = buffer_data_2[2415:2408];
        layer2[45][31:24] = buffer_data_2[2423:2416];
        layer2[45][39:32] = buffer_data_2[2431:2424];
        layer3[45][7:0] = buffer_data_1[2399:2392];
        layer3[45][15:8] = buffer_data_1[2407:2400];
        layer3[45][23:16] = buffer_data_1[2415:2408];
        layer3[45][31:24] = buffer_data_1[2423:2416];
        layer3[45][39:32] = buffer_data_1[2431:2424];
        layer4[45][7:0] = buffer_data_0[2399:2392];
        layer4[45][15:8] = buffer_data_0[2407:2400];
        layer4[45][23:16] = buffer_data_0[2415:2408];
        layer4[45][31:24] = buffer_data_0[2423:2416];
        layer4[45][39:32] = buffer_data_0[2431:2424];
        layer0[46][7:0] = buffer_data_4[2407:2400];
        layer0[46][15:8] = buffer_data_4[2415:2408];
        layer0[46][23:16] = buffer_data_4[2423:2416];
        layer0[46][31:24] = buffer_data_4[2431:2424];
        layer0[46][39:32] = buffer_data_4[2439:2432];
        layer1[46][7:0] = buffer_data_3[2407:2400];
        layer1[46][15:8] = buffer_data_3[2415:2408];
        layer1[46][23:16] = buffer_data_3[2423:2416];
        layer1[46][31:24] = buffer_data_3[2431:2424];
        layer1[46][39:32] = buffer_data_3[2439:2432];
        layer2[46][7:0] = buffer_data_2[2407:2400];
        layer2[46][15:8] = buffer_data_2[2415:2408];
        layer2[46][23:16] = buffer_data_2[2423:2416];
        layer2[46][31:24] = buffer_data_2[2431:2424];
        layer2[46][39:32] = buffer_data_2[2439:2432];
        layer3[46][7:0] = buffer_data_1[2407:2400];
        layer3[46][15:8] = buffer_data_1[2415:2408];
        layer3[46][23:16] = buffer_data_1[2423:2416];
        layer3[46][31:24] = buffer_data_1[2431:2424];
        layer3[46][39:32] = buffer_data_1[2439:2432];
        layer4[46][7:0] = buffer_data_0[2407:2400];
        layer4[46][15:8] = buffer_data_0[2415:2408];
        layer4[46][23:16] = buffer_data_0[2423:2416];
        layer4[46][31:24] = buffer_data_0[2431:2424];
        layer4[46][39:32] = buffer_data_0[2439:2432];
        layer0[47][7:0] = buffer_data_4[2415:2408];
        layer0[47][15:8] = buffer_data_4[2423:2416];
        layer0[47][23:16] = buffer_data_4[2431:2424];
        layer0[47][31:24] = buffer_data_4[2439:2432];
        layer0[47][39:32] = buffer_data_4[2447:2440];
        layer1[47][7:0] = buffer_data_3[2415:2408];
        layer1[47][15:8] = buffer_data_3[2423:2416];
        layer1[47][23:16] = buffer_data_3[2431:2424];
        layer1[47][31:24] = buffer_data_3[2439:2432];
        layer1[47][39:32] = buffer_data_3[2447:2440];
        layer2[47][7:0] = buffer_data_2[2415:2408];
        layer2[47][15:8] = buffer_data_2[2423:2416];
        layer2[47][23:16] = buffer_data_2[2431:2424];
        layer2[47][31:24] = buffer_data_2[2439:2432];
        layer2[47][39:32] = buffer_data_2[2447:2440];
        layer3[47][7:0] = buffer_data_1[2415:2408];
        layer3[47][15:8] = buffer_data_1[2423:2416];
        layer3[47][23:16] = buffer_data_1[2431:2424];
        layer3[47][31:24] = buffer_data_1[2439:2432];
        layer3[47][39:32] = buffer_data_1[2447:2440];
        layer4[47][7:0] = buffer_data_0[2415:2408];
        layer4[47][15:8] = buffer_data_0[2423:2416];
        layer4[47][23:16] = buffer_data_0[2431:2424];
        layer4[47][31:24] = buffer_data_0[2439:2432];
        layer4[47][39:32] = buffer_data_0[2447:2440];
        layer0[48][7:0] = buffer_data_4[2423:2416];
        layer0[48][15:8] = buffer_data_4[2431:2424];
        layer0[48][23:16] = buffer_data_4[2439:2432];
        layer0[48][31:24] = buffer_data_4[2447:2440];
        layer0[48][39:32] = buffer_data_4[2455:2448];
        layer1[48][7:0] = buffer_data_3[2423:2416];
        layer1[48][15:8] = buffer_data_3[2431:2424];
        layer1[48][23:16] = buffer_data_3[2439:2432];
        layer1[48][31:24] = buffer_data_3[2447:2440];
        layer1[48][39:32] = buffer_data_3[2455:2448];
        layer2[48][7:0] = buffer_data_2[2423:2416];
        layer2[48][15:8] = buffer_data_2[2431:2424];
        layer2[48][23:16] = buffer_data_2[2439:2432];
        layer2[48][31:24] = buffer_data_2[2447:2440];
        layer2[48][39:32] = buffer_data_2[2455:2448];
        layer3[48][7:0] = buffer_data_1[2423:2416];
        layer3[48][15:8] = buffer_data_1[2431:2424];
        layer3[48][23:16] = buffer_data_1[2439:2432];
        layer3[48][31:24] = buffer_data_1[2447:2440];
        layer3[48][39:32] = buffer_data_1[2455:2448];
        layer4[48][7:0] = buffer_data_0[2423:2416];
        layer4[48][15:8] = buffer_data_0[2431:2424];
        layer4[48][23:16] = buffer_data_0[2439:2432];
        layer4[48][31:24] = buffer_data_0[2447:2440];
        layer4[48][39:32] = buffer_data_0[2455:2448];
        layer0[49][7:0] = buffer_data_4[2431:2424];
        layer0[49][15:8] = buffer_data_4[2439:2432];
        layer0[49][23:16] = buffer_data_4[2447:2440];
        layer0[49][31:24] = buffer_data_4[2455:2448];
        layer0[49][39:32] = buffer_data_4[2463:2456];
        layer1[49][7:0] = buffer_data_3[2431:2424];
        layer1[49][15:8] = buffer_data_3[2439:2432];
        layer1[49][23:16] = buffer_data_3[2447:2440];
        layer1[49][31:24] = buffer_data_3[2455:2448];
        layer1[49][39:32] = buffer_data_3[2463:2456];
        layer2[49][7:0] = buffer_data_2[2431:2424];
        layer2[49][15:8] = buffer_data_2[2439:2432];
        layer2[49][23:16] = buffer_data_2[2447:2440];
        layer2[49][31:24] = buffer_data_2[2455:2448];
        layer2[49][39:32] = buffer_data_2[2463:2456];
        layer3[49][7:0] = buffer_data_1[2431:2424];
        layer3[49][15:8] = buffer_data_1[2439:2432];
        layer3[49][23:16] = buffer_data_1[2447:2440];
        layer3[49][31:24] = buffer_data_1[2455:2448];
        layer3[49][39:32] = buffer_data_1[2463:2456];
        layer4[49][7:0] = buffer_data_0[2431:2424];
        layer4[49][15:8] = buffer_data_0[2439:2432];
        layer4[49][23:16] = buffer_data_0[2447:2440];
        layer4[49][31:24] = buffer_data_0[2455:2448];
        layer4[49][39:32] = buffer_data_0[2463:2456];
        layer0[50][7:0] = buffer_data_4[2439:2432];
        layer0[50][15:8] = buffer_data_4[2447:2440];
        layer0[50][23:16] = buffer_data_4[2455:2448];
        layer0[50][31:24] = buffer_data_4[2463:2456];
        layer0[50][39:32] = buffer_data_4[2471:2464];
        layer1[50][7:0] = buffer_data_3[2439:2432];
        layer1[50][15:8] = buffer_data_3[2447:2440];
        layer1[50][23:16] = buffer_data_3[2455:2448];
        layer1[50][31:24] = buffer_data_3[2463:2456];
        layer1[50][39:32] = buffer_data_3[2471:2464];
        layer2[50][7:0] = buffer_data_2[2439:2432];
        layer2[50][15:8] = buffer_data_2[2447:2440];
        layer2[50][23:16] = buffer_data_2[2455:2448];
        layer2[50][31:24] = buffer_data_2[2463:2456];
        layer2[50][39:32] = buffer_data_2[2471:2464];
        layer3[50][7:0] = buffer_data_1[2439:2432];
        layer3[50][15:8] = buffer_data_1[2447:2440];
        layer3[50][23:16] = buffer_data_1[2455:2448];
        layer3[50][31:24] = buffer_data_1[2463:2456];
        layer3[50][39:32] = buffer_data_1[2471:2464];
        layer4[50][7:0] = buffer_data_0[2439:2432];
        layer4[50][15:8] = buffer_data_0[2447:2440];
        layer4[50][23:16] = buffer_data_0[2455:2448];
        layer4[50][31:24] = buffer_data_0[2463:2456];
        layer4[50][39:32] = buffer_data_0[2471:2464];
        layer0[51][7:0] = buffer_data_4[2447:2440];
        layer0[51][15:8] = buffer_data_4[2455:2448];
        layer0[51][23:16] = buffer_data_4[2463:2456];
        layer0[51][31:24] = buffer_data_4[2471:2464];
        layer0[51][39:32] = buffer_data_4[2479:2472];
        layer1[51][7:0] = buffer_data_3[2447:2440];
        layer1[51][15:8] = buffer_data_3[2455:2448];
        layer1[51][23:16] = buffer_data_3[2463:2456];
        layer1[51][31:24] = buffer_data_3[2471:2464];
        layer1[51][39:32] = buffer_data_3[2479:2472];
        layer2[51][7:0] = buffer_data_2[2447:2440];
        layer2[51][15:8] = buffer_data_2[2455:2448];
        layer2[51][23:16] = buffer_data_2[2463:2456];
        layer2[51][31:24] = buffer_data_2[2471:2464];
        layer2[51][39:32] = buffer_data_2[2479:2472];
        layer3[51][7:0] = buffer_data_1[2447:2440];
        layer3[51][15:8] = buffer_data_1[2455:2448];
        layer3[51][23:16] = buffer_data_1[2463:2456];
        layer3[51][31:24] = buffer_data_1[2471:2464];
        layer3[51][39:32] = buffer_data_1[2479:2472];
        layer4[51][7:0] = buffer_data_0[2447:2440];
        layer4[51][15:8] = buffer_data_0[2455:2448];
        layer4[51][23:16] = buffer_data_0[2463:2456];
        layer4[51][31:24] = buffer_data_0[2471:2464];
        layer4[51][39:32] = buffer_data_0[2479:2472];
        layer0[52][7:0] = buffer_data_4[2455:2448];
        layer0[52][15:8] = buffer_data_4[2463:2456];
        layer0[52][23:16] = buffer_data_4[2471:2464];
        layer0[52][31:24] = buffer_data_4[2479:2472];
        layer0[52][39:32] = buffer_data_4[2487:2480];
        layer1[52][7:0] = buffer_data_3[2455:2448];
        layer1[52][15:8] = buffer_data_3[2463:2456];
        layer1[52][23:16] = buffer_data_3[2471:2464];
        layer1[52][31:24] = buffer_data_3[2479:2472];
        layer1[52][39:32] = buffer_data_3[2487:2480];
        layer2[52][7:0] = buffer_data_2[2455:2448];
        layer2[52][15:8] = buffer_data_2[2463:2456];
        layer2[52][23:16] = buffer_data_2[2471:2464];
        layer2[52][31:24] = buffer_data_2[2479:2472];
        layer2[52][39:32] = buffer_data_2[2487:2480];
        layer3[52][7:0] = buffer_data_1[2455:2448];
        layer3[52][15:8] = buffer_data_1[2463:2456];
        layer3[52][23:16] = buffer_data_1[2471:2464];
        layer3[52][31:24] = buffer_data_1[2479:2472];
        layer3[52][39:32] = buffer_data_1[2487:2480];
        layer4[52][7:0] = buffer_data_0[2455:2448];
        layer4[52][15:8] = buffer_data_0[2463:2456];
        layer4[52][23:16] = buffer_data_0[2471:2464];
        layer4[52][31:24] = buffer_data_0[2479:2472];
        layer4[52][39:32] = buffer_data_0[2487:2480];
        layer0[53][7:0] = buffer_data_4[2463:2456];
        layer0[53][15:8] = buffer_data_4[2471:2464];
        layer0[53][23:16] = buffer_data_4[2479:2472];
        layer0[53][31:24] = buffer_data_4[2487:2480];
        layer0[53][39:32] = buffer_data_4[2495:2488];
        layer1[53][7:0] = buffer_data_3[2463:2456];
        layer1[53][15:8] = buffer_data_3[2471:2464];
        layer1[53][23:16] = buffer_data_3[2479:2472];
        layer1[53][31:24] = buffer_data_3[2487:2480];
        layer1[53][39:32] = buffer_data_3[2495:2488];
        layer2[53][7:0] = buffer_data_2[2463:2456];
        layer2[53][15:8] = buffer_data_2[2471:2464];
        layer2[53][23:16] = buffer_data_2[2479:2472];
        layer2[53][31:24] = buffer_data_2[2487:2480];
        layer2[53][39:32] = buffer_data_2[2495:2488];
        layer3[53][7:0] = buffer_data_1[2463:2456];
        layer3[53][15:8] = buffer_data_1[2471:2464];
        layer3[53][23:16] = buffer_data_1[2479:2472];
        layer3[53][31:24] = buffer_data_1[2487:2480];
        layer3[53][39:32] = buffer_data_1[2495:2488];
        layer4[53][7:0] = buffer_data_0[2463:2456];
        layer4[53][15:8] = buffer_data_0[2471:2464];
        layer4[53][23:16] = buffer_data_0[2479:2472];
        layer4[53][31:24] = buffer_data_0[2487:2480];
        layer4[53][39:32] = buffer_data_0[2495:2488];
        layer0[54][7:0] = buffer_data_4[2471:2464];
        layer0[54][15:8] = buffer_data_4[2479:2472];
        layer0[54][23:16] = buffer_data_4[2487:2480];
        layer0[54][31:24] = buffer_data_4[2495:2488];
        layer0[54][39:32] = buffer_data_4[2503:2496];
        layer1[54][7:0] = buffer_data_3[2471:2464];
        layer1[54][15:8] = buffer_data_3[2479:2472];
        layer1[54][23:16] = buffer_data_3[2487:2480];
        layer1[54][31:24] = buffer_data_3[2495:2488];
        layer1[54][39:32] = buffer_data_3[2503:2496];
        layer2[54][7:0] = buffer_data_2[2471:2464];
        layer2[54][15:8] = buffer_data_2[2479:2472];
        layer2[54][23:16] = buffer_data_2[2487:2480];
        layer2[54][31:24] = buffer_data_2[2495:2488];
        layer2[54][39:32] = buffer_data_2[2503:2496];
        layer3[54][7:0] = buffer_data_1[2471:2464];
        layer3[54][15:8] = buffer_data_1[2479:2472];
        layer3[54][23:16] = buffer_data_1[2487:2480];
        layer3[54][31:24] = buffer_data_1[2495:2488];
        layer3[54][39:32] = buffer_data_1[2503:2496];
        layer4[54][7:0] = buffer_data_0[2471:2464];
        layer4[54][15:8] = buffer_data_0[2479:2472];
        layer4[54][23:16] = buffer_data_0[2487:2480];
        layer4[54][31:24] = buffer_data_0[2495:2488];
        layer4[54][39:32] = buffer_data_0[2503:2496];
        layer0[55][7:0] = buffer_data_4[2479:2472];
        layer0[55][15:8] = buffer_data_4[2487:2480];
        layer0[55][23:16] = buffer_data_4[2495:2488];
        layer0[55][31:24] = buffer_data_4[2503:2496];
        layer0[55][39:32] = buffer_data_4[2511:2504];
        layer1[55][7:0] = buffer_data_3[2479:2472];
        layer1[55][15:8] = buffer_data_3[2487:2480];
        layer1[55][23:16] = buffer_data_3[2495:2488];
        layer1[55][31:24] = buffer_data_3[2503:2496];
        layer1[55][39:32] = buffer_data_3[2511:2504];
        layer2[55][7:0] = buffer_data_2[2479:2472];
        layer2[55][15:8] = buffer_data_2[2487:2480];
        layer2[55][23:16] = buffer_data_2[2495:2488];
        layer2[55][31:24] = buffer_data_2[2503:2496];
        layer2[55][39:32] = buffer_data_2[2511:2504];
        layer3[55][7:0] = buffer_data_1[2479:2472];
        layer3[55][15:8] = buffer_data_1[2487:2480];
        layer3[55][23:16] = buffer_data_1[2495:2488];
        layer3[55][31:24] = buffer_data_1[2503:2496];
        layer3[55][39:32] = buffer_data_1[2511:2504];
        layer4[55][7:0] = buffer_data_0[2479:2472];
        layer4[55][15:8] = buffer_data_0[2487:2480];
        layer4[55][23:16] = buffer_data_0[2495:2488];
        layer4[55][31:24] = buffer_data_0[2503:2496];
        layer4[55][39:32] = buffer_data_0[2511:2504];
        layer0[56][7:0] = buffer_data_4[2487:2480];
        layer0[56][15:8] = buffer_data_4[2495:2488];
        layer0[56][23:16] = buffer_data_4[2503:2496];
        layer0[56][31:24] = buffer_data_4[2511:2504];
        layer0[56][39:32] = buffer_data_4[2519:2512];
        layer1[56][7:0] = buffer_data_3[2487:2480];
        layer1[56][15:8] = buffer_data_3[2495:2488];
        layer1[56][23:16] = buffer_data_3[2503:2496];
        layer1[56][31:24] = buffer_data_3[2511:2504];
        layer1[56][39:32] = buffer_data_3[2519:2512];
        layer2[56][7:0] = buffer_data_2[2487:2480];
        layer2[56][15:8] = buffer_data_2[2495:2488];
        layer2[56][23:16] = buffer_data_2[2503:2496];
        layer2[56][31:24] = buffer_data_2[2511:2504];
        layer2[56][39:32] = buffer_data_2[2519:2512];
        layer3[56][7:0] = buffer_data_1[2487:2480];
        layer3[56][15:8] = buffer_data_1[2495:2488];
        layer3[56][23:16] = buffer_data_1[2503:2496];
        layer3[56][31:24] = buffer_data_1[2511:2504];
        layer3[56][39:32] = buffer_data_1[2519:2512];
        layer4[56][7:0] = buffer_data_0[2487:2480];
        layer4[56][15:8] = buffer_data_0[2495:2488];
        layer4[56][23:16] = buffer_data_0[2503:2496];
        layer4[56][31:24] = buffer_data_0[2511:2504];
        layer4[56][39:32] = buffer_data_0[2519:2512];
        layer0[57][7:0] = buffer_data_4[2495:2488];
        layer0[57][15:8] = buffer_data_4[2503:2496];
        layer0[57][23:16] = buffer_data_4[2511:2504];
        layer0[57][31:24] = buffer_data_4[2519:2512];
        layer0[57][39:32] = buffer_data_4[2527:2520];
        layer1[57][7:0] = buffer_data_3[2495:2488];
        layer1[57][15:8] = buffer_data_3[2503:2496];
        layer1[57][23:16] = buffer_data_3[2511:2504];
        layer1[57][31:24] = buffer_data_3[2519:2512];
        layer1[57][39:32] = buffer_data_3[2527:2520];
        layer2[57][7:0] = buffer_data_2[2495:2488];
        layer2[57][15:8] = buffer_data_2[2503:2496];
        layer2[57][23:16] = buffer_data_2[2511:2504];
        layer2[57][31:24] = buffer_data_2[2519:2512];
        layer2[57][39:32] = buffer_data_2[2527:2520];
        layer3[57][7:0] = buffer_data_1[2495:2488];
        layer3[57][15:8] = buffer_data_1[2503:2496];
        layer3[57][23:16] = buffer_data_1[2511:2504];
        layer3[57][31:24] = buffer_data_1[2519:2512];
        layer3[57][39:32] = buffer_data_1[2527:2520];
        layer4[57][7:0] = buffer_data_0[2495:2488];
        layer4[57][15:8] = buffer_data_0[2503:2496];
        layer4[57][23:16] = buffer_data_0[2511:2504];
        layer4[57][31:24] = buffer_data_0[2519:2512];
        layer4[57][39:32] = buffer_data_0[2527:2520];
        layer0[58][7:0] = buffer_data_4[2503:2496];
        layer0[58][15:8] = buffer_data_4[2511:2504];
        layer0[58][23:16] = buffer_data_4[2519:2512];
        layer0[58][31:24] = buffer_data_4[2527:2520];
        layer0[58][39:32] = buffer_data_4[2535:2528];
        layer1[58][7:0] = buffer_data_3[2503:2496];
        layer1[58][15:8] = buffer_data_3[2511:2504];
        layer1[58][23:16] = buffer_data_3[2519:2512];
        layer1[58][31:24] = buffer_data_3[2527:2520];
        layer1[58][39:32] = buffer_data_3[2535:2528];
        layer2[58][7:0] = buffer_data_2[2503:2496];
        layer2[58][15:8] = buffer_data_2[2511:2504];
        layer2[58][23:16] = buffer_data_2[2519:2512];
        layer2[58][31:24] = buffer_data_2[2527:2520];
        layer2[58][39:32] = buffer_data_2[2535:2528];
        layer3[58][7:0] = buffer_data_1[2503:2496];
        layer3[58][15:8] = buffer_data_1[2511:2504];
        layer3[58][23:16] = buffer_data_1[2519:2512];
        layer3[58][31:24] = buffer_data_1[2527:2520];
        layer3[58][39:32] = buffer_data_1[2535:2528];
        layer4[58][7:0] = buffer_data_0[2503:2496];
        layer4[58][15:8] = buffer_data_0[2511:2504];
        layer4[58][23:16] = buffer_data_0[2519:2512];
        layer4[58][31:24] = buffer_data_0[2527:2520];
        layer4[58][39:32] = buffer_data_0[2535:2528];
        layer0[59][7:0] = buffer_data_4[2511:2504];
        layer0[59][15:8] = buffer_data_4[2519:2512];
        layer0[59][23:16] = buffer_data_4[2527:2520];
        layer0[59][31:24] = buffer_data_4[2535:2528];
        layer0[59][39:32] = buffer_data_4[2543:2536];
        layer1[59][7:0] = buffer_data_3[2511:2504];
        layer1[59][15:8] = buffer_data_3[2519:2512];
        layer1[59][23:16] = buffer_data_3[2527:2520];
        layer1[59][31:24] = buffer_data_3[2535:2528];
        layer1[59][39:32] = buffer_data_3[2543:2536];
        layer2[59][7:0] = buffer_data_2[2511:2504];
        layer2[59][15:8] = buffer_data_2[2519:2512];
        layer2[59][23:16] = buffer_data_2[2527:2520];
        layer2[59][31:24] = buffer_data_2[2535:2528];
        layer2[59][39:32] = buffer_data_2[2543:2536];
        layer3[59][7:0] = buffer_data_1[2511:2504];
        layer3[59][15:8] = buffer_data_1[2519:2512];
        layer3[59][23:16] = buffer_data_1[2527:2520];
        layer3[59][31:24] = buffer_data_1[2535:2528];
        layer3[59][39:32] = buffer_data_1[2543:2536];
        layer4[59][7:0] = buffer_data_0[2511:2504];
        layer4[59][15:8] = buffer_data_0[2519:2512];
        layer4[59][23:16] = buffer_data_0[2527:2520];
        layer4[59][31:24] = buffer_data_0[2535:2528];
        layer4[59][39:32] = buffer_data_0[2543:2536];
        layer0[60][7:0] = buffer_data_4[2519:2512];
        layer0[60][15:8] = buffer_data_4[2527:2520];
        layer0[60][23:16] = buffer_data_4[2535:2528];
        layer0[60][31:24] = buffer_data_4[2543:2536];
        layer0[60][39:32] = buffer_data_4[2551:2544];
        layer1[60][7:0] = buffer_data_3[2519:2512];
        layer1[60][15:8] = buffer_data_3[2527:2520];
        layer1[60][23:16] = buffer_data_3[2535:2528];
        layer1[60][31:24] = buffer_data_3[2543:2536];
        layer1[60][39:32] = buffer_data_3[2551:2544];
        layer2[60][7:0] = buffer_data_2[2519:2512];
        layer2[60][15:8] = buffer_data_2[2527:2520];
        layer2[60][23:16] = buffer_data_2[2535:2528];
        layer2[60][31:24] = buffer_data_2[2543:2536];
        layer2[60][39:32] = buffer_data_2[2551:2544];
        layer3[60][7:0] = buffer_data_1[2519:2512];
        layer3[60][15:8] = buffer_data_1[2527:2520];
        layer3[60][23:16] = buffer_data_1[2535:2528];
        layer3[60][31:24] = buffer_data_1[2543:2536];
        layer3[60][39:32] = buffer_data_1[2551:2544];
        layer4[60][7:0] = buffer_data_0[2519:2512];
        layer4[60][15:8] = buffer_data_0[2527:2520];
        layer4[60][23:16] = buffer_data_0[2535:2528];
        layer4[60][31:24] = buffer_data_0[2543:2536];
        layer4[60][39:32] = buffer_data_0[2551:2544];
        layer0[61][7:0] = buffer_data_4[2527:2520];
        layer0[61][15:8] = buffer_data_4[2535:2528];
        layer0[61][23:16] = buffer_data_4[2543:2536];
        layer0[61][31:24] = buffer_data_4[2551:2544];
        layer0[61][39:32] = buffer_data_4[2559:2552];
        layer1[61][7:0] = buffer_data_3[2527:2520];
        layer1[61][15:8] = buffer_data_3[2535:2528];
        layer1[61][23:16] = buffer_data_3[2543:2536];
        layer1[61][31:24] = buffer_data_3[2551:2544];
        layer1[61][39:32] = buffer_data_3[2559:2552];
        layer2[61][7:0] = buffer_data_2[2527:2520];
        layer2[61][15:8] = buffer_data_2[2535:2528];
        layer2[61][23:16] = buffer_data_2[2543:2536];
        layer2[61][31:24] = buffer_data_2[2551:2544];
        layer2[61][39:32] = buffer_data_2[2559:2552];
        layer3[61][7:0] = buffer_data_1[2527:2520];
        layer3[61][15:8] = buffer_data_1[2535:2528];
        layer3[61][23:16] = buffer_data_1[2543:2536];
        layer3[61][31:24] = buffer_data_1[2551:2544];
        layer3[61][39:32] = buffer_data_1[2559:2552];
        layer4[61][7:0] = buffer_data_0[2527:2520];
        layer4[61][15:8] = buffer_data_0[2535:2528];
        layer4[61][23:16] = buffer_data_0[2543:2536];
        layer4[61][31:24] = buffer_data_0[2551:2544];
        layer4[61][39:32] = buffer_data_0[2559:2552];
        layer0[62][7:0] = buffer_data_4[2535:2528];
        layer0[62][15:8] = buffer_data_4[2543:2536];
        layer0[62][23:16] = buffer_data_4[2551:2544];
        layer0[62][31:24] = buffer_data_4[2559:2552];
        layer0[62][39:32] = buffer_data_4[2567:2560];
        layer1[62][7:0] = buffer_data_3[2535:2528];
        layer1[62][15:8] = buffer_data_3[2543:2536];
        layer1[62][23:16] = buffer_data_3[2551:2544];
        layer1[62][31:24] = buffer_data_3[2559:2552];
        layer1[62][39:32] = buffer_data_3[2567:2560];
        layer2[62][7:0] = buffer_data_2[2535:2528];
        layer2[62][15:8] = buffer_data_2[2543:2536];
        layer2[62][23:16] = buffer_data_2[2551:2544];
        layer2[62][31:24] = buffer_data_2[2559:2552];
        layer2[62][39:32] = buffer_data_2[2567:2560];
        layer3[62][7:0] = buffer_data_1[2535:2528];
        layer3[62][15:8] = buffer_data_1[2543:2536];
        layer3[62][23:16] = buffer_data_1[2551:2544];
        layer3[62][31:24] = buffer_data_1[2559:2552];
        layer3[62][39:32] = buffer_data_1[2567:2560];
        layer4[62][7:0] = buffer_data_0[2535:2528];
        layer4[62][15:8] = buffer_data_0[2543:2536];
        layer4[62][23:16] = buffer_data_0[2551:2544];
        layer4[62][31:24] = buffer_data_0[2559:2552];
        layer4[62][39:32] = buffer_data_0[2567:2560];
        layer0[63][7:0] = buffer_data_4[2543:2536];
        layer0[63][15:8] = buffer_data_4[2551:2544];
        layer0[63][23:16] = buffer_data_4[2559:2552];
        layer0[63][31:24] = buffer_data_4[2567:2560];
        layer0[63][39:32] = buffer_data_4[2575:2568];
        layer1[63][7:0] = buffer_data_3[2543:2536];
        layer1[63][15:8] = buffer_data_3[2551:2544];
        layer1[63][23:16] = buffer_data_3[2559:2552];
        layer1[63][31:24] = buffer_data_3[2567:2560];
        layer1[63][39:32] = buffer_data_3[2575:2568];
        layer2[63][7:0] = buffer_data_2[2543:2536];
        layer2[63][15:8] = buffer_data_2[2551:2544];
        layer2[63][23:16] = buffer_data_2[2559:2552];
        layer2[63][31:24] = buffer_data_2[2567:2560];
        layer2[63][39:32] = buffer_data_2[2575:2568];
        layer3[63][7:0] = buffer_data_1[2543:2536];
        layer3[63][15:8] = buffer_data_1[2551:2544];
        layer3[63][23:16] = buffer_data_1[2559:2552];
        layer3[63][31:24] = buffer_data_1[2567:2560];
        layer3[63][39:32] = buffer_data_1[2575:2568];
        layer4[63][7:0] = buffer_data_0[2543:2536];
        layer4[63][15:8] = buffer_data_0[2551:2544];
        layer4[63][23:16] = buffer_data_0[2559:2552];
        layer4[63][31:24] = buffer_data_0[2567:2560];
        layer4[63][39:32] = buffer_data_0[2575:2568];
    end
    ST_GAUSSIAN_5: begin
        layer0[0][7:0] = buffer_data_4[2551:2544];
        layer0[0][15:8] = buffer_data_4[2559:2552];
        layer0[0][23:16] = buffer_data_4[2567:2560];
        layer0[0][31:24] = buffer_data_4[2575:2568];
        layer0[0][39:32] = buffer_data_4[2583:2576];
        layer1[0][7:0] = buffer_data_3[2551:2544];
        layer1[0][15:8] = buffer_data_3[2559:2552];
        layer1[0][23:16] = buffer_data_3[2567:2560];
        layer1[0][31:24] = buffer_data_3[2575:2568];
        layer1[0][39:32] = buffer_data_3[2583:2576];
        layer2[0][7:0] = buffer_data_2[2551:2544];
        layer2[0][15:8] = buffer_data_2[2559:2552];
        layer2[0][23:16] = buffer_data_2[2567:2560];
        layer2[0][31:24] = buffer_data_2[2575:2568];
        layer2[0][39:32] = buffer_data_2[2583:2576];
        layer3[0][7:0] = buffer_data_1[2551:2544];
        layer3[0][15:8] = buffer_data_1[2559:2552];
        layer3[0][23:16] = buffer_data_1[2567:2560];
        layer3[0][31:24] = buffer_data_1[2575:2568];
        layer3[0][39:32] = buffer_data_1[2583:2576];
        layer4[0][7:0] = buffer_data_0[2551:2544];
        layer4[0][15:8] = buffer_data_0[2559:2552];
        layer4[0][23:16] = buffer_data_0[2567:2560];
        layer4[0][31:24] = buffer_data_0[2575:2568];
        layer4[0][39:32] = buffer_data_0[2583:2576];
        layer0[1][7:0] = buffer_data_4[2559:2552];
        layer0[1][15:8] = buffer_data_4[2567:2560];
        layer0[1][23:16] = buffer_data_4[2575:2568];
        layer0[1][31:24] = buffer_data_4[2583:2576];
        layer0[1][39:32] = buffer_data_4[2591:2584];
        layer1[1][7:0] = buffer_data_3[2559:2552];
        layer1[1][15:8] = buffer_data_3[2567:2560];
        layer1[1][23:16] = buffer_data_3[2575:2568];
        layer1[1][31:24] = buffer_data_3[2583:2576];
        layer1[1][39:32] = buffer_data_3[2591:2584];
        layer2[1][7:0] = buffer_data_2[2559:2552];
        layer2[1][15:8] = buffer_data_2[2567:2560];
        layer2[1][23:16] = buffer_data_2[2575:2568];
        layer2[1][31:24] = buffer_data_2[2583:2576];
        layer2[1][39:32] = buffer_data_2[2591:2584];
        layer3[1][7:0] = buffer_data_1[2559:2552];
        layer3[1][15:8] = buffer_data_1[2567:2560];
        layer3[1][23:16] = buffer_data_1[2575:2568];
        layer3[1][31:24] = buffer_data_1[2583:2576];
        layer3[1][39:32] = buffer_data_1[2591:2584];
        layer4[1][7:0] = buffer_data_0[2559:2552];
        layer4[1][15:8] = buffer_data_0[2567:2560];
        layer4[1][23:16] = buffer_data_0[2575:2568];
        layer4[1][31:24] = buffer_data_0[2583:2576];
        layer4[1][39:32] = buffer_data_0[2591:2584];
        layer0[2][7:0] = buffer_data_4[2567:2560];
        layer0[2][15:8] = buffer_data_4[2575:2568];
        layer0[2][23:16] = buffer_data_4[2583:2576];
        layer0[2][31:24] = buffer_data_4[2591:2584];
        layer0[2][39:32] = buffer_data_4[2599:2592];
        layer1[2][7:0] = buffer_data_3[2567:2560];
        layer1[2][15:8] = buffer_data_3[2575:2568];
        layer1[2][23:16] = buffer_data_3[2583:2576];
        layer1[2][31:24] = buffer_data_3[2591:2584];
        layer1[2][39:32] = buffer_data_3[2599:2592];
        layer2[2][7:0] = buffer_data_2[2567:2560];
        layer2[2][15:8] = buffer_data_2[2575:2568];
        layer2[2][23:16] = buffer_data_2[2583:2576];
        layer2[2][31:24] = buffer_data_2[2591:2584];
        layer2[2][39:32] = buffer_data_2[2599:2592];
        layer3[2][7:0] = buffer_data_1[2567:2560];
        layer3[2][15:8] = buffer_data_1[2575:2568];
        layer3[2][23:16] = buffer_data_1[2583:2576];
        layer3[2][31:24] = buffer_data_1[2591:2584];
        layer3[2][39:32] = buffer_data_1[2599:2592];
        layer4[2][7:0] = buffer_data_0[2567:2560];
        layer4[2][15:8] = buffer_data_0[2575:2568];
        layer4[2][23:16] = buffer_data_0[2583:2576];
        layer4[2][31:24] = buffer_data_0[2591:2584];
        layer4[2][39:32] = buffer_data_0[2599:2592];
        layer0[3][7:0] = buffer_data_4[2575:2568];
        layer0[3][15:8] = buffer_data_4[2583:2576];
        layer0[3][23:16] = buffer_data_4[2591:2584];
        layer0[3][31:24] = buffer_data_4[2599:2592];
        layer0[3][39:32] = buffer_data_4[2607:2600];
        layer1[3][7:0] = buffer_data_3[2575:2568];
        layer1[3][15:8] = buffer_data_3[2583:2576];
        layer1[3][23:16] = buffer_data_3[2591:2584];
        layer1[3][31:24] = buffer_data_3[2599:2592];
        layer1[3][39:32] = buffer_data_3[2607:2600];
        layer2[3][7:0] = buffer_data_2[2575:2568];
        layer2[3][15:8] = buffer_data_2[2583:2576];
        layer2[3][23:16] = buffer_data_2[2591:2584];
        layer2[3][31:24] = buffer_data_2[2599:2592];
        layer2[3][39:32] = buffer_data_2[2607:2600];
        layer3[3][7:0] = buffer_data_1[2575:2568];
        layer3[3][15:8] = buffer_data_1[2583:2576];
        layer3[3][23:16] = buffer_data_1[2591:2584];
        layer3[3][31:24] = buffer_data_1[2599:2592];
        layer3[3][39:32] = buffer_data_1[2607:2600];
        layer4[3][7:0] = buffer_data_0[2575:2568];
        layer4[3][15:8] = buffer_data_0[2583:2576];
        layer4[3][23:16] = buffer_data_0[2591:2584];
        layer4[3][31:24] = buffer_data_0[2599:2592];
        layer4[3][39:32] = buffer_data_0[2607:2600];
        layer0[4][7:0] = buffer_data_4[2583:2576];
        layer0[4][15:8] = buffer_data_4[2591:2584];
        layer0[4][23:16] = buffer_data_4[2599:2592];
        layer0[4][31:24] = buffer_data_4[2607:2600];
        layer0[4][39:32] = buffer_data_4[2615:2608];
        layer1[4][7:0] = buffer_data_3[2583:2576];
        layer1[4][15:8] = buffer_data_3[2591:2584];
        layer1[4][23:16] = buffer_data_3[2599:2592];
        layer1[4][31:24] = buffer_data_3[2607:2600];
        layer1[4][39:32] = buffer_data_3[2615:2608];
        layer2[4][7:0] = buffer_data_2[2583:2576];
        layer2[4][15:8] = buffer_data_2[2591:2584];
        layer2[4][23:16] = buffer_data_2[2599:2592];
        layer2[4][31:24] = buffer_data_2[2607:2600];
        layer2[4][39:32] = buffer_data_2[2615:2608];
        layer3[4][7:0] = buffer_data_1[2583:2576];
        layer3[4][15:8] = buffer_data_1[2591:2584];
        layer3[4][23:16] = buffer_data_1[2599:2592];
        layer3[4][31:24] = buffer_data_1[2607:2600];
        layer3[4][39:32] = buffer_data_1[2615:2608];
        layer4[4][7:0] = buffer_data_0[2583:2576];
        layer4[4][15:8] = buffer_data_0[2591:2584];
        layer4[4][23:16] = buffer_data_0[2599:2592];
        layer4[4][31:24] = buffer_data_0[2607:2600];
        layer4[4][39:32] = buffer_data_0[2615:2608];
        layer0[5][7:0] = buffer_data_4[2591:2584];
        layer0[5][15:8] = buffer_data_4[2599:2592];
        layer0[5][23:16] = buffer_data_4[2607:2600];
        layer0[5][31:24] = buffer_data_4[2615:2608];
        layer0[5][39:32] = buffer_data_4[2623:2616];
        layer1[5][7:0] = buffer_data_3[2591:2584];
        layer1[5][15:8] = buffer_data_3[2599:2592];
        layer1[5][23:16] = buffer_data_3[2607:2600];
        layer1[5][31:24] = buffer_data_3[2615:2608];
        layer1[5][39:32] = buffer_data_3[2623:2616];
        layer2[5][7:0] = buffer_data_2[2591:2584];
        layer2[5][15:8] = buffer_data_2[2599:2592];
        layer2[5][23:16] = buffer_data_2[2607:2600];
        layer2[5][31:24] = buffer_data_2[2615:2608];
        layer2[5][39:32] = buffer_data_2[2623:2616];
        layer3[5][7:0] = buffer_data_1[2591:2584];
        layer3[5][15:8] = buffer_data_1[2599:2592];
        layer3[5][23:16] = buffer_data_1[2607:2600];
        layer3[5][31:24] = buffer_data_1[2615:2608];
        layer3[5][39:32] = buffer_data_1[2623:2616];
        layer4[5][7:0] = buffer_data_0[2591:2584];
        layer4[5][15:8] = buffer_data_0[2599:2592];
        layer4[5][23:16] = buffer_data_0[2607:2600];
        layer4[5][31:24] = buffer_data_0[2615:2608];
        layer4[5][39:32] = buffer_data_0[2623:2616];
        layer0[6][7:0] = buffer_data_4[2599:2592];
        layer0[6][15:8] = buffer_data_4[2607:2600];
        layer0[6][23:16] = buffer_data_4[2615:2608];
        layer0[6][31:24] = buffer_data_4[2623:2616];
        layer0[6][39:32] = buffer_data_4[2631:2624];
        layer1[6][7:0] = buffer_data_3[2599:2592];
        layer1[6][15:8] = buffer_data_3[2607:2600];
        layer1[6][23:16] = buffer_data_3[2615:2608];
        layer1[6][31:24] = buffer_data_3[2623:2616];
        layer1[6][39:32] = buffer_data_3[2631:2624];
        layer2[6][7:0] = buffer_data_2[2599:2592];
        layer2[6][15:8] = buffer_data_2[2607:2600];
        layer2[6][23:16] = buffer_data_2[2615:2608];
        layer2[6][31:24] = buffer_data_2[2623:2616];
        layer2[6][39:32] = buffer_data_2[2631:2624];
        layer3[6][7:0] = buffer_data_1[2599:2592];
        layer3[6][15:8] = buffer_data_1[2607:2600];
        layer3[6][23:16] = buffer_data_1[2615:2608];
        layer3[6][31:24] = buffer_data_1[2623:2616];
        layer3[6][39:32] = buffer_data_1[2631:2624];
        layer4[6][7:0] = buffer_data_0[2599:2592];
        layer4[6][15:8] = buffer_data_0[2607:2600];
        layer4[6][23:16] = buffer_data_0[2615:2608];
        layer4[6][31:24] = buffer_data_0[2623:2616];
        layer4[6][39:32] = buffer_data_0[2631:2624];
        layer0[7][7:0] = buffer_data_4[2607:2600];
        layer0[7][15:8] = buffer_data_4[2615:2608];
        layer0[7][23:16] = buffer_data_4[2623:2616];
        layer0[7][31:24] = buffer_data_4[2631:2624];
        layer0[7][39:32] = buffer_data_4[2639:2632];
        layer1[7][7:0] = buffer_data_3[2607:2600];
        layer1[7][15:8] = buffer_data_3[2615:2608];
        layer1[7][23:16] = buffer_data_3[2623:2616];
        layer1[7][31:24] = buffer_data_3[2631:2624];
        layer1[7][39:32] = buffer_data_3[2639:2632];
        layer2[7][7:0] = buffer_data_2[2607:2600];
        layer2[7][15:8] = buffer_data_2[2615:2608];
        layer2[7][23:16] = buffer_data_2[2623:2616];
        layer2[7][31:24] = buffer_data_2[2631:2624];
        layer2[7][39:32] = buffer_data_2[2639:2632];
        layer3[7][7:0] = buffer_data_1[2607:2600];
        layer3[7][15:8] = buffer_data_1[2615:2608];
        layer3[7][23:16] = buffer_data_1[2623:2616];
        layer3[7][31:24] = buffer_data_1[2631:2624];
        layer3[7][39:32] = buffer_data_1[2639:2632];
        layer4[7][7:0] = buffer_data_0[2607:2600];
        layer4[7][15:8] = buffer_data_0[2615:2608];
        layer4[7][23:16] = buffer_data_0[2623:2616];
        layer4[7][31:24] = buffer_data_0[2631:2624];
        layer4[7][39:32] = buffer_data_0[2639:2632];
        layer0[8][7:0] = buffer_data_4[2615:2608];
        layer0[8][15:8] = buffer_data_4[2623:2616];
        layer0[8][23:16] = buffer_data_4[2631:2624];
        layer0[8][31:24] = buffer_data_4[2639:2632];
        layer0[8][39:32] = buffer_data_4[2647:2640];
        layer1[8][7:0] = buffer_data_3[2615:2608];
        layer1[8][15:8] = buffer_data_3[2623:2616];
        layer1[8][23:16] = buffer_data_3[2631:2624];
        layer1[8][31:24] = buffer_data_3[2639:2632];
        layer1[8][39:32] = buffer_data_3[2647:2640];
        layer2[8][7:0] = buffer_data_2[2615:2608];
        layer2[8][15:8] = buffer_data_2[2623:2616];
        layer2[8][23:16] = buffer_data_2[2631:2624];
        layer2[8][31:24] = buffer_data_2[2639:2632];
        layer2[8][39:32] = buffer_data_2[2647:2640];
        layer3[8][7:0] = buffer_data_1[2615:2608];
        layer3[8][15:8] = buffer_data_1[2623:2616];
        layer3[8][23:16] = buffer_data_1[2631:2624];
        layer3[8][31:24] = buffer_data_1[2639:2632];
        layer3[8][39:32] = buffer_data_1[2647:2640];
        layer4[8][7:0] = buffer_data_0[2615:2608];
        layer4[8][15:8] = buffer_data_0[2623:2616];
        layer4[8][23:16] = buffer_data_0[2631:2624];
        layer4[8][31:24] = buffer_data_0[2639:2632];
        layer4[8][39:32] = buffer_data_0[2647:2640];
        layer0[9][7:0] = buffer_data_4[2623:2616];
        layer0[9][15:8] = buffer_data_4[2631:2624];
        layer0[9][23:16] = buffer_data_4[2639:2632];
        layer0[9][31:24] = buffer_data_4[2647:2640];
        layer0[9][39:32] = buffer_data_4[2655:2648];
        layer1[9][7:0] = buffer_data_3[2623:2616];
        layer1[9][15:8] = buffer_data_3[2631:2624];
        layer1[9][23:16] = buffer_data_3[2639:2632];
        layer1[9][31:24] = buffer_data_3[2647:2640];
        layer1[9][39:32] = buffer_data_3[2655:2648];
        layer2[9][7:0] = buffer_data_2[2623:2616];
        layer2[9][15:8] = buffer_data_2[2631:2624];
        layer2[9][23:16] = buffer_data_2[2639:2632];
        layer2[9][31:24] = buffer_data_2[2647:2640];
        layer2[9][39:32] = buffer_data_2[2655:2648];
        layer3[9][7:0] = buffer_data_1[2623:2616];
        layer3[9][15:8] = buffer_data_1[2631:2624];
        layer3[9][23:16] = buffer_data_1[2639:2632];
        layer3[9][31:24] = buffer_data_1[2647:2640];
        layer3[9][39:32] = buffer_data_1[2655:2648];
        layer4[9][7:0] = buffer_data_0[2623:2616];
        layer4[9][15:8] = buffer_data_0[2631:2624];
        layer4[9][23:16] = buffer_data_0[2639:2632];
        layer4[9][31:24] = buffer_data_0[2647:2640];
        layer4[9][39:32] = buffer_data_0[2655:2648];
        layer0[10][7:0] = buffer_data_4[2631:2624];
        layer0[10][15:8] = buffer_data_4[2639:2632];
        layer0[10][23:16] = buffer_data_4[2647:2640];
        layer0[10][31:24] = buffer_data_4[2655:2648];
        layer0[10][39:32] = buffer_data_4[2663:2656];
        layer1[10][7:0] = buffer_data_3[2631:2624];
        layer1[10][15:8] = buffer_data_3[2639:2632];
        layer1[10][23:16] = buffer_data_3[2647:2640];
        layer1[10][31:24] = buffer_data_3[2655:2648];
        layer1[10][39:32] = buffer_data_3[2663:2656];
        layer2[10][7:0] = buffer_data_2[2631:2624];
        layer2[10][15:8] = buffer_data_2[2639:2632];
        layer2[10][23:16] = buffer_data_2[2647:2640];
        layer2[10][31:24] = buffer_data_2[2655:2648];
        layer2[10][39:32] = buffer_data_2[2663:2656];
        layer3[10][7:0] = buffer_data_1[2631:2624];
        layer3[10][15:8] = buffer_data_1[2639:2632];
        layer3[10][23:16] = buffer_data_1[2647:2640];
        layer3[10][31:24] = buffer_data_1[2655:2648];
        layer3[10][39:32] = buffer_data_1[2663:2656];
        layer4[10][7:0] = buffer_data_0[2631:2624];
        layer4[10][15:8] = buffer_data_0[2639:2632];
        layer4[10][23:16] = buffer_data_0[2647:2640];
        layer4[10][31:24] = buffer_data_0[2655:2648];
        layer4[10][39:32] = buffer_data_0[2663:2656];
        layer0[11][7:0] = buffer_data_4[2639:2632];
        layer0[11][15:8] = buffer_data_4[2647:2640];
        layer0[11][23:16] = buffer_data_4[2655:2648];
        layer0[11][31:24] = buffer_data_4[2663:2656];
        layer0[11][39:32] = buffer_data_4[2671:2664];
        layer1[11][7:0] = buffer_data_3[2639:2632];
        layer1[11][15:8] = buffer_data_3[2647:2640];
        layer1[11][23:16] = buffer_data_3[2655:2648];
        layer1[11][31:24] = buffer_data_3[2663:2656];
        layer1[11][39:32] = buffer_data_3[2671:2664];
        layer2[11][7:0] = buffer_data_2[2639:2632];
        layer2[11][15:8] = buffer_data_2[2647:2640];
        layer2[11][23:16] = buffer_data_2[2655:2648];
        layer2[11][31:24] = buffer_data_2[2663:2656];
        layer2[11][39:32] = buffer_data_2[2671:2664];
        layer3[11][7:0] = buffer_data_1[2639:2632];
        layer3[11][15:8] = buffer_data_1[2647:2640];
        layer3[11][23:16] = buffer_data_1[2655:2648];
        layer3[11][31:24] = buffer_data_1[2663:2656];
        layer3[11][39:32] = buffer_data_1[2671:2664];
        layer4[11][7:0] = buffer_data_0[2639:2632];
        layer4[11][15:8] = buffer_data_0[2647:2640];
        layer4[11][23:16] = buffer_data_0[2655:2648];
        layer4[11][31:24] = buffer_data_0[2663:2656];
        layer4[11][39:32] = buffer_data_0[2671:2664];
        layer0[12][7:0] = buffer_data_4[2647:2640];
        layer0[12][15:8] = buffer_data_4[2655:2648];
        layer0[12][23:16] = buffer_data_4[2663:2656];
        layer0[12][31:24] = buffer_data_4[2671:2664];
        layer0[12][39:32] = buffer_data_4[2679:2672];
        layer1[12][7:0] = buffer_data_3[2647:2640];
        layer1[12][15:8] = buffer_data_3[2655:2648];
        layer1[12][23:16] = buffer_data_3[2663:2656];
        layer1[12][31:24] = buffer_data_3[2671:2664];
        layer1[12][39:32] = buffer_data_3[2679:2672];
        layer2[12][7:0] = buffer_data_2[2647:2640];
        layer2[12][15:8] = buffer_data_2[2655:2648];
        layer2[12][23:16] = buffer_data_2[2663:2656];
        layer2[12][31:24] = buffer_data_2[2671:2664];
        layer2[12][39:32] = buffer_data_2[2679:2672];
        layer3[12][7:0] = buffer_data_1[2647:2640];
        layer3[12][15:8] = buffer_data_1[2655:2648];
        layer3[12][23:16] = buffer_data_1[2663:2656];
        layer3[12][31:24] = buffer_data_1[2671:2664];
        layer3[12][39:32] = buffer_data_1[2679:2672];
        layer4[12][7:0] = buffer_data_0[2647:2640];
        layer4[12][15:8] = buffer_data_0[2655:2648];
        layer4[12][23:16] = buffer_data_0[2663:2656];
        layer4[12][31:24] = buffer_data_0[2671:2664];
        layer4[12][39:32] = buffer_data_0[2679:2672];
        layer0[13][7:0] = buffer_data_4[2655:2648];
        layer0[13][15:8] = buffer_data_4[2663:2656];
        layer0[13][23:16] = buffer_data_4[2671:2664];
        layer0[13][31:24] = buffer_data_4[2679:2672];
        layer0[13][39:32] = buffer_data_4[2687:2680];
        layer1[13][7:0] = buffer_data_3[2655:2648];
        layer1[13][15:8] = buffer_data_3[2663:2656];
        layer1[13][23:16] = buffer_data_3[2671:2664];
        layer1[13][31:24] = buffer_data_3[2679:2672];
        layer1[13][39:32] = buffer_data_3[2687:2680];
        layer2[13][7:0] = buffer_data_2[2655:2648];
        layer2[13][15:8] = buffer_data_2[2663:2656];
        layer2[13][23:16] = buffer_data_2[2671:2664];
        layer2[13][31:24] = buffer_data_2[2679:2672];
        layer2[13][39:32] = buffer_data_2[2687:2680];
        layer3[13][7:0] = buffer_data_1[2655:2648];
        layer3[13][15:8] = buffer_data_1[2663:2656];
        layer3[13][23:16] = buffer_data_1[2671:2664];
        layer3[13][31:24] = buffer_data_1[2679:2672];
        layer3[13][39:32] = buffer_data_1[2687:2680];
        layer4[13][7:0] = buffer_data_0[2655:2648];
        layer4[13][15:8] = buffer_data_0[2663:2656];
        layer4[13][23:16] = buffer_data_0[2671:2664];
        layer4[13][31:24] = buffer_data_0[2679:2672];
        layer4[13][39:32] = buffer_data_0[2687:2680];
        layer0[14][7:0] = buffer_data_4[2663:2656];
        layer0[14][15:8] = buffer_data_4[2671:2664];
        layer0[14][23:16] = buffer_data_4[2679:2672];
        layer0[14][31:24] = buffer_data_4[2687:2680];
        layer0[14][39:32] = buffer_data_4[2695:2688];
        layer1[14][7:0] = buffer_data_3[2663:2656];
        layer1[14][15:8] = buffer_data_3[2671:2664];
        layer1[14][23:16] = buffer_data_3[2679:2672];
        layer1[14][31:24] = buffer_data_3[2687:2680];
        layer1[14][39:32] = buffer_data_3[2695:2688];
        layer2[14][7:0] = buffer_data_2[2663:2656];
        layer2[14][15:8] = buffer_data_2[2671:2664];
        layer2[14][23:16] = buffer_data_2[2679:2672];
        layer2[14][31:24] = buffer_data_2[2687:2680];
        layer2[14][39:32] = buffer_data_2[2695:2688];
        layer3[14][7:0] = buffer_data_1[2663:2656];
        layer3[14][15:8] = buffer_data_1[2671:2664];
        layer3[14][23:16] = buffer_data_1[2679:2672];
        layer3[14][31:24] = buffer_data_1[2687:2680];
        layer3[14][39:32] = buffer_data_1[2695:2688];
        layer4[14][7:0] = buffer_data_0[2663:2656];
        layer4[14][15:8] = buffer_data_0[2671:2664];
        layer4[14][23:16] = buffer_data_0[2679:2672];
        layer4[14][31:24] = buffer_data_0[2687:2680];
        layer4[14][39:32] = buffer_data_0[2695:2688];
        layer0[15][7:0] = buffer_data_4[2671:2664];
        layer0[15][15:8] = buffer_data_4[2679:2672];
        layer0[15][23:16] = buffer_data_4[2687:2680];
        layer0[15][31:24] = buffer_data_4[2695:2688];
        layer0[15][39:32] = buffer_data_4[2703:2696];
        layer1[15][7:0] = buffer_data_3[2671:2664];
        layer1[15][15:8] = buffer_data_3[2679:2672];
        layer1[15][23:16] = buffer_data_3[2687:2680];
        layer1[15][31:24] = buffer_data_3[2695:2688];
        layer1[15][39:32] = buffer_data_3[2703:2696];
        layer2[15][7:0] = buffer_data_2[2671:2664];
        layer2[15][15:8] = buffer_data_2[2679:2672];
        layer2[15][23:16] = buffer_data_2[2687:2680];
        layer2[15][31:24] = buffer_data_2[2695:2688];
        layer2[15][39:32] = buffer_data_2[2703:2696];
        layer3[15][7:0] = buffer_data_1[2671:2664];
        layer3[15][15:8] = buffer_data_1[2679:2672];
        layer3[15][23:16] = buffer_data_1[2687:2680];
        layer3[15][31:24] = buffer_data_1[2695:2688];
        layer3[15][39:32] = buffer_data_1[2703:2696];
        layer4[15][7:0] = buffer_data_0[2671:2664];
        layer4[15][15:8] = buffer_data_0[2679:2672];
        layer4[15][23:16] = buffer_data_0[2687:2680];
        layer4[15][31:24] = buffer_data_0[2695:2688];
        layer4[15][39:32] = buffer_data_0[2703:2696];
        layer0[16][7:0] = buffer_data_4[2679:2672];
        layer0[16][15:8] = buffer_data_4[2687:2680];
        layer0[16][23:16] = buffer_data_4[2695:2688];
        layer0[16][31:24] = buffer_data_4[2703:2696];
        layer0[16][39:32] = buffer_data_4[2711:2704];
        layer1[16][7:0] = buffer_data_3[2679:2672];
        layer1[16][15:8] = buffer_data_3[2687:2680];
        layer1[16][23:16] = buffer_data_3[2695:2688];
        layer1[16][31:24] = buffer_data_3[2703:2696];
        layer1[16][39:32] = buffer_data_3[2711:2704];
        layer2[16][7:0] = buffer_data_2[2679:2672];
        layer2[16][15:8] = buffer_data_2[2687:2680];
        layer2[16][23:16] = buffer_data_2[2695:2688];
        layer2[16][31:24] = buffer_data_2[2703:2696];
        layer2[16][39:32] = buffer_data_2[2711:2704];
        layer3[16][7:0] = buffer_data_1[2679:2672];
        layer3[16][15:8] = buffer_data_1[2687:2680];
        layer3[16][23:16] = buffer_data_1[2695:2688];
        layer3[16][31:24] = buffer_data_1[2703:2696];
        layer3[16][39:32] = buffer_data_1[2711:2704];
        layer4[16][7:0] = buffer_data_0[2679:2672];
        layer4[16][15:8] = buffer_data_0[2687:2680];
        layer4[16][23:16] = buffer_data_0[2695:2688];
        layer4[16][31:24] = buffer_data_0[2703:2696];
        layer4[16][39:32] = buffer_data_0[2711:2704];
        layer0[17][7:0] = buffer_data_4[2687:2680];
        layer0[17][15:8] = buffer_data_4[2695:2688];
        layer0[17][23:16] = buffer_data_4[2703:2696];
        layer0[17][31:24] = buffer_data_4[2711:2704];
        layer0[17][39:32] = buffer_data_4[2719:2712];
        layer1[17][7:0] = buffer_data_3[2687:2680];
        layer1[17][15:8] = buffer_data_3[2695:2688];
        layer1[17][23:16] = buffer_data_3[2703:2696];
        layer1[17][31:24] = buffer_data_3[2711:2704];
        layer1[17][39:32] = buffer_data_3[2719:2712];
        layer2[17][7:0] = buffer_data_2[2687:2680];
        layer2[17][15:8] = buffer_data_2[2695:2688];
        layer2[17][23:16] = buffer_data_2[2703:2696];
        layer2[17][31:24] = buffer_data_2[2711:2704];
        layer2[17][39:32] = buffer_data_2[2719:2712];
        layer3[17][7:0] = buffer_data_1[2687:2680];
        layer3[17][15:8] = buffer_data_1[2695:2688];
        layer3[17][23:16] = buffer_data_1[2703:2696];
        layer3[17][31:24] = buffer_data_1[2711:2704];
        layer3[17][39:32] = buffer_data_1[2719:2712];
        layer4[17][7:0] = buffer_data_0[2687:2680];
        layer4[17][15:8] = buffer_data_0[2695:2688];
        layer4[17][23:16] = buffer_data_0[2703:2696];
        layer4[17][31:24] = buffer_data_0[2711:2704];
        layer4[17][39:32] = buffer_data_0[2719:2712];
        layer0[18][7:0] = buffer_data_4[2695:2688];
        layer0[18][15:8] = buffer_data_4[2703:2696];
        layer0[18][23:16] = buffer_data_4[2711:2704];
        layer0[18][31:24] = buffer_data_4[2719:2712];
        layer0[18][39:32] = buffer_data_4[2727:2720];
        layer1[18][7:0] = buffer_data_3[2695:2688];
        layer1[18][15:8] = buffer_data_3[2703:2696];
        layer1[18][23:16] = buffer_data_3[2711:2704];
        layer1[18][31:24] = buffer_data_3[2719:2712];
        layer1[18][39:32] = buffer_data_3[2727:2720];
        layer2[18][7:0] = buffer_data_2[2695:2688];
        layer2[18][15:8] = buffer_data_2[2703:2696];
        layer2[18][23:16] = buffer_data_2[2711:2704];
        layer2[18][31:24] = buffer_data_2[2719:2712];
        layer2[18][39:32] = buffer_data_2[2727:2720];
        layer3[18][7:0] = buffer_data_1[2695:2688];
        layer3[18][15:8] = buffer_data_1[2703:2696];
        layer3[18][23:16] = buffer_data_1[2711:2704];
        layer3[18][31:24] = buffer_data_1[2719:2712];
        layer3[18][39:32] = buffer_data_1[2727:2720];
        layer4[18][7:0] = buffer_data_0[2695:2688];
        layer4[18][15:8] = buffer_data_0[2703:2696];
        layer4[18][23:16] = buffer_data_0[2711:2704];
        layer4[18][31:24] = buffer_data_0[2719:2712];
        layer4[18][39:32] = buffer_data_0[2727:2720];
        layer0[19][7:0] = buffer_data_4[2703:2696];
        layer0[19][15:8] = buffer_data_4[2711:2704];
        layer0[19][23:16] = buffer_data_4[2719:2712];
        layer0[19][31:24] = buffer_data_4[2727:2720];
        layer0[19][39:32] = buffer_data_4[2735:2728];
        layer1[19][7:0] = buffer_data_3[2703:2696];
        layer1[19][15:8] = buffer_data_3[2711:2704];
        layer1[19][23:16] = buffer_data_3[2719:2712];
        layer1[19][31:24] = buffer_data_3[2727:2720];
        layer1[19][39:32] = buffer_data_3[2735:2728];
        layer2[19][7:0] = buffer_data_2[2703:2696];
        layer2[19][15:8] = buffer_data_2[2711:2704];
        layer2[19][23:16] = buffer_data_2[2719:2712];
        layer2[19][31:24] = buffer_data_2[2727:2720];
        layer2[19][39:32] = buffer_data_2[2735:2728];
        layer3[19][7:0] = buffer_data_1[2703:2696];
        layer3[19][15:8] = buffer_data_1[2711:2704];
        layer3[19][23:16] = buffer_data_1[2719:2712];
        layer3[19][31:24] = buffer_data_1[2727:2720];
        layer3[19][39:32] = buffer_data_1[2735:2728];
        layer4[19][7:0] = buffer_data_0[2703:2696];
        layer4[19][15:8] = buffer_data_0[2711:2704];
        layer4[19][23:16] = buffer_data_0[2719:2712];
        layer4[19][31:24] = buffer_data_0[2727:2720];
        layer4[19][39:32] = buffer_data_0[2735:2728];
        layer0[20][7:0] = buffer_data_4[2711:2704];
        layer0[20][15:8] = buffer_data_4[2719:2712];
        layer0[20][23:16] = buffer_data_4[2727:2720];
        layer0[20][31:24] = buffer_data_4[2735:2728];
        layer0[20][39:32] = buffer_data_4[2743:2736];
        layer1[20][7:0] = buffer_data_3[2711:2704];
        layer1[20][15:8] = buffer_data_3[2719:2712];
        layer1[20][23:16] = buffer_data_3[2727:2720];
        layer1[20][31:24] = buffer_data_3[2735:2728];
        layer1[20][39:32] = buffer_data_3[2743:2736];
        layer2[20][7:0] = buffer_data_2[2711:2704];
        layer2[20][15:8] = buffer_data_2[2719:2712];
        layer2[20][23:16] = buffer_data_2[2727:2720];
        layer2[20][31:24] = buffer_data_2[2735:2728];
        layer2[20][39:32] = buffer_data_2[2743:2736];
        layer3[20][7:0] = buffer_data_1[2711:2704];
        layer3[20][15:8] = buffer_data_1[2719:2712];
        layer3[20][23:16] = buffer_data_1[2727:2720];
        layer3[20][31:24] = buffer_data_1[2735:2728];
        layer3[20][39:32] = buffer_data_1[2743:2736];
        layer4[20][7:0] = buffer_data_0[2711:2704];
        layer4[20][15:8] = buffer_data_0[2719:2712];
        layer4[20][23:16] = buffer_data_0[2727:2720];
        layer4[20][31:24] = buffer_data_0[2735:2728];
        layer4[20][39:32] = buffer_data_0[2743:2736];
        layer0[21][7:0] = buffer_data_4[2719:2712];
        layer0[21][15:8] = buffer_data_4[2727:2720];
        layer0[21][23:16] = buffer_data_4[2735:2728];
        layer0[21][31:24] = buffer_data_4[2743:2736];
        layer0[21][39:32] = buffer_data_4[2751:2744];
        layer1[21][7:0] = buffer_data_3[2719:2712];
        layer1[21][15:8] = buffer_data_3[2727:2720];
        layer1[21][23:16] = buffer_data_3[2735:2728];
        layer1[21][31:24] = buffer_data_3[2743:2736];
        layer1[21][39:32] = buffer_data_3[2751:2744];
        layer2[21][7:0] = buffer_data_2[2719:2712];
        layer2[21][15:8] = buffer_data_2[2727:2720];
        layer2[21][23:16] = buffer_data_2[2735:2728];
        layer2[21][31:24] = buffer_data_2[2743:2736];
        layer2[21][39:32] = buffer_data_2[2751:2744];
        layer3[21][7:0] = buffer_data_1[2719:2712];
        layer3[21][15:8] = buffer_data_1[2727:2720];
        layer3[21][23:16] = buffer_data_1[2735:2728];
        layer3[21][31:24] = buffer_data_1[2743:2736];
        layer3[21][39:32] = buffer_data_1[2751:2744];
        layer4[21][7:0] = buffer_data_0[2719:2712];
        layer4[21][15:8] = buffer_data_0[2727:2720];
        layer4[21][23:16] = buffer_data_0[2735:2728];
        layer4[21][31:24] = buffer_data_0[2743:2736];
        layer4[21][39:32] = buffer_data_0[2751:2744];
        layer0[22][7:0] = buffer_data_4[2727:2720];
        layer0[22][15:8] = buffer_data_4[2735:2728];
        layer0[22][23:16] = buffer_data_4[2743:2736];
        layer0[22][31:24] = buffer_data_4[2751:2744];
        layer0[22][39:32] = buffer_data_4[2759:2752];
        layer1[22][7:0] = buffer_data_3[2727:2720];
        layer1[22][15:8] = buffer_data_3[2735:2728];
        layer1[22][23:16] = buffer_data_3[2743:2736];
        layer1[22][31:24] = buffer_data_3[2751:2744];
        layer1[22][39:32] = buffer_data_3[2759:2752];
        layer2[22][7:0] = buffer_data_2[2727:2720];
        layer2[22][15:8] = buffer_data_2[2735:2728];
        layer2[22][23:16] = buffer_data_2[2743:2736];
        layer2[22][31:24] = buffer_data_2[2751:2744];
        layer2[22][39:32] = buffer_data_2[2759:2752];
        layer3[22][7:0] = buffer_data_1[2727:2720];
        layer3[22][15:8] = buffer_data_1[2735:2728];
        layer3[22][23:16] = buffer_data_1[2743:2736];
        layer3[22][31:24] = buffer_data_1[2751:2744];
        layer3[22][39:32] = buffer_data_1[2759:2752];
        layer4[22][7:0] = buffer_data_0[2727:2720];
        layer4[22][15:8] = buffer_data_0[2735:2728];
        layer4[22][23:16] = buffer_data_0[2743:2736];
        layer4[22][31:24] = buffer_data_0[2751:2744];
        layer4[22][39:32] = buffer_data_0[2759:2752];
        layer0[23][7:0] = buffer_data_4[2735:2728];
        layer0[23][15:8] = buffer_data_4[2743:2736];
        layer0[23][23:16] = buffer_data_4[2751:2744];
        layer0[23][31:24] = buffer_data_4[2759:2752];
        layer0[23][39:32] = buffer_data_4[2767:2760];
        layer1[23][7:0] = buffer_data_3[2735:2728];
        layer1[23][15:8] = buffer_data_3[2743:2736];
        layer1[23][23:16] = buffer_data_3[2751:2744];
        layer1[23][31:24] = buffer_data_3[2759:2752];
        layer1[23][39:32] = buffer_data_3[2767:2760];
        layer2[23][7:0] = buffer_data_2[2735:2728];
        layer2[23][15:8] = buffer_data_2[2743:2736];
        layer2[23][23:16] = buffer_data_2[2751:2744];
        layer2[23][31:24] = buffer_data_2[2759:2752];
        layer2[23][39:32] = buffer_data_2[2767:2760];
        layer3[23][7:0] = buffer_data_1[2735:2728];
        layer3[23][15:8] = buffer_data_1[2743:2736];
        layer3[23][23:16] = buffer_data_1[2751:2744];
        layer3[23][31:24] = buffer_data_1[2759:2752];
        layer3[23][39:32] = buffer_data_1[2767:2760];
        layer4[23][7:0] = buffer_data_0[2735:2728];
        layer4[23][15:8] = buffer_data_0[2743:2736];
        layer4[23][23:16] = buffer_data_0[2751:2744];
        layer4[23][31:24] = buffer_data_0[2759:2752];
        layer4[23][39:32] = buffer_data_0[2767:2760];
        layer0[24][7:0] = buffer_data_4[2743:2736];
        layer0[24][15:8] = buffer_data_4[2751:2744];
        layer0[24][23:16] = buffer_data_4[2759:2752];
        layer0[24][31:24] = buffer_data_4[2767:2760];
        layer0[24][39:32] = buffer_data_4[2775:2768];
        layer1[24][7:0] = buffer_data_3[2743:2736];
        layer1[24][15:8] = buffer_data_3[2751:2744];
        layer1[24][23:16] = buffer_data_3[2759:2752];
        layer1[24][31:24] = buffer_data_3[2767:2760];
        layer1[24][39:32] = buffer_data_3[2775:2768];
        layer2[24][7:0] = buffer_data_2[2743:2736];
        layer2[24][15:8] = buffer_data_2[2751:2744];
        layer2[24][23:16] = buffer_data_2[2759:2752];
        layer2[24][31:24] = buffer_data_2[2767:2760];
        layer2[24][39:32] = buffer_data_2[2775:2768];
        layer3[24][7:0] = buffer_data_1[2743:2736];
        layer3[24][15:8] = buffer_data_1[2751:2744];
        layer3[24][23:16] = buffer_data_1[2759:2752];
        layer3[24][31:24] = buffer_data_1[2767:2760];
        layer3[24][39:32] = buffer_data_1[2775:2768];
        layer4[24][7:0] = buffer_data_0[2743:2736];
        layer4[24][15:8] = buffer_data_0[2751:2744];
        layer4[24][23:16] = buffer_data_0[2759:2752];
        layer4[24][31:24] = buffer_data_0[2767:2760];
        layer4[24][39:32] = buffer_data_0[2775:2768];
        layer0[25][7:0] = buffer_data_4[2751:2744];
        layer0[25][15:8] = buffer_data_4[2759:2752];
        layer0[25][23:16] = buffer_data_4[2767:2760];
        layer0[25][31:24] = buffer_data_4[2775:2768];
        layer0[25][39:32] = buffer_data_4[2783:2776];
        layer1[25][7:0] = buffer_data_3[2751:2744];
        layer1[25][15:8] = buffer_data_3[2759:2752];
        layer1[25][23:16] = buffer_data_3[2767:2760];
        layer1[25][31:24] = buffer_data_3[2775:2768];
        layer1[25][39:32] = buffer_data_3[2783:2776];
        layer2[25][7:0] = buffer_data_2[2751:2744];
        layer2[25][15:8] = buffer_data_2[2759:2752];
        layer2[25][23:16] = buffer_data_2[2767:2760];
        layer2[25][31:24] = buffer_data_2[2775:2768];
        layer2[25][39:32] = buffer_data_2[2783:2776];
        layer3[25][7:0] = buffer_data_1[2751:2744];
        layer3[25][15:8] = buffer_data_1[2759:2752];
        layer3[25][23:16] = buffer_data_1[2767:2760];
        layer3[25][31:24] = buffer_data_1[2775:2768];
        layer3[25][39:32] = buffer_data_1[2783:2776];
        layer4[25][7:0] = buffer_data_0[2751:2744];
        layer4[25][15:8] = buffer_data_0[2759:2752];
        layer4[25][23:16] = buffer_data_0[2767:2760];
        layer4[25][31:24] = buffer_data_0[2775:2768];
        layer4[25][39:32] = buffer_data_0[2783:2776];
        layer0[26][7:0] = buffer_data_4[2759:2752];
        layer0[26][15:8] = buffer_data_4[2767:2760];
        layer0[26][23:16] = buffer_data_4[2775:2768];
        layer0[26][31:24] = buffer_data_4[2783:2776];
        layer0[26][39:32] = buffer_data_4[2791:2784];
        layer1[26][7:0] = buffer_data_3[2759:2752];
        layer1[26][15:8] = buffer_data_3[2767:2760];
        layer1[26][23:16] = buffer_data_3[2775:2768];
        layer1[26][31:24] = buffer_data_3[2783:2776];
        layer1[26][39:32] = buffer_data_3[2791:2784];
        layer2[26][7:0] = buffer_data_2[2759:2752];
        layer2[26][15:8] = buffer_data_2[2767:2760];
        layer2[26][23:16] = buffer_data_2[2775:2768];
        layer2[26][31:24] = buffer_data_2[2783:2776];
        layer2[26][39:32] = buffer_data_2[2791:2784];
        layer3[26][7:0] = buffer_data_1[2759:2752];
        layer3[26][15:8] = buffer_data_1[2767:2760];
        layer3[26][23:16] = buffer_data_1[2775:2768];
        layer3[26][31:24] = buffer_data_1[2783:2776];
        layer3[26][39:32] = buffer_data_1[2791:2784];
        layer4[26][7:0] = buffer_data_0[2759:2752];
        layer4[26][15:8] = buffer_data_0[2767:2760];
        layer4[26][23:16] = buffer_data_0[2775:2768];
        layer4[26][31:24] = buffer_data_0[2783:2776];
        layer4[26][39:32] = buffer_data_0[2791:2784];
        layer0[27][7:0] = buffer_data_4[2767:2760];
        layer0[27][15:8] = buffer_data_4[2775:2768];
        layer0[27][23:16] = buffer_data_4[2783:2776];
        layer0[27][31:24] = buffer_data_4[2791:2784];
        layer0[27][39:32] = buffer_data_4[2799:2792];
        layer1[27][7:0] = buffer_data_3[2767:2760];
        layer1[27][15:8] = buffer_data_3[2775:2768];
        layer1[27][23:16] = buffer_data_3[2783:2776];
        layer1[27][31:24] = buffer_data_3[2791:2784];
        layer1[27][39:32] = buffer_data_3[2799:2792];
        layer2[27][7:0] = buffer_data_2[2767:2760];
        layer2[27][15:8] = buffer_data_2[2775:2768];
        layer2[27][23:16] = buffer_data_2[2783:2776];
        layer2[27][31:24] = buffer_data_2[2791:2784];
        layer2[27][39:32] = buffer_data_2[2799:2792];
        layer3[27][7:0] = buffer_data_1[2767:2760];
        layer3[27][15:8] = buffer_data_1[2775:2768];
        layer3[27][23:16] = buffer_data_1[2783:2776];
        layer3[27][31:24] = buffer_data_1[2791:2784];
        layer3[27][39:32] = buffer_data_1[2799:2792];
        layer4[27][7:0] = buffer_data_0[2767:2760];
        layer4[27][15:8] = buffer_data_0[2775:2768];
        layer4[27][23:16] = buffer_data_0[2783:2776];
        layer4[27][31:24] = buffer_data_0[2791:2784];
        layer4[27][39:32] = buffer_data_0[2799:2792];
        layer0[28][7:0] = buffer_data_4[2775:2768];
        layer0[28][15:8] = buffer_data_4[2783:2776];
        layer0[28][23:16] = buffer_data_4[2791:2784];
        layer0[28][31:24] = buffer_data_4[2799:2792];
        layer0[28][39:32] = buffer_data_4[2807:2800];
        layer1[28][7:0] = buffer_data_3[2775:2768];
        layer1[28][15:8] = buffer_data_3[2783:2776];
        layer1[28][23:16] = buffer_data_3[2791:2784];
        layer1[28][31:24] = buffer_data_3[2799:2792];
        layer1[28][39:32] = buffer_data_3[2807:2800];
        layer2[28][7:0] = buffer_data_2[2775:2768];
        layer2[28][15:8] = buffer_data_2[2783:2776];
        layer2[28][23:16] = buffer_data_2[2791:2784];
        layer2[28][31:24] = buffer_data_2[2799:2792];
        layer2[28][39:32] = buffer_data_2[2807:2800];
        layer3[28][7:0] = buffer_data_1[2775:2768];
        layer3[28][15:8] = buffer_data_1[2783:2776];
        layer3[28][23:16] = buffer_data_1[2791:2784];
        layer3[28][31:24] = buffer_data_1[2799:2792];
        layer3[28][39:32] = buffer_data_1[2807:2800];
        layer4[28][7:0] = buffer_data_0[2775:2768];
        layer4[28][15:8] = buffer_data_0[2783:2776];
        layer4[28][23:16] = buffer_data_0[2791:2784];
        layer4[28][31:24] = buffer_data_0[2799:2792];
        layer4[28][39:32] = buffer_data_0[2807:2800];
        layer0[29][7:0] = buffer_data_4[2783:2776];
        layer0[29][15:8] = buffer_data_4[2791:2784];
        layer0[29][23:16] = buffer_data_4[2799:2792];
        layer0[29][31:24] = buffer_data_4[2807:2800];
        layer0[29][39:32] = buffer_data_4[2815:2808];
        layer1[29][7:0] = buffer_data_3[2783:2776];
        layer1[29][15:8] = buffer_data_3[2791:2784];
        layer1[29][23:16] = buffer_data_3[2799:2792];
        layer1[29][31:24] = buffer_data_3[2807:2800];
        layer1[29][39:32] = buffer_data_3[2815:2808];
        layer2[29][7:0] = buffer_data_2[2783:2776];
        layer2[29][15:8] = buffer_data_2[2791:2784];
        layer2[29][23:16] = buffer_data_2[2799:2792];
        layer2[29][31:24] = buffer_data_2[2807:2800];
        layer2[29][39:32] = buffer_data_2[2815:2808];
        layer3[29][7:0] = buffer_data_1[2783:2776];
        layer3[29][15:8] = buffer_data_1[2791:2784];
        layer3[29][23:16] = buffer_data_1[2799:2792];
        layer3[29][31:24] = buffer_data_1[2807:2800];
        layer3[29][39:32] = buffer_data_1[2815:2808];
        layer4[29][7:0] = buffer_data_0[2783:2776];
        layer4[29][15:8] = buffer_data_0[2791:2784];
        layer4[29][23:16] = buffer_data_0[2799:2792];
        layer4[29][31:24] = buffer_data_0[2807:2800];
        layer4[29][39:32] = buffer_data_0[2815:2808];
        layer0[30][7:0] = buffer_data_4[2791:2784];
        layer0[30][15:8] = buffer_data_4[2799:2792];
        layer0[30][23:16] = buffer_data_4[2807:2800];
        layer0[30][31:24] = buffer_data_4[2815:2808];
        layer0[30][39:32] = buffer_data_4[2823:2816];
        layer1[30][7:0] = buffer_data_3[2791:2784];
        layer1[30][15:8] = buffer_data_3[2799:2792];
        layer1[30][23:16] = buffer_data_3[2807:2800];
        layer1[30][31:24] = buffer_data_3[2815:2808];
        layer1[30][39:32] = buffer_data_3[2823:2816];
        layer2[30][7:0] = buffer_data_2[2791:2784];
        layer2[30][15:8] = buffer_data_2[2799:2792];
        layer2[30][23:16] = buffer_data_2[2807:2800];
        layer2[30][31:24] = buffer_data_2[2815:2808];
        layer2[30][39:32] = buffer_data_2[2823:2816];
        layer3[30][7:0] = buffer_data_1[2791:2784];
        layer3[30][15:8] = buffer_data_1[2799:2792];
        layer3[30][23:16] = buffer_data_1[2807:2800];
        layer3[30][31:24] = buffer_data_1[2815:2808];
        layer3[30][39:32] = buffer_data_1[2823:2816];
        layer4[30][7:0] = buffer_data_0[2791:2784];
        layer4[30][15:8] = buffer_data_0[2799:2792];
        layer4[30][23:16] = buffer_data_0[2807:2800];
        layer4[30][31:24] = buffer_data_0[2815:2808];
        layer4[30][39:32] = buffer_data_0[2823:2816];
        layer0[31][7:0] = buffer_data_4[2799:2792];
        layer0[31][15:8] = buffer_data_4[2807:2800];
        layer0[31][23:16] = buffer_data_4[2815:2808];
        layer0[31][31:24] = buffer_data_4[2823:2816];
        layer0[31][39:32] = buffer_data_4[2831:2824];
        layer1[31][7:0] = buffer_data_3[2799:2792];
        layer1[31][15:8] = buffer_data_3[2807:2800];
        layer1[31][23:16] = buffer_data_3[2815:2808];
        layer1[31][31:24] = buffer_data_3[2823:2816];
        layer1[31][39:32] = buffer_data_3[2831:2824];
        layer2[31][7:0] = buffer_data_2[2799:2792];
        layer2[31][15:8] = buffer_data_2[2807:2800];
        layer2[31][23:16] = buffer_data_2[2815:2808];
        layer2[31][31:24] = buffer_data_2[2823:2816];
        layer2[31][39:32] = buffer_data_2[2831:2824];
        layer3[31][7:0] = buffer_data_1[2799:2792];
        layer3[31][15:8] = buffer_data_1[2807:2800];
        layer3[31][23:16] = buffer_data_1[2815:2808];
        layer3[31][31:24] = buffer_data_1[2823:2816];
        layer3[31][39:32] = buffer_data_1[2831:2824];
        layer4[31][7:0] = buffer_data_0[2799:2792];
        layer4[31][15:8] = buffer_data_0[2807:2800];
        layer4[31][23:16] = buffer_data_0[2815:2808];
        layer4[31][31:24] = buffer_data_0[2823:2816];
        layer4[31][39:32] = buffer_data_0[2831:2824];
        layer0[32][7:0] = buffer_data_4[2807:2800];
        layer0[32][15:8] = buffer_data_4[2815:2808];
        layer0[32][23:16] = buffer_data_4[2823:2816];
        layer0[32][31:24] = buffer_data_4[2831:2824];
        layer0[32][39:32] = buffer_data_4[2839:2832];
        layer1[32][7:0] = buffer_data_3[2807:2800];
        layer1[32][15:8] = buffer_data_3[2815:2808];
        layer1[32][23:16] = buffer_data_3[2823:2816];
        layer1[32][31:24] = buffer_data_3[2831:2824];
        layer1[32][39:32] = buffer_data_3[2839:2832];
        layer2[32][7:0] = buffer_data_2[2807:2800];
        layer2[32][15:8] = buffer_data_2[2815:2808];
        layer2[32][23:16] = buffer_data_2[2823:2816];
        layer2[32][31:24] = buffer_data_2[2831:2824];
        layer2[32][39:32] = buffer_data_2[2839:2832];
        layer3[32][7:0] = buffer_data_1[2807:2800];
        layer3[32][15:8] = buffer_data_1[2815:2808];
        layer3[32][23:16] = buffer_data_1[2823:2816];
        layer3[32][31:24] = buffer_data_1[2831:2824];
        layer3[32][39:32] = buffer_data_1[2839:2832];
        layer4[32][7:0] = buffer_data_0[2807:2800];
        layer4[32][15:8] = buffer_data_0[2815:2808];
        layer4[32][23:16] = buffer_data_0[2823:2816];
        layer4[32][31:24] = buffer_data_0[2831:2824];
        layer4[32][39:32] = buffer_data_0[2839:2832];
        layer0[33][7:0] = buffer_data_4[2815:2808];
        layer0[33][15:8] = buffer_data_4[2823:2816];
        layer0[33][23:16] = buffer_data_4[2831:2824];
        layer0[33][31:24] = buffer_data_4[2839:2832];
        layer0[33][39:32] = buffer_data_4[2847:2840];
        layer1[33][7:0] = buffer_data_3[2815:2808];
        layer1[33][15:8] = buffer_data_3[2823:2816];
        layer1[33][23:16] = buffer_data_3[2831:2824];
        layer1[33][31:24] = buffer_data_3[2839:2832];
        layer1[33][39:32] = buffer_data_3[2847:2840];
        layer2[33][7:0] = buffer_data_2[2815:2808];
        layer2[33][15:8] = buffer_data_2[2823:2816];
        layer2[33][23:16] = buffer_data_2[2831:2824];
        layer2[33][31:24] = buffer_data_2[2839:2832];
        layer2[33][39:32] = buffer_data_2[2847:2840];
        layer3[33][7:0] = buffer_data_1[2815:2808];
        layer3[33][15:8] = buffer_data_1[2823:2816];
        layer3[33][23:16] = buffer_data_1[2831:2824];
        layer3[33][31:24] = buffer_data_1[2839:2832];
        layer3[33][39:32] = buffer_data_1[2847:2840];
        layer4[33][7:0] = buffer_data_0[2815:2808];
        layer4[33][15:8] = buffer_data_0[2823:2816];
        layer4[33][23:16] = buffer_data_0[2831:2824];
        layer4[33][31:24] = buffer_data_0[2839:2832];
        layer4[33][39:32] = buffer_data_0[2847:2840];
        layer0[34][7:0] = buffer_data_4[2823:2816];
        layer0[34][15:8] = buffer_data_4[2831:2824];
        layer0[34][23:16] = buffer_data_4[2839:2832];
        layer0[34][31:24] = buffer_data_4[2847:2840];
        layer0[34][39:32] = buffer_data_4[2855:2848];
        layer1[34][7:0] = buffer_data_3[2823:2816];
        layer1[34][15:8] = buffer_data_3[2831:2824];
        layer1[34][23:16] = buffer_data_3[2839:2832];
        layer1[34][31:24] = buffer_data_3[2847:2840];
        layer1[34][39:32] = buffer_data_3[2855:2848];
        layer2[34][7:0] = buffer_data_2[2823:2816];
        layer2[34][15:8] = buffer_data_2[2831:2824];
        layer2[34][23:16] = buffer_data_2[2839:2832];
        layer2[34][31:24] = buffer_data_2[2847:2840];
        layer2[34][39:32] = buffer_data_2[2855:2848];
        layer3[34][7:0] = buffer_data_1[2823:2816];
        layer3[34][15:8] = buffer_data_1[2831:2824];
        layer3[34][23:16] = buffer_data_1[2839:2832];
        layer3[34][31:24] = buffer_data_1[2847:2840];
        layer3[34][39:32] = buffer_data_1[2855:2848];
        layer4[34][7:0] = buffer_data_0[2823:2816];
        layer4[34][15:8] = buffer_data_0[2831:2824];
        layer4[34][23:16] = buffer_data_0[2839:2832];
        layer4[34][31:24] = buffer_data_0[2847:2840];
        layer4[34][39:32] = buffer_data_0[2855:2848];
        layer0[35][7:0] = buffer_data_4[2831:2824];
        layer0[35][15:8] = buffer_data_4[2839:2832];
        layer0[35][23:16] = buffer_data_4[2847:2840];
        layer0[35][31:24] = buffer_data_4[2855:2848];
        layer0[35][39:32] = buffer_data_4[2863:2856];
        layer1[35][7:0] = buffer_data_3[2831:2824];
        layer1[35][15:8] = buffer_data_3[2839:2832];
        layer1[35][23:16] = buffer_data_3[2847:2840];
        layer1[35][31:24] = buffer_data_3[2855:2848];
        layer1[35][39:32] = buffer_data_3[2863:2856];
        layer2[35][7:0] = buffer_data_2[2831:2824];
        layer2[35][15:8] = buffer_data_2[2839:2832];
        layer2[35][23:16] = buffer_data_2[2847:2840];
        layer2[35][31:24] = buffer_data_2[2855:2848];
        layer2[35][39:32] = buffer_data_2[2863:2856];
        layer3[35][7:0] = buffer_data_1[2831:2824];
        layer3[35][15:8] = buffer_data_1[2839:2832];
        layer3[35][23:16] = buffer_data_1[2847:2840];
        layer3[35][31:24] = buffer_data_1[2855:2848];
        layer3[35][39:32] = buffer_data_1[2863:2856];
        layer4[35][7:0] = buffer_data_0[2831:2824];
        layer4[35][15:8] = buffer_data_0[2839:2832];
        layer4[35][23:16] = buffer_data_0[2847:2840];
        layer4[35][31:24] = buffer_data_0[2855:2848];
        layer4[35][39:32] = buffer_data_0[2863:2856];
        layer0[36][7:0] = buffer_data_4[2839:2832];
        layer0[36][15:8] = buffer_data_4[2847:2840];
        layer0[36][23:16] = buffer_data_4[2855:2848];
        layer0[36][31:24] = buffer_data_4[2863:2856];
        layer0[36][39:32] = buffer_data_4[2871:2864];
        layer1[36][7:0] = buffer_data_3[2839:2832];
        layer1[36][15:8] = buffer_data_3[2847:2840];
        layer1[36][23:16] = buffer_data_3[2855:2848];
        layer1[36][31:24] = buffer_data_3[2863:2856];
        layer1[36][39:32] = buffer_data_3[2871:2864];
        layer2[36][7:0] = buffer_data_2[2839:2832];
        layer2[36][15:8] = buffer_data_2[2847:2840];
        layer2[36][23:16] = buffer_data_2[2855:2848];
        layer2[36][31:24] = buffer_data_2[2863:2856];
        layer2[36][39:32] = buffer_data_2[2871:2864];
        layer3[36][7:0] = buffer_data_1[2839:2832];
        layer3[36][15:8] = buffer_data_1[2847:2840];
        layer3[36][23:16] = buffer_data_1[2855:2848];
        layer3[36][31:24] = buffer_data_1[2863:2856];
        layer3[36][39:32] = buffer_data_1[2871:2864];
        layer4[36][7:0] = buffer_data_0[2839:2832];
        layer4[36][15:8] = buffer_data_0[2847:2840];
        layer4[36][23:16] = buffer_data_0[2855:2848];
        layer4[36][31:24] = buffer_data_0[2863:2856];
        layer4[36][39:32] = buffer_data_0[2871:2864];
        layer0[37][7:0] = buffer_data_4[2847:2840];
        layer0[37][15:8] = buffer_data_4[2855:2848];
        layer0[37][23:16] = buffer_data_4[2863:2856];
        layer0[37][31:24] = buffer_data_4[2871:2864];
        layer0[37][39:32] = buffer_data_4[2879:2872];
        layer1[37][7:0] = buffer_data_3[2847:2840];
        layer1[37][15:8] = buffer_data_3[2855:2848];
        layer1[37][23:16] = buffer_data_3[2863:2856];
        layer1[37][31:24] = buffer_data_3[2871:2864];
        layer1[37][39:32] = buffer_data_3[2879:2872];
        layer2[37][7:0] = buffer_data_2[2847:2840];
        layer2[37][15:8] = buffer_data_2[2855:2848];
        layer2[37][23:16] = buffer_data_2[2863:2856];
        layer2[37][31:24] = buffer_data_2[2871:2864];
        layer2[37][39:32] = buffer_data_2[2879:2872];
        layer3[37][7:0] = buffer_data_1[2847:2840];
        layer3[37][15:8] = buffer_data_1[2855:2848];
        layer3[37][23:16] = buffer_data_1[2863:2856];
        layer3[37][31:24] = buffer_data_1[2871:2864];
        layer3[37][39:32] = buffer_data_1[2879:2872];
        layer4[37][7:0] = buffer_data_0[2847:2840];
        layer4[37][15:8] = buffer_data_0[2855:2848];
        layer4[37][23:16] = buffer_data_0[2863:2856];
        layer4[37][31:24] = buffer_data_0[2871:2864];
        layer4[37][39:32] = buffer_data_0[2879:2872];
        layer0[38][7:0] = buffer_data_4[2855:2848];
        layer0[38][15:8] = buffer_data_4[2863:2856];
        layer0[38][23:16] = buffer_data_4[2871:2864];
        layer0[38][31:24] = buffer_data_4[2879:2872];
        layer0[38][39:32] = buffer_data_4[2887:2880];
        layer1[38][7:0] = buffer_data_3[2855:2848];
        layer1[38][15:8] = buffer_data_3[2863:2856];
        layer1[38][23:16] = buffer_data_3[2871:2864];
        layer1[38][31:24] = buffer_data_3[2879:2872];
        layer1[38][39:32] = buffer_data_3[2887:2880];
        layer2[38][7:0] = buffer_data_2[2855:2848];
        layer2[38][15:8] = buffer_data_2[2863:2856];
        layer2[38][23:16] = buffer_data_2[2871:2864];
        layer2[38][31:24] = buffer_data_2[2879:2872];
        layer2[38][39:32] = buffer_data_2[2887:2880];
        layer3[38][7:0] = buffer_data_1[2855:2848];
        layer3[38][15:8] = buffer_data_1[2863:2856];
        layer3[38][23:16] = buffer_data_1[2871:2864];
        layer3[38][31:24] = buffer_data_1[2879:2872];
        layer3[38][39:32] = buffer_data_1[2887:2880];
        layer4[38][7:0] = buffer_data_0[2855:2848];
        layer4[38][15:8] = buffer_data_0[2863:2856];
        layer4[38][23:16] = buffer_data_0[2871:2864];
        layer4[38][31:24] = buffer_data_0[2879:2872];
        layer4[38][39:32] = buffer_data_0[2887:2880];
        layer0[39][7:0] = buffer_data_4[2863:2856];
        layer0[39][15:8] = buffer_data_4[2871:2864];
        layer0[39][23:16] = buffer_data_4[2879:2872];
        layer0[39][31:24] = buffer_data_4[2887:2880];
        layer0[39][39:32] = buffer_data_4[2895:2888];
        layer1[39][7:0] = buffer_data_3[2863:2856];
        layer1[39][15:8] = buffer_data_3[2871:2864];
        layer1[39][23:16] = buffer_data_3[2879:2872];
        layer1[39][31:24] = buffer_data_3[2887:2880];
        layer1[39][39:32] = buffer_data_3[2895:2888];
        layer2[39][7:0] = buffer_data_2[2863:2856];
        layer2[39][15:8] = buffer_data_2[2871:2864];
        layer2[39][23:16] = buffer_data_2[2879:2872];
        layer2[39][31:24] = buffer_data_2[2887:2880];
        layer2[39][39:32] = buffer_data_2[2895:2888];
        layer3[39][7:0] = buffer_data_1[2863:2856];
        layer3[39][15:8] = buffer_data_1[2871:2864];
        layer3[39][23:16] = buffer_data_1[2879:2872];
        layer3[39][31:24] = buffer_data_1[2887:2880];
        layer3[39][39:32] = buffer_data_1[2895:2888];
        layer4[39][7:0] = buffer_data_0[2863:2856];
        layer4[39][15:8] = buffer_data_0[2871:2864];
        layer4[39][23:16] = buffer_data_0[2879:2872];
        layer4[39][31:24] = buffer_data_0[2887:2880];
        layer4[39][39:32] = buffer_data_0[2895:2888];
        layer0[40][7:0] = buffer_data_4[2871:2864];
        layer0[40][15:8] = buffer_data_4[2879:2872];
        layer0[40][23:16] = buffer_data_4[2887:2880];
        layer0[40][31:24] = buffer_data_4[2895:2888];
        layer0[40][39:32] = buffer_data_4[2903:2896];
        layer1[40][7:0] = buffer_data_3[2871:2864];
        layer1[40][15:8] = buffer_data_3[2879:2872];
        layer1[40][23:16] = buffer_data_3[2887:2880];
        layer1[40][31:24] = buffer_data_3[2895:2888];
        layer1[40][39:32] = buffer_data_3[2903:2896];
        layer2[40][7:0] = buffer_data_2[2871:2864];
        layer2[40][15:8] = buffer_data_2[2879:2872];
        layer2[40][23:16] = buffer_data_2[2887:2880];
        layer2[40][31:24] = buffer_data_2[2895:2888];
        layer2[40][39:32] = buffer_data_2[2903:2896];
        layer3[40][7:0] = buffer_data_1[2871:2864];
        layer3[40][15:8] = buffer_data_1[2879:2872];
        layer3[40][23:16] = buffer_data_1[2887:2880];
        layer3[40][31:24] = buffer_data_1[2895:2888];
        layer3[40][39:32] = buffer_data_1[2903:2896];
        layer4[40][7:0] = buffer_data_0[2871:2864];
        layer4[40][15:8] = buffer_data_0[2879:2872];
        layer4[40][23:16] = buffer_data_0[2887:2880];
        layer4[40][31:24] = buffer_data_0[2895:2888];
        layer4[40][39:32] = buffer_data_0[2903:2896];
        layer0[41][7:0] = buffer_data_4[2879:2872];
        layer0[41][15:8] = buffer_data_4[2887:2880];
        layer0[41][23:16] = buffer_data_4[2895:2888];
        layer0[41][31:24] = buffer_data_4[2903:2896];
        layer0[41][39:32] = buffer_data_4[2911:2904];
        layer1[41][7:0] = buffer_data_3[2879:2872];
        layer1[41][15:8] = buffer_data_3[2887:2880];
        layer1[41][23:16] = buffer_data_3[2895:2888];
        layer1[41][31:24] = buffer_data_3[2903:2896];
        layer1[41][39:32] = buffer_data_3[2911:2904];
        layer2[41][7:0] = buffer_data_2[2879:2872];
        layer2[41][15:8] = buffer_data_2[2887:2880];
        layer2[41][23:16] = buffer_data_2[2895:2888];
        layer2[41][31:24] = buffer_data_2[2903:2896];
        layer2[41][39:32] = buffer_data_2[2911:2904];
        layer3[41][7:0] = buffer_data_1[2879:2872];
        layer3[41][15:8] = buffer_data_1[2887:2880];
        layer3[41][23:16] = buffer_data_1[2895:2888];
        layer3[41][31:24] = buffer_data_1[2903:2896];
        layer3[41][39:32] = buffer_data_1[2911:2904];
        layer4[41][7:0] = buffer_data_0[2879:2872];
        layer4[41][15:8] = buffer_data_0[2887:2880];
        layer4[41][23:16] = buffer_data_0[2895:2888];
        layer4[41][31:24] = buffer_data_0[2903:2896];
        layer4[41][39:32] = buffer_data_0[2911:2904];
        layer0[42][7:0] = buffer_data_4[2887:2880];
        layer0[42][15:8] = buffer_data_4[2895:2888];
        layer0[42][23:16] = buffer_data_4[2903:2896];
        layer0[42][31:24] = buffer_data_4[2911:2904];
        layer0[42][39:32] = buffer_data_4[2919:2912];
        layer1[42][7:0] = buffer_data_3[2887:2880];
        layer1[42][15:8] = buffer_data_3[2895:2888];
        layer1[42][23:16] = buffer_data_3[2903:2896];
        layer1[42][31:24] = buffer_data_3[2911:2904];
        layer1[42][39:32] = buffer_data_3[2919:2912];
        layer2[42][7:0] = buffer_data_2[2887:2880];
        layer2[42][15:8] = buffer_data_2[2895:2888];
        layer2[42][23:16] = buffer_data_2[2903:2896];
        layer2[42][31:24] = buffer_data_2[2911:2904];
        layer2[42][39:32] = buffer_data_2[2919:2912];
        layer3[42][7:0] = buffer_data_1[2887:2880];
        layer3[42][15:8] = buffer_data_1[2895:2888];
        layer3[42][23:16] = buffer_data_1[2903:2896];
        layer3[42][31:24] = buffer_data_1[2911:2904];
        layer3[42][39:32] = buffer_data_1[2919:2912];
        layer4[42][7:0] = buffer_data_0[2887:2880];
        layer4[42][15:8] = buffer_data_0[2895:2888];
        layer4[42][23:16] = buffer_data_0[2903:2896];
        layer4[42][31:24] = buffer_data_0[2911:2904];
        layer4[42][39:32] = buffer_data_0[2919:2912];
        layer0[43][7:0] = buffer_data_4[2895:2888];
        layer0[43][15:8] = buffer_data_4[2903:2896];
        layer0[43][23:16] = buffer_data_4[2911:2904];
        layer0[43][31:24] = buffer_data_4[2919:2912];
        layer0[43][39:32] = buffer_data_4[2927:2920];
        layer1[43][7:0] = buffer_data_3[2895:2888];
        layer1[43][15:8] = buffer_data_3[2903:2896];
        layer1[43][23:16] = buffer_data_3[2911:2904];
        layer1[43][31:24] = buffer_data_3[2919:2912];
        layer1[43][39:32] = buffer_data_3[2927:2920];
        layer2[43][7:0] = buffer_data_2[2895:2888];
        layer2[43][15:8] = buffer_data_2[2903:2896];
        layer2[43][23:16] = buffer_data_2[2911:2904];
        layer2[43][31:24] = buffer_data_2[2919:2912];
        layer2[43][39:32] = buffer_data_2[2927:2920];
        layer3[43][7:0] = buffer_data_1[2895:2888];
        layer3[43][15:8] = buffer_data_1[2903:2896];
        layer3[43][23:16] = buffer_data_1[2911:2904];
        layer3[43][31:24] = buffer_data_1[2919:2912];
        layer3[43][39:32] = buffer_data_1[2927:2920];
        layer4[43][7:0] = buffer_data_0[2895:2888];
        layer4[43][15:8] = buffer_data_0[2903:2896];
        layer4[43][23:16] = buffer_data_0[2911:2904];
        layer4[43][31:24] = buffer_data_0[2919:2912];
        layer4[43][39:32] = buffer_data_0[2927:2920];
        layer0[44][7:0] = buffer_data_4[2903:2896];
        layer0[44][15:8] = buffer_data_4[2911:2904];
        layer0[44][23:16] = buffer_data_4[2919:2912];
        layer0[44][31:24] = buffer_data_4[2927:2920];
        layer0[44][39:32] = buffer_data_4[2935:2928];
        layer1[44][7:0] = buffer_data_3[2903:2896];
        layer1[44][15:8] = buffer_data_3[2911:2904];
        layer1[44][23:16] = buffer_data_3[2919:2912];
        layer1[44][31:24] = buffer_data_3[2927:2920];
        layer1[44][39:32] = buffer_data_3[2935:2928];
        layer2[44][7:0] = buffer_data_2[2903:2896];
        layer2[44][15:8] = buffer_data_2[2911:2904];
        layer2[44][23:16] = buffer_data_2[2919:2912];
        layer2[44][31:24] = buffer_data_2[2927:2920];
        layer2[44][39:32] = buffer_data_2[2935:2928];
        layer3[44][7:0] = buffer_data_1[2903:2896];
        layer3[44][15:8] = buffer_data_1[2911:2904];
        layer3[44][23:16] = buffer_data_1[2919:2912];
        layer3[44][31:24] = buffer_data_1[2927:2920];
        layer3[44][39:32] = buffer_data_1[2935:2928];
        layer4[44][7:0] = buffer_data_0[2903:2896];
        layer4[44][15:8] = buffer_data_0[2911:2904];
        layer4[44][23:16] = buffer_data_0[2919:2912];
        layer4[44][31:24] = buffer_data_0[2927:2920];
        layer4[44][39:32] = buffer_data_0[2935:2928];
        layer0[45][7:0] = buffer_data_4[2911:2904];
        layer0[45][15:8] = buffer_data_4[2919:2912];
        layer0[45][23:16] = buffer_data_4[2927:2920];
        layer0[45][31:24] = buffer_data_4[2935:2928];
        layer0[45][39:32] = buffer_data_4[2943:2936];
        layer1[45][7:0] = buffer_data_3[2911:2904];
        layer1[45][15:8] = buffer_data_3[2919:2912];
        layer1[45][23:16] = buffer_data_3[2927:2920];
        layer1[45][31:24] = buffer_data_3[2935:2928];
        layer1[45][39:32] = buffer_data_3[2943:2936];
        layer2[45][7:0] = buffer_data_2[2911:2904];
        layer2[45][15:8] = buffer_data_2[2919:2912];
        layer2[45][23:16] = buffer_data_2[2927:2920];
        layer2[45][31:24] = buffer_data_2[2935:2928];
        layer2[45][39:32] = buffer_data_2[2943:2936];
        layer3[45][7:0] = buffer_data_1[2911:2904];
        layer3[45][15:8] = buffer_data_1[2919:2912];
        layer3[45][23:16] = buffer_data_1[2927:2920];
        layer3[45][31:24] = buffer_data_1[2935:2928];
        layer3[45][39:32] = buffer_data_1[2943:2936];
        layer4[45][7:0] = buffer_data_0[2911:2904];
        layer4[45][15:8] = buffer_data_0[2919:2912];
        layer4[45][23:16] = buffer_data_0[2927:2920];
        layer4[45][31:24] = buffer_data_0[2935:2928];
        layer4[45][39:32] = buffer_data_0[2943:2936];
        layer0[46][7:0] = buffer_data_4[2919:2912];
        layer0[46][15:8] = buffer_data_4[2927:2920];
        layer0[46][23:16] = buffer_data_4[2935:2928];
        layer0[46][31:24] = buffer_data_4[2943:2936];
        layer0[46][39:32] = buffer_data_4[2951:2944];
        layer1[46][7:0] = buffer_data_3[2919:2912];
        layer1[46][15:8] = buffer_data_3[2927:2920];
        layer1[46][23:16] = buffer_data_3[2935:2928];
        layer1[46][31:24] = buffer_data_3[2943:2936];
        layer1[46][39:32] = buffer_data_3[2951:2944];
        layer2[46][7:0] = buffer_data_2[2919:2912];
        layer2[46][15:8] = buffer_data_2[2927:2920];
        layer2[46][23:16] = buffer_data_2[2935:2928];
        layer2[46][31:24] = buffer_data_2[2943:2936];
        layer2[46][39:32] = buffer_data_2[2951:2944];
        layer3[46][7:0] = buffer_data_1[2919:2912];
        layer3[46][15:8] = buffer_data_1[2927:2920];
        layer3[46][23:16] = buffer_data_1[2935:2928];
        layer3[46][31:24] = buffer_data_1[2943:2936];
        layer3[46][39:32] = buffer_data_1[2951:2944];
        layer4[46][7:0] = buffer_data_0[2919:2912];
        layer4[46][15:8] = buffer_data_0[2927:2920];
        layer4[46][23:16] = buffer_data_0[2935:2928];
        layer4[46][31:24] = buffer_data_0[2943:2936];
        layer4[46][39:32] = buffer_data_0[2951:2944];
        layer0[47][7:0] = buffer_data_4[2927:2920];
        layer0[47][15:8] = buffer_data_4[2935:2928];
        layer0[47][23:16] = buffer_data_4[2943:2936];
        layer0[47][31:24] = buffer_data_4[2951:2944];
        layer0[47][39:32] = buffer_data_4[2959:2952];
        layer1[47][7:0] = buffer_data_3[2927:2920];
        layer1[47][15:8] = buffer_data_3[2935:2928];
        layer1[47][23:16] = buffer_data_3[2943:2936];
        layer1[47][31:24] = buffer_data_3[2951:2944];
        layer1[47][39:32] = buffer_data_3[2959:2952];
        layer2[47][7:0] = buffer_data_2[2927:2920];
        layer2[47][15:8] = buffer_data_2[2935:2928];
        layer2[47][23:16] = buffer_data_2[2943:2936];
        layer2[47][31:24] = buffer_data_2[2951:2944];
        layer2[47][39:32] = buffer_data_2[2959:2952];
        layer3[47][7:0] = buffer_data_1[2927:2920];
        layer3[47][15:8] = buffer_data_1[2935:2928];
        layer3[47][23:16] = buffer_data_1[2943:2936];
        layer3[47][31:24] = buffer_data_1[2951:2944];
        layer3[47][39:32] = buffer_data_1[2959:2952];
        layer4[47][7:0] = buffer_data_0[2927:2920];
        layer4[47][15:8] = buffer_data_0[2935:2928];
        layer4[47][23:16] = buffer_data_0[2943:2936];
        layer4[47][31:24] = buffer_data_0[2951:2944];
        layer4[47][39:32] = buffer_data_0[2959:2952];
        layer0[48][7:0] = buffer_data_4[2935:2928];
        layer0[48][15:8] = buffer_data_4[2943:2936];
        layer0[48][23:16] = buffer_data_4[2951:2944];
        layer0[48][31:24] = buffer_data_4[2959:2952];
        layer0[48][39:32] = buffer_data_4[2967:2960];
        layer1[48][7:0] = buffer_data_3[2935:2928];
        layer1[48][15:8] = buffer_data_3[2943:2936];
        layer1[48][23:16] = buffer_data_3[2951:2944];
        layer1[48][31:24] = buffer_data_3[2959:2952];
        layer1[48][39:32] = buffer_data_3[2967:2960];
        layer2[48][7:0] = buffer_data_2[2935:2928];
        layer2[48][15:8] = buffer_data_2[2943:2936];
        layer2[48][23:16] = buffer_data_2[2951:2944];
        layer2[48][31:24] = buffer_data_2[2959:2952];
        layer2[48][39:32] = buffer_data_2[2967:2960];
        layer3[48][7:0] = buffer_data_1[2935:2928];
        layer3[48][15:8] = buffer_data_1[2943:2936];
        layer3[48][23:16] = buffer_data_1[2951:2944];
        layer3[48][31:24] = buffer_data_1[2959:2952];
        layer3[48][39:32] = buffer_data_1[2967:2960];
        layer4[48][7:0] = buffer_data_0[2935:2928];
        layer4[48][15:8] = buffer_data_0[2943:2936];
        layer4[48][23:16] = buffer_data_0[2951:2944];
        layer4[48][31:24] = buffer_data_0[2959:2952];
        layer4[48][39:32] = buffer_data_0[2967:2960];
        layer0[49][7:0] = buffer_data_4[2943:2936];
        layer0[49][15:8] = buffer_data_4[2951:2944];
        layer0[49][23:16] = buffer_data_4[2959:2952];
        layer0[49][31:24] = buffer_data_4[2967:2960];
        layer0[49][39:32] = buffer_data_4[2975:2968];
        layer1[49][7:0] = buffer_data_3[2943:2936];
        layer1[49][15:8] = buffer_data_3[2951:2944];
        layer1[49][23:16] = buffer_data_3[2959:2952];
        layer1[49][31:24] = buffer_data_3[2967:2960];
        layer1[49][39:32] = buffer_data_3[2975:2968];
        layer2[49][7:0] = buffer_data_2[2943:2936];
        layer2[49][15:8] = buffer_data_2[2951:2944];
        layer2[49][23:16] = buffer_data_2[2959:2952];
        layer2[49][31:24] = buffer_data_2[2967:2960];
        layer2[49][39:32] = buffer_data_2[2975:2968];
        layer3[49][7:0] = buffer_data_1[2943:2936];
        layer3[49][15:8] = buffer_data_1[2951:2944];
        layer3[49][23:16] = buffer_data_1[2959:2952];
        layer3[49][31:24] = buffer_data_1[2967:2960];
        layer3[49][39:32] = buffer_data_1[2975:2968];
        layer4[49][7:0] = buffer_data_0[2943:2936];
        layer4[49][15:8] = buffer_data_0[2951:2944];
        layer4[49][23:16] = buffer_data_0[2959:2952];
        layer4[49][31:24] = buffer_data_0[2967:2960];
        layer4[49][39:32] = buffer_data_0[2975:2968];
        layer0[50][7:0] = buffer_data_4[2951:2944];
        layer0[50][15:8] = buffer_data_4[2959:2952];
        layer0[50][23:16] = buffer_data_4[2967:2960];
        layer0[50][31:24] = buffer_data_4[2975:2968];
        layer0[50][39:32] = buffer_data_4[2983:2976];
        layer1[50][7:0] = buffer_data_3[2951:2944];
        layer1[50][15:8] = buffer_data_3[2959:2952];
        layer1[50][23:16] = buffer_data_3[2967:2960];
        layer1[50][31:24] = buffer_data_3[2975:2968];
        layer1[50][39:32] = buffer_data_3[2983:2976];
        layer2[50][7:0] = buffer_data_2[2951:2944];
        layer2[50][15:8] = buffer_data_2[2959:2952];
        layer2[50][23:16] = buffer_data_2[2967:2960];
        layer2[50][31:24] = buffer_data_2[2975:2968];
        layer2[50][39:32] = buffer_data_2[2983:2976];
        layer3[50][7:0] = buffer_data_1[2951:2944];
        layer3[50][15:8] = buffer_data_1[2959:2952];
        layer3[50][23:16] = buffer_data_1[2967:2960];
        layer3[50][31:24] = buffer_data_1[2975:2968];
        layer3[50][39:32] = buffer_data_1[2983:2976];
        layer4[50][7:0] = buffer_data_0[2951:2944];
        layer4[50][15:8] = buffer_data_0[2959:2952];
        layer4[50][23:16] = buffer_data_0[2967:2960];
        layer4[50][31:24] = buffer_data_0[2975:2968];
        layer4[50][39:32] = buffer_data_0[2983:2976];
        layer0[51][7:0] = buffer_data_4[2959:2952];
        layer0[51][15:8] = buffer_data_4[2967:2960];
        layer0[51][23:16] = buffer_data_4[2975:2968];
        layer0[51][31:24] = buffer_data_4[2983:2976];
        layer0[51][39:32] = buffer_data_4[2991:2984];
        layer1[51][7:0] = buffer_data_3[2959:2952];
        layer1[51][15:8] = buffer_data_3[2967:2960];
        layer1[51][23:16] = buffer_data_3[2975:2968];
        layer1[51][31:24] = buffer_data_3[2983:2976];
        layer1[51][39:32] = buffer_data_3[2991:2984];
        layer2[51][7:0] = buffer_data_2[2959:2952];
        layer2[51][15:8] = buffer_data_2[2967:2960];
        layer2[51][23:16] = buffer_data_2[2975:2968];
        layer2[51][31:24] = buffer_data_2[2983:2976];
        layer2[51][39:32] = buffer_data_2[2991:2984];
        layer3[51][7:0] = buffer_data_1[2959:2952];
        layer3[51][15:8] = buffer_data_1[2967:2960];
        layer3[51][23:16] = buffer_data_1[2975:2968];
        layer3[51][31:24] = buffer_data_1[2983:2976];
        layer3[51][39:32] = buffer_data_1[2991:2984];
        layer4[51][7:0] = buffer_data_0[2959:2952];
        layer4[51][15:8] = buffer_data_0[2967:2960];
        layer4[51][23:16] = buffer_data_0[2975:2968];
        layer4[51][31:24] = buffer_data_0[2983:2976];
        layer4[51][39:32] = buffer_data_0[2991:2984];
        layer0[52][7:0] = buffer_data_4[2967:2960];
        layer0[52][15:8] = buffer_data_4[2975:2968];
        layer0[52][23:16] = buffer_data_4[2983:2976];
        layer0[52][31:24] = buffer_data_4[2991:2984];
        layer0[52][39:32] = buffer_data_4[2999:2992];
        layer1[52][7:0] = buffer_data_3[2967:2960];
        layer1[52][15:8] = buffer_data_3[2975:2968];
        layer1[52][23:16] = buffer_data_3[2983:2976];
        layer1[52][31:24] = buffer_data_3[2991:2984];
        layer1[52][39:32] = buffer_data_3[2999:2992];
        layer2[52][7:0] = buffer_data_2[2967:2960];
        layer2[52][15:8] = buffer_data_2[2975:2968];
        layer2[52][23:16] = buffer_data_2[2983:2976];
        layer2[52][31:24] = buffer_data_2[2991:2984];
        layer2[52][39:32] = buffer_data_2[2999:2992];
        layer3[52][7:0] = buffer_data_1[2967:2960];
        layer3[52][15:8] = buffer_data_1[2975:2968];
        layer3[52][23:16] = buffer_data_1[2983:2976];
        layer3[52][31:24] = buffer_data_1[2991:2984];
        layer3[52][39:32] = buffer_data_1[2999:2992];
        layer4[52][7:0] = buffer_data_0[2967:2960];
        layer4[52][15:8] = buffer_data_0[2975:2968];
        layer4[52][23:16] = buffer_data_0[2983:2976];
        layer4[52][31:24] = buffer_data_0[2991:2984];
        layer4[52][39:32] = buffer_data_0[2999:2992];
        layer0[53][7:0] = buffer_data_4[2975:2968];
        layer0[53][15:8] = buffer_data_4[2983:2976];
        layer0[53][23:16] = buffer_data_4[2991:2984];
        layer0[53][31:24] = buffer_data_4[2999:2992];
        layer0[53][39:32] = buffer_data_4[3007:3000];
        layer1[53][7:0] = buffer_data_3[2975:2968];
        layer1[53][15:8] = buffer_data_3[2983:2976];
        layer1[53][23:16] = buffer_data_3[2991:2984];
        layer1[53][31:24] = buffer_data_3[2999:2992];
        layer1[53][39:32] = buffer_data_3[3007:3000];
        layer2[53][7:0] = buffer_data_2[2975:2968];
        layer2[53][15:8] = buffer_data_2[2983:2976];
        layer2[53][23:16] = buffer_data_2[2991:2984];
        layer2[53][31:24] = buffer_data_2[2999:2992];
        layer2[53][39:32] = buffer_data_2[3007:3000];
        layer3[53][7:0] = buffer_data_1[2975:2968];
        layer3[53][15:8] = buffer_data_1[2983:2976];
        layer3[53][23:16] = buffer_data_1[2991:2984];
        layer3[53][31:24] = buffer_data_1[2999:2992];
        layer3[53][39:32] = buffer_data_1[3007:3000];
        layer4[53][7:0] = buffer_data_0[2975:2968];
        layer4[53][15:8] = buffer_data_0[2983:2976];
        layer4[53][23:16] = buffer_data_0[2991:2984];
        layer4[53][31:24] = buffer_data_0[2999:2992];
        layer4[53][39:32] = buffer_data_0[3007:3000];
        layer0[54][7:0] = buffer_data_4[2983:2976];
        layer0[54][15:8] = buffer_data_4[2991:2984];
        layer0[54][23:16] = buffer_data_4[2999:2992];
        layer0[54][31:24] = buffer_data_4[3007:3000];
        layer0[54][39:32] = buffer_data_4[3015:3008];
        layer1[54][7:0] = buffer_data_3[2983:2976];
        layer1[54][15:8] = buffer_data_3[2991:2984];
        layer1[54][23:16] = buffer_data_3[2999:2992];
        layer1[54][31:24] = buffer_data_3[3007:3000];
        layer1[54][39:32] = buffer_data_3[3015:3008];
        layer2[54][7:0] = buffer_data_2[2983:2976];
        layer2[54][15:8] = buffer_data_2[2991:2984];
        layer2[54][23:16] = buffer_data_2[2999:2992];
        layer2[54][31:24] = buffer_data_2[3007:3000];
        layer2[54][39:32] = buffer_data_2[3015:3008];
        layer3[54][7:0] = buffer_data_1[2983:2976];
        layer3[54][15:8] = buffer_data_1[2991:2984];
        layer3[54][23:16] = buffer_data_1[2999:2992];
        layer3[54][31:24] = buffer_data_1[3007:3000];
        layer3[54][39:32] = buffer_data_1[3015:3008];
        layer4[54][7:0] = buffer_data_0[2983:2976];
        layer4[54][15:8] = buffer_data_0[2991:2984];
        layer4[54][23:16] = buffer_data_0[2999:2992];
        layer4[54][31:24] = buffer_data_0[3007:3000];
        layer4[54][39:32] = buffer_data_0[3015:3008];
        layer0[55][7:0] = buffer_data_4[2991:2984];
        layer0[55][15:8] = buffer_data_4[2999:2992];
        layer0[55][23:16] = buffer_data_4[3007:3000];
        layer0[55][31:24] = buffer_data_4[3015:3008];
        layer0[55][39:32] = buffer_data_4[3023:3016];
        layer1[55][7:0] = buffer_data_3[2991:2984];
        layer1[55][15:8] = buffer_data_3[2999:2992];
        layer1[55][23:16] = buffer_data_3[3007:3000];
        layer1[55][31:24] = buffer_data_3[3015:3008];
        layer1[55][39:32] = buffer_data_3[3023:3016];
        layer2[55][7:0] = buffer_data_2[2991:2984];
        layer2[55][15:8] = buffer_data_2[2999:2992];
        layer2[55][23:16] = buffer_data_2[3007:3000];
        layer2[55][31:24] = buffer_data_2[3015:3008];
        layer2[55][39:32] = buffer_data_2[3023:3016];
        layer3[55][7:0] = buffer_data_1[2991:2984];
        layer3[55][15:8] = buffer_data_1[2999:2992];
        layer3[55][23:16] = buffer_data_1[3007:3000];
        layer3[55][31:24] = buffer_data_1[3015:3008];
        layer3[55][39:32] = buffer_data_1[3023:3016];
        layer4[55][7:0] = buffer_data_0[2991:2984];
        layer4[55][15:8] = buffer_data_0[2999:2992];
        layer4[55][23:16] = buffer_data_0[3007:3000];
        layer4[55][31:24] = buffer_data_0[3015:3008];
        layer4[55][39:32] = buffer_data_0[3023:3016];
        layer0[56][7:0] = buffer_data_4[2999:2992];
        layer0[56][15:8] = buffer_data_4[3007:3000];
        layer0[56][23:16] = buffer_data_4[3015:3008];
        layer0[56][31:24] = buffer_data_4[3023:3016];
        layer0[56][39:32] = buffer_data_4[3031:3024];
        layer1[56][7:0] = buffer_data_3[2999:2992];
        layer1[56][15:8] = buffer_data_3[3007:3000];
        layer1[56][23:16] = buffer_data_3[3015:3008];
        layer1[56][31:24] = buffer_data_3[3023:3016];
        layer1[56][39:32] = buffer_data_3[3031:3024];
        layer2[56][7:0] = buffer_data_2[2999:2992];
        layer2[56][15:8] = buffer_data_2[3007:3000];
        layer2[56][23:16] = buffer_data_2[3015:3008];
        layer2[56][31:24] = buffer_data_2[3023:3016];
        layer2[56][39:32] = buffer_data_2[3031:3024];
        layer3[56][7:0] = buffer_data_1[2999:2992];
        layer3[56][15:8] = buffer_data_1[3007:3000];
        layer3[56][23:16] = buffer_data_1[3015:3008];
        layer3[56][31:24] = buffer_data_1[3023:3016];
        layer3[56][39:32] = buffer_data_1[3031:3024];
        layer4[56][7:0] = buffer_data_0[2999:2992];
        layer4[56][15:8] = buffer_data_0[3007:3000];
        layer4[56][23:16] = buffer_data_0[3015:3008];
        layer4[56][31:24] = buffer_data_0[3023:3016];
        layer4[56][39:32] = buffer_data_0[3031:3024];
        layer0[57][7:0] = buffer_data_4[3007:3000];
        layer0[57][15:8] = buffer_data_4[3015:3008];
        layer0[57][23:16] = buffer_data_4[3023:3016];
        layer0[57][31:24] = buffer_data_4[3031:3024];
        layer0[57][39:32] = buffer_data_4[3039:3032];
        layer1[57][7:0] = buffer_data_3[3007:3000];
        layer1[57][15:8] = buffer_data_3[3015:3008];
        layer1[57][23:16] = buffer_data_3[3023:3016];
        layer1[57][31:24] = buffer_data_3[3031:3024];
        layer1[57][39:32] = buffer_data_3[3039:3032];
        layer2[57][7:0] = buffer_data_2[3007:3000];
        layer2[57][15:8] = buffer_data_2[3015:3008];
        layer2[57][23:16] = buffer_data_2[3023:3016];
        layer2[57][31:24] = buffer_data_2[3031:3024];
        layer2[57][39:32] = buffer_data_2[3039:3032];
        layer3[57][7:0] = buffer_data_1[3007:3000];
        layer3[57][15:8] = buffer_data_1[3015:3008];
        layer3[57][23:16] = buffer_data_1[3023:3016];
        layer3[57][31:24] = buffer_data_1[3031:3024];
        layer3[57][39:32] = buffer_data_1[3039:3032];
        layer4[57][7:0] = buffer_data_0[3007:3000];
        layer4[57][15:8] = buffer_data_0[3015:3008];
        layer4[57][23:16] = buffer_data_0[3023:3016];
        layer4[57][31:24] = buffer_data_0[3031:3024];
        layer4[57][39:32] = buffer_data_0[3039:3032];
        layer0[58][7:0] = buffer_data_4[3015:3008];
        layer0[58][15:8] = buffer_data_4[3023:3016];
        layer0[58][23:16] = buffer_data_4[3031:3024];
        layer0[58][31:24] = buffer_data_4[3039:3032];
        layer0[58][39:32] = buffer_data_4[3047:3040];
        layer1[58][7:0] = buffer_data_3[3015:3008];
        layer1[58][15:8] = buffer_data_3[3023:3016];
        layer1[58][23:16] = buffer_data_3[3031:3024];
        layer1[58][31:24] = buffer_data_3[3039:3032];
        layer1[58][39:32] = buffer_data_3[3047:3040];
        layer2[58][7:0] = buffer_data_2[3015:3008];
        layer2[58][15:8] = buffer_data_2[3023:3016];
        layer2[58][23:16] = buffer_data_2[3031:3024];
        layer2[58][31:24] = buffer_data_2[3039:3032];
        layer2[58][39:32] = buffer_data_2[3047:3040];
        layer3[58][7:0] = buffer_data_1[3015:3008];
        layer3[58][15:8] = buffer_data_1[3023:3016];
        layer3[58][23:16] = buffer_data_1[3031:3024];
        layer3[58][31:24] = buffer_data_1[3039:3032];
        layer3[58][39:32] = buffer_data_1[3047:3040];
        layer4[58][7:0] = buffer_data_0[3015:3008];
        layer4[58][15:8] = buffer_data_0[3023:3016];
        layer4[58][23:16] = buffer_data_0[3031:3024];
        layer4[58][31:24] = buffer_data_0[3039:3032];
        layer4[58][39:32] = buffer_data_0[3047:3040];
        layer0[59][7:0] = buffer_data_4[3023:3016];
        layer0[59][15:8] = buffer_data_4[3031:3024];
        layer0[59][23:16] = buffer_data_4[3039:3032];
        layer0[59][31:24] = buffer_data_4[3047:3040];
        layer0[59][39:32] = buffer_data_4[3055:3048];
        layer1[59][7:0] = buffer_data_3[3023:3016];
        layer1[59][15:8] = buffer_data_3[3031:3024];
        layer1[59][23:16] = buffer_data_3[3039:3032];
        layer1[59][31:24] = buffer_data_3[3047:3040];
        layer1[59][39:32] = buffer_data_3[3055:3048];
        layer2[59][7:0] = buffer_data_2[3023:3016];
        layer2[59][15:8] = buffer_data_2[3031:3024];
        layer2[59][23:16] = buffer_data_2[3039:3032];
        layer2[59][31:24] = buffer_data_2[3047:3040];
        layer2[59][39:32] = buffer_data_2[3055:3048];
        layer3[59][7:0] = buffer_data_1[3023:3016];
        layer3[59][15:8] = buffer_data_1[3031:3024];
        layer3[59][23:16] = buffer_data_1[3039:3032];
        layer3[59][31:24] = buffer_data_1[3047:3040];
        layer3[59][39:32] = buffer_data_1[3055:3048];
        layer4[59][7:0] = buffer_data_0[3023:3016];
        layer4[59][15:8] = buffer_data_0[3031:3024];
        layer4[59][23:16] = buffer_data_0[3039:3032];
        layer4[59][31:24] = buffer_data_0[3047:3040];
        layer4[59][39:32] = buffer_data_0[3055:3048];
        layer0[60][7:0] = buffer_data_4[3031:3024];
        layer0[60][15:8] = buffer_data_4[3039:3032];
        layer0[60][23:16] = buffer_data_4[3047:3040];
        layer0[60][31:24] = buffer_data_4[3055:3048];
        layer0[60][39:32] = buffer_data_4[3063:3056];
        layer1[60][7:0] = buffer_data_3[3031:3024];
        layer1[60][15:8] = buffer_data_3[3039:3032];
        layer1[60][23:16] = buffer_data_3[3047:3040];
        layer1[60][31:24] = buffer_data_3[3055:3048];
        layer1[60][39:32] = buffer_data_3[3063:3056];
        layer2[60][7:0] = buffer_data_2[3031:3024];
        layer2[60][15:8] = buffer_data_2[3039:3032];
        layer2[60][23:16] = buffer_data_2[3047:3040];
        layer2[60][31:24] = buffer_data_2[3055:3048];
        layer2[60][39:32] = buffer_data_2[3063:3056];
        layer3[60][7:0] = buffer_data_1[3031:3024];
        layer3[60][15:8] = buffer_data_1[3039:3032];
        layer3[60][23:16] = buffer_data_1[3047:3040];
        layer3[60][31:24] = buffer_data_1[3055:3048];
        layer3[60][39:32] = buffer_data_1[3063:3056];
        layer4[60][7:0] = buffer_data_0[3031:3024];
        layer4[60][15:8] = buffer_data_0[3039:3032];
        layer4[60][23:16] = buffer_data_0[3047:3040];
        layer4[60][31:24] = buffer_data_0[3055:3048];
        layer4[60][39:32] = buffer_data_0[3063:3056];
        layer0[61][7:0] = buffer_data_4[3039:3032];
        layer0[61][15:8] = buffer_data_4[3047:3040];
        layer0[61][23:16] = buffer_data_4[3055:3048];
        layer0[61][31:24] = buffer_data_4[3063:3056];
        layer0[61][39:32] = buffer_data_4[3071:3064];
        layer1[61][7:0] = buffer_data_3[3039:3032];
        layer1[61][15:8] = buffer_data_3[3047:3040];
        layer1[61][23:16] = buffer_data_3[3055:3048];
        layer1[61][31:24] = buffer_data_3[3063:3056];
        layer1[61][39:32] = buffer_data_3[3071:3064];
        layer2[61][7:0] = buffer_data_2[3039:3032];
        layer2[61][15:8] = buffer_data_2[3047:3040];
        layer2[61][23:16] = buffer_data_2[3055:3048];
        layer2[61][31:24] = buffer_data_2[3063:3056];
        layer2[61][39:32] = buffer_data_2[3071:3064];
        layer3[61][7:0] = buffer_data_1[3039:3032];
        layer3[61][15:8] = buffer_data_1[3047:3040];
        layer3[61][23:16] = buffer_data_1[3055:3048];
        layer3[61][31:24] = buffer_data_1[3063:3056];
        layer3[61][39:32] = buffer_data_1[3071:3064];
        layer4[61][7:0] = buffer_data_0[3039:3032];
        layer4[61][15:8] = buffer_data_0[3047:3040];
        layer4[61][23:16] = buffer_data_0[3055:3048];
        layer4[61][31:24] = buffer_data_0[3063:3056];
        layer4[61][39:32] = buffer_data_0[3071:3064];
        layer0[62][7:0] = buffer_data_4[3047:3040];
        layer0[62][15:8] = buffer_data_4[3055:3048];
        layer0[62][23:16] = buffer_data_4[3063:3056];
        layer0[62][31:24] = buffer_data_4[3071:3064];
        layer0[62][39:32] = buffer_data_4[3079:3072];
        layer1[62][7:0] = buffer_data_3[3047:3040];
        layer1[62][15:8] = buffer_data_3[3055:3048];
        layer1[62][23:16] = buffer_data_3[3063:3056];
        layer1[62][31:24] = buffer_data_3[3071:3064];
        layer1[62][39:32] = buffer_data_3[3079:3072];
        layer2[62][7:0] = buffer_data_2[3047:3040];
        layer2[62][15:8] = buffer_data_2[3055:3048];
        layer2[62][23:16] = buffer_data_2[3063:3056];
        layer2[62][31:24] = buffer_data_2[3071:3064];
        layer2[62][39:32] = buffer_data_2[3079:3072];
        layer3[62][7:0] = buffer_data_1[3047:3040];
        layer3[62][15:8] = buffer_data_1[3055:3048];
        layer3[62][23:16] = buffer_data_1[3063:3056];
        layer3[62][31:24] = buffer_data_1[3071:3064];
        layer3[62][39:32] = buffer_data_1[3079:3072];
        layer4[62][7:0] = buffer_data_0[3047:3040];
        layer4[62][15:8] = buffer_data_0[3055:3048];
        layer4[62][23:16] = buffer_data_0[3063:3056];
        layer4[62][31:24] = buffer_data_0[3071:3064];
        layer4[62][39:32] = buffer_data_0[3079:3072];
        layer0[63][7:0] = buffer_data_4[3055:3048];
        layer0[63][15:8] = buffer_data_4[3063:3056];
        layer0[63][23:16] = buffer_data_4[3071:3064];
        layer0[63][31:24] = buffer_data_4[3079:3072];
        layer0[63][39:32] = buffer_data_4[3087:3080];
        layer1[63][7:0] = buffer_data_3[3055:3048];
        layer1[63][15:8] = buffer_data_3[3063:3056];
        layer1[63][23:16] = buffer_data_3[3071:3064];
        layer1[63][31:24] = buffer_data_3[3079:3072];
        layer1[63][39:32] = buffer_data_3[3087:3080];
        layer2[63][7:0] = buffer_data_2[3055:3048];
        layer2[63][15:8] = buffer_data_2[3063:3056];
        layer2[63][23:16] = buffer_data_2[3071:3064];
        layer2[63][31:24] = buffer_data_2[3079:3072];
        layer2[63][39:32] = buffer_data_2[3087:3080];
        layer3[63][7:0] = buffer_data_1[3055:3048];
        layer3[63][15:8] = buffer_data_1[3063:3056];
        layer3[63][23:16] = buffer_data_1[3071:3064];
        layer3[63][31:24] = buffer_data_1[3079:3072];
        layer3[63][39:32] = buffer_data_1[3087:3080];
        layer4[63][7:0] = buffer_data_0[3055:3048];
        layer4[63][15:8] = buffer_data_0[3063:3056];
        layer4[63][23:16] = buffer_data_0[3071:3064];
        layer4[63][31:24] = buffer_data_0[3079:3072];
        layer4[63][39:32] = buffer_data_0[3087:3080];
    end
    ST_GAUSSIAN_6: begin
        layer0[0][7:0] = buffer_data_4[3063:3056];
        layer0[0][15:8] = buffer_data_4[3071:3064];
        layer0[0][23:16] = buffer_data_4[3079:3072];
        layer0[0][31:24] = buffer_data_4[3087:3080];
        layer0[0][39:32] = buffer_data_4[3095:3088];
        layer1[0][7:0] = buffer_data_3[3063:3056];
        layer1[0][15:8] = buffer_data_3[3071:3064];
        layer1[0][23:16] = buffer_data_3[3079:3072];
        layer1[0][31:24] = buffer_data_3[3087:3080];
        layer1[0][39:32] = buffer_data_3[3095:3088];
        layer2[0][7:0] = buffer_data_2[3063:3056];
        layer2[0][15:8] = buffer_data_2[3071:3064];
        layer2[0][23:16] = buffer_data_2[3079:3072];
        layer2[0][31:24] = buffer_data_2[3087:3080];
        layer2[0][39:32] = buffer_data_2[3095:3088];
        layer3[0][7:0] = buffer_data_1[3063:3056];
        layer3[0][15:8] = buffer_data_1[3071:3064];
        layer3[0][23:16] = buffer_data_1[3079:3072];
        layer3[0][31:24] = buffer_data_1[3087:3080];
        layer3[0][39:32] = buffer_data_1[3095:3088];
        layer4[0][7:0] = buffer_data_0[3063:3056];
        layer4[0][15:8] = buffer_data_0[3071:3064];
        layer4[0][23:16] = buffer_data_0[3079:3072];
        layer4[0][31:24] = buffer_data_0[3087:3080];
        layer4[0][39:32] = buffer_data_0[3095:3088];
        layer0[1][7:0] = buffer_data_4[3071:3064];
        layer0[1][15:8] = buffer_data_4[3079:3072];
        layer0[1][23:16] = buffer_data_4[3087:3080];
        layer0[1][31:24] = buffer_data_4[3095:3088];
        layer0[1][39:32] = buffer_data_4[3103:3096];
        layer1[1][7:0] = buffer_data_3[3071:3064];
        layer1[1][15:8] = buffer_data_3[3079:3072];
        layer1[1][23:16] = buffer_data_3[3087:3080];
        layer1[1][31:24] = buffer_data_3[3095:3088];
        layer1[1][39:32] = buffer_data_3[3103:3096];
        layer2[1][7:0] = buffer_data_2[3071:3064];
        layer2[1][15:8] = buffer_data_2[3079:3072];
        layer2[1][23:16] = buffer_data_2[3087:3080];
        layer2[1][31:24] = buffer_data_2[3095:3088];
        layer2[1][39:32] = buffer_data_2[3103:3096];
        layer3[1][7:0] = buffer_data_1[3071:3064];
        layer3[1][15:8] = buffer_data_1[3079:3072];
        layer3[1][23:16] = buffer_data_1[3087:3080];
        layer3[1][31:24] = buffer_data_1[3095:3088];
        layer3[1][39:32] = buffer_data_1[3103:3096];
        layer4[1][7:0] = buffer_data_0[3071:3064];
        layer4[1][15:8] = buffer_data_0[3079:3072];
        layer4[1][23:16] = buffer_data_0[3087:3080];
        layer4[1][31:24] = buffer_data_0[3095:3088];
        layer4[1][39:32] = buffer_data_0[3103:3096];
        layer0[2][7:0] = buffer_data_4[3079:3072];
        layer0[2][15:8] = buffer_data_4[3087:3080];
        layer0[2][23:16] = buffer_data_4[3095:3088];
        layer0[2][31:24] = buffer_data_4[3103:3096];
        layer0[2][39:32] = buffer_data_4[3111:3104];
        layer1[2][7:0] = buffer_data_3[3079:3072];
        layer1[2][15:8] = buffer_data_3[3087:3080];
        layer1[2][23:16] = buffer_data_3[3095:3088];
        layer1[2][31:24] = buffer_data_3[3103:3096];
        layer1[2][39:32] = buffer_data_3[3111:3104];
        layer2[2][7:0] = buffer_data_2[3079:3072];
        layer2[2][15:8] = buffer_data_2[3087:3080];
        layer2[2][23:16] = buffer_data_2[3095:3088];
        layer2[2][31:24] = buffer_data_2[3103:3096];
        layer2[2][39:32] = buffer_data_2[3111:3104];
        layer3[2][7:0] = buffer_data_1[3079:3072];
        layer3[2][15:8] = buffer_data_1[3087:3080];
        layer3[2][23:16] = buffer_data_1[3095:3088];
        layer3[2][31:24] = buffer_data_1[3103:3096];
        layer3[2][39:32] = buffer_data_1[3111:3104];
        layer4[2][7:0] = buffer_data_0[3079:3072];
        layer4[2][15:8] = buffer_data_0[3087:3080];
        layer4[2][23:16] = buffer_data_0[3095:3088];
        layer4[2][31:24] = buffer_data_0[3103:3096];
        layer4[2][39:32] = buffer_data_0[3111:3104];
        layer0[3][7:0] = buffer_data_4[3087:3080];
        layer0[3][15:8] = buffer_data_4[3095:3088];
        layer0[3][23:16] = buffer_data_4[3103:3096];
        layer0[3][31:24] = buffer_data_4[3111:3104];
        layer0[3][39:32] = buffer_data_4[3119:3112];
        layer1[3][7:0] = buffer_data_3[3087:3080];
        layer1[3][15:8] = buffer_data_3[3095:3088];
        layer1[3][23:16] = buffer_data_3[3103:3096];
        layer1[3][31:24] = buffer_data_3[3111:3104];
        layer1[3][39:32] = buffer_data_3[3119:3112];
        layer2[3][7:0] = buffer_data_2[3087:3080];
        layer2[3][15:8] = buffer_data_2[3095:3088];
        layer2[3][23:16] = buffer_data_2[3103:3096];
        layer2[3][31:24] = buffer_data_2[3111:3104];
        layer2[3][39:32] = buffer_data_2[3119:3112];
        layer3[3][7:0] = buffer_data_1[3087:3080];
        layer3[3][15:8] = buffer_data_1[3095:3088];
        layer3[3][23:16] = buffer_data_1[3103:3096];
        layer3[3][31:24] = buffer_data_1[3111:3104];
        layer3[3][39:32] = buffer_data_1[3119:3112];
        layer4[3][7:0] = buffer_data_0[3087:3080];
        layer4[3][15:8] = buffer_data_0[3095:3088];
        layer4[3][23:16] = buffer_data_0[3103:3096];
        layer4[3][31:24] = buffer_data_0[3111:3104];
        layer4[3][39:32] = buffer_data_0[3119:3112];
        layer0[4][7:0] = buffer_data_4[3095:3088];
        layer0[4][15:8] = buffer_data_4[3103:3096];
        layer0[4][23:16] = buffer_data_4[3111:3104];
        layer0[4][31:24] = buffer_data_4[3119:3112];
        layer0[4][39:32] = buffer_data_4[3127:3120];
        layer1[4][7:0] = buffer_data_3[3095:3088];
        layer1[4][15:8] = buffer_data_3[3103:3096];
        layer1[4][23:16] = buffer_data_3[3111:3104];
        layer1[4][31:24] = buffer_data_3[3119:3112];
        layer1[4][39:32] = buffer_data_3[3127:3120];
        layer2[4][7:0] = buffer_data_2[3095:3088];
        layer2[4][15:8] = buffer_data_2[3103:3096];
        layer2[4][23:16] = buffer_data_2[3111:3104];
        layer2[4][31:24] = buffer_data_2[3119:3112];
        layer2[4][39:32] = buffer_data_2[3127:3120];
        layer3[4][7:0] = buffer_data_1[3095:3088];
        layer3[4][15:8] = buffer_data_1[3103:3096];
        layer3[4][23:16] = buffer_data_1[3111:3104];
        layer3[4][31:24] = buffer_data_1[3119:3112];
        layer3[4][39:32] = buffer_data_1[3127:3120];
        layer4[4][7:0] = buffer_data_0[3095:3088];
        layer4[4][15:8] = buffer_data_0[3103:3096];
        layer4[4][23:16] = buffer_data_0[3111:3104];
        layer4[4][31:24] = buffer_data_0[3119:3112];
        layer4[4][39:32] = buffer_data_0[3127:3120];
        layer0[5][7:0] = buffer_data_4[3103:3096];
        layer0[5][15:8] = buffer_data_4[3111:3104];
        layer0[5][23:16] = buffer_data_4[3119:3112];
        layer0[5][31:24] = buffer_data_4[3127:3120];
        layer0[5][39:32] = buffer_data_4[3135:3128];
        layer1[5][7:0] = buffer_data_3[3103:3096];
        layer1[5][15:8] = buffer_data_3[3111:3104];
        layer1[5][23:16] = buffer_data_3[3119:3112];
        layer1[5][31:24] = buffer_data_3[3127:3120];
        layer1[5][39:32] = buffer_data_3[3135:3128];
        layer2[5][7:0] = buffer_data_2[3103:3096];
        layer2[5][15:8] = buffer_data_2[3111:3104];
        layer2[5][23:16] = buffer_data_2[3119:3112];
        layer2[5][31:24] = buffer_data_2[3127:3120];
        layer2[5][39:32] = buffer_data_2[3135:3128];
        layer3[5][7:0] = buffer_data_1[3103:3096];
        layer3[5][15:8] = buffer_data_1[3111:3104];
        layer3[5][23:16] = buffer_data_1[3119:3112];
        layer3[5][31:24] = buffer_data_1[3127:3120];
        layer3[5][39:32] = buffer_data_1[3135:3128];
        layer4[5][7:0] = buffer_data_0[3103:3096];
        layer4[5][15:8] = buffer_data_0[3111:3104];
        layer4[5][23:16] = buffer_data_0[3119:3112];
        layer4[5][31:24] = buffer_data_0[3127:3120];
        layer4[5][39:32] = buffer_data_0[3135:3128];
        layer0[6][7:0] = buffer_data_4[3111:3104];
        layer0[6][15:8] = buffer_data_4[3119:3112];
        layer0[6][23:16] = buffer_data_4[3127:3120];
        layer0[6][31:24] = buffer_data_4[3135:3128];
        layer0[6][39:32] = buffer_data_4[3143:3136];
        layer1[6][7:0] = buffer_data_3[3111:3104];
        layer1[6][15:8] = buffer_data_3[3119:3112];
        layer1[6][23:16] = buffer_data_3[3127:3120];
        layer1[6][31:24] = buffer_data_3[3135:3128];
        layer1[6][39:32] = buffer_data_3[3143:3136];
        layer2[6][7:0] = buffer_data_2[3111:3104];
        layer2[6][15:8] = buffer_data_2[3119:3112];
        layer2[6][23:16] = buffer_data_2[3127:3120];
        layer2[6][31:24] = buffer_data_2[3135:3128];
        layer2[6][39:32] = buffer_data_2[3143:3136];
        layer3[6][7:0] = buffer_data_1[3111:3104];
        layer3[6][15:8] = buffer_data_1[3119:3112];
        layer3[6][23:16] = buffer_data_1[3127:3120];
        layer3[6][31:24] = buffer_data_1[3135:3128];
        layer3[6][39:32] = buffer_data_1[3143:3136];
        layer4[6][7:0] = buffer_data_0[3111:3104];
        layer4[6][15:8] = buffer_data_0[3119:3112];
        layer4[6][23:16] = buffer_data_0[3127:3120];
        layer4[6][31:24] = buffer_data_0[3135:3128];
        layer4[6][39:32] = buffer_data_0[3143:3136];
        layer0[7][7:0] = buffer_data_4[3119:3112];
        layer0[7][15:8] = buffer_data_4[3127:3120];
        layer0[7][23:16] = buffer_data_4[3135:3128];
        layer0[7][31:24] = buffer_data_4[3143:3136];
        layer0[7][39:32] = buffer_data_4[3151:3144];
        layer1[7][7:0] = buffer_data_3[3119:3112];
        layer1[7][15:8] = buffer_data_3[3127:3120];
        layer1[7][23:16] = buffer_data_3[3135:3128];
        layer1[7][31:24] = buffer_data_3[3143:3136];
        layer1[7][39:32] = buffer_data_3[3151:3144];
        layer2[7][7:0] = buffer_data_2[3119:3112];
        layer2[7][15:8] = buffer_data_2[3127:3120];
        layer2[7][23:16] = buffer_data_2[3135:3128];
        layer2[7][31:24] = buffer_data_2[3143:3136];
        layer2[7][39:32] = buffer_data_2[3151:3144];
        layer3[7][7:0] = buffer_data_1[3119:3112];
        layer3[7][15:8] = buffer_data_1[3127:3120];
        layer3[7][23:16] = buffer_data_1[3135:3128];
        layer3[7][31:24] = buffer_data_1[3143:3136];
        layer3[7][39:32] = buffer_data_1[3151:3144];
        layer4[7][7:0] = buffer_data_0[3119:3112];
        layer4[7][15:8] = buffer_data_0[3127:3120];
        layer4[7][23:16] = buffer_data_0[3135:3128];
        layer4[7][31:24] = buffer_data_0[3143:3136];
        layer4[7][39:32] = buffer_data_0[3151:3144];
        layer0[8][7:0] = buffer_data_4[3127:3120];
        layer0[8][15:8] = buffer_data_4[3135:3128];
        layer0[8][23:16] = buffer_data_4[3143:3136];
        layer0[8][31:24] = buffer_data_4[3151:3144];
        layer0[8][39:32] = buffer_data_4[3159:3152];
        layer1[8][7:0] = buffer_data_3[3127:3120];
        layer1[8][15:8] = buffer_data_3[3135:3128];
        layer1[8][23:16] = buffer_data_3[3143:3136];
        layer1[8][31:24] = buffer_data_3[3151:3144];
        layer1[8][39:32] = buffer_data_3[3159:3152];
        layer2[8][7:0] = buffer_data_2[3127:3120];
        layer2[8][15:8] = buffer_data_2[3135:3128];
        layer2[8][23:16] = buffer_data_2[3143:3136];
        layer2[8][31:24] = buffer_data_2[3151:3144];
        layer2[8][39:32] = buffer_data_2[3159:3152];
        layer3[8][7:0] = buffer_data_1[3127:3120];
        layer3[8][15:8] = buffer_data_1[3135:3128];
        layer3[8][23:16] = buffer_data_1[3143:3136];
        layer3[8][31:24] = buffer_data_1[3151:3144];
        layer3[8][39:32] = buffer_data_1[3159:3152];
        layer4[8][7:0] = buffer_data_0[3127:3120];
        layer4[8][15:8] = buffer_data_0[3135:3128];
        layer4[8][23:16] = buffer_data_0[3143:3136];
        layer4[8][31:24] = buffer_data_0[3151:3144];
        layer4[8][39:32] = buffer_data_0[3159:3152];
        layer0[9][7:0] = buffer_data_4[3135:3128];
        layer0[9][15:8] = buffer_data_4[3143:3136];
        layer0[9][23:16] = buffer_data_4[3151:3144];
        layer0[9][31:24] = buffer_data_4[3159:3152];
        layer0[9][39:32] = buffer_data_4[3167:3160];
        layer1[9][7:0] = buffer_data_3[3135:3128];
        layer1[9][15:8] = buffer_data_3[3143:3136];
        layer1[9][23:16] = buffer_data_3[3151:3144];
        layer1[9][31:24] = buffer_data_3[3159:3152];
        layer1[9][39:32] = buffer_data_3[3167:3160];
        layer2[9][7:0] = buffer_data_2[3135:3128];
        layer2[9][15:8] = buffer_data_2[3143:3136];
        layer2[9][23:16] = buffer_data_2[3151:3144];
        layer2[9][31:24] = buffer_data_2[3159:3152];
        layer2[9][39:32] = buffer_data_2[3167:3160];
        layer3[9][7:0] = buffer_data_1[3135:3128];
        layer3[9][15:8] = buffer_data_1[3143:3136];
        layer3[9][23:16] = buffer_data_1[3151:3144];
        layer3[9][31:24] = buffer_data_1[3159:3152];
        layer3[9][39:32] = buffer_data_1[3167:3160];
        layer4[9][7:0] = buffer_data_0[3135:3128];
        layer4[9][15:8] = buffer_data_0[3143:3136];
        layer4[9][23:16] = buffer_data_0[3151:3144];
        layer4[9][31:24] = buffer_data_0[3159:3152];
        layer4[9][39:32] = buffer_data_0[3167:3160];
        layer0[10][7:0] = buffer_data_4[3143:3136];
        layer0[10][15:8] = buffer_data_4[3151:3144];
        layer0[10][23:16] = buffer_data_4[3159:3152];
        layer0[10][31:24] = buffer_data_4[3167:3160];
        layer0[10][39:32] = buffer_data_4[3175:3168];
        layer1[10][7:0] = buffer_data_3[3143:3136];
        layer1[10][15:8] = buffer_data_3[3151:3144];
        layer1[10][23:16] = buffer_data_3[3159:3152];
        layer1[10][31:24] = buffer_data_3[3167:3160];
        layer1[10][39:32] = buffer_data_3[3175:3168];
        layer2[10][7:0] = buffer_data_2[3143:3136];
        layer2[10][15:8] = buffer_data_2[3151:3144];
        layer2[10][23:16] = buffer_data_2[3159:3152];
        layer2[10][31:24] = buffer_data_2[3167:3160];
        layer2[10][39:32] = buffer_data_2[3175:3168];
        layer3[10][7:0] = buffer_data_1[3143:3136];
        layer3[10][15:8] = buffer_data_1[3151:3144];
        layer3[10][23:16] = buffer_data_1[3159:3152];
        layer3[10][31:24] = buffer_data_1[3167:3160];
        layer3[10][39:32] = buffer_data_1[3175:3168];
        layer4[10][7:0] = buffer_data_0[3143:3136];
        layer4[10][15:8] = buffer_data_0[3151:3144];
        layer4[10][23:16] = buffer_data_0[3159:3152];
        layer4[10][31:24] = buffer_data_0[3167:3160];
        layer4[10][39:32] = buffer_data_0[3175:3168];
        layer0[11][7:0] = buffer_data_4[3151:3144];
        layer0[11][15:8] = buffer_data_4[3159:3152];
        layer0[11][23:16] = buffer_data_4[3167:3160];
        layer0[11][31:24] = buffer_data_4[3175:3168];
        layer0[11][39:32] = buffer_data_4[3183:3176];
        layer1[11][7:0] = buffer_data_3[3151:3144];
        layer1[11][15:8] = buffer_data_3[3159:3152];
        layer1[11][23:16] = buffer_data_3[3167:3160];
        layer1[11][31:24] = buffer_data_3[3175:3168];
        layer1[11][39:32] = buffer_data_3[3183:3176];
        layer2[11][7:0] = buffer_data_2[3151:3144];
        layer2[11][15:8] = buffer_data_2[3159:3152];
        layer2[11][23:16] = buffer_data_2[3167:3160];
        layer2[11][31:24] = buffer_data_2[3175:3168];
        layer2[11][39:32] = buffer_data_2[3183:3176];
        layer3[11][7:0] = buffer_data_1[3151:3144];
        layer3[11][15:8] = buffer_data_1[3159:3152];
        layer3[11][23:16] = buffer_data_1[3167:3160];
        layer3[11][31:24] = buffer_data_1[3175:3168];
        layer3[11][39:32] = buffer_data_1[3183:3176];
        layer4[11][7:0] = buffer_data_0[3151:3144];
        layer4[11][15:8] = buffer_data_0[3159:3152];
        layer4[11][23:16] = buffer_data_0[3167:3160];
        layer4[11][31:24] = buffer_data_0[3175:3168];
        layer4[11][39:32] = buffer_data_0[3183:3176];
        layer0[12][7:0] = buffer_data_4[3159:3152];
        layer0[12][15:8] = buffer_data_4[3167:3160];
        layer0[12][23:16] = buffer_data_4[3175:3168];
        layer0[12][31:24] = buffer_data_4[3183:3176];
        layer0[12][39:32] = buffer_data_4[3191:3184];
        layer1[12][7:0] = buffer_data_3[3159:3152];
        layer1[12][15:8] = buffer_data_3[3167:3160];
        layer1[12][23:16] = buffer_data_3[3175:3168];
        layer1[12][31:24] = buffer_data_3[3183:3176];
        layer1[12][39:32] = buffer_data_3[3191:3184];
        layer2[12][7:0] = buffer_data_2[3159:3152];
        layer2[12][15:8] = buffer_data_2[3167:3160];
        layer2[12][23:16] = buffer_data_2[3175:3168];
        layer2[12][31:24] = buffer_data_2[3183:3176];
        layer2[12][39:32] = buffer_data_2[3191:3184];
        layer3[12][7:0] = buffer_data_1[3159:3152];
        layer3[12][15:8] = buffer_data_1[3167:3160];
        layer3[12][23:16] = buffer_data_1[3175:3168];
        layer3[12][31:24] = buffer_data_1[3183:3176];
        layer3[12][39:32] = buffer_data_1[3191:3184];
        layer4[12][7:0] = buffer_data_0[3159:3152];
        layer4[12][15:8] = buffer_data_0[3167:3160];
        layer4[12][23:16] = buffer_data_0[3175:3168];
        layer4[12][31:24] = buffer_data_0[3183:3176];
        layer4[12][39:32] = buffer_data_0[3191:3184];
        layer0[13][7:0] = buffer_data_4[3167:3160];
        layer0[13][15:8] = buffer_data_4[3175:3168];
        layer0[13][23:16] = buffer_data_4[3183:3176];
        layer0[13][31:24] = buffer_data_4[3191:3184];
        layer0[13][39:32] = buffer_data_4[3199:3192];
        layer1[13][7:0] = buffer_data_3[3167:3160];
        layer1[13][15:8] = buffer_data_3[3175:3168];
        layer1[13][23:16] = buffer_data_3[3183:3176];
        layer1[13][31:24] = buffer_data_3[3191:3184];
        layer1[13][39:32] = buffer_data_3[3199:3192];
        layer2[13][7:0] = buffer_data_2[3167:3160];
        layer2[13][15:8] = buffer_data_2[3175:3168];
        layer2[13][23:16] = buffer_data_2[3183:3176];
        layer2[13][31:24] = buffer_data_2[3191:3184];
        layer2[13][39:32] = buffer_data_2[3199:3192];
        layer3[13][7:0] = buffer_data_1[3167:3160];
        layer3[13][15:8] = buffer_data_1[3175:3168];
        layer3[13][23:16] = buffer_data_1[3183:3176];
        layer3[13][31:24] = buffer_data_1[3191:3184];
        layer3[13][39:32] = buffer_data_1[3199:3192];
        layer4[13][7:0] = buffer_data_0[3167:3160];
        layer4[13][15:8] = buffer_data_0[3175:3168];
        layer4[13][23:16] = buffer_data_0[3183:3176];
        layer4[13][31:24] = buffer_data_0[3191:3184];
        layer4[13][39:32] = buffer_data_0[3199:3192];
        layer0[14][7:0] = buffer_data_4[3175:3168];
        layer0[14][15:8] = buffer_data_4[3183:3176];
        layer0[14][23:16] = buffer_data_4[3191:3184];
        layer0[14][31:24] = buffer_data_4[3199:3192];
        layer0[14][39:32] = buffer_data_4[3207:3200];
        layer1[14][7:0] = buffer_data_3[3175:3168];
        layer1[14][15:8] = buffer_data_3[3183:3176];
        layer1[14][23:16] = buffer_data_3[3191:3184];
        layer1[14][31:24] = buffer_data_3[3199:3192];
        layer1[14][39:32] = buffer_data_3[3207:3200];
        layer2[14][7:0] = buffer_data_2[3175:3168];
        layer2[14][15:8] = buffer_data_2[3183:3176];
        layer2[14][23:16] = buffer_data_2[3191:3184];
        layer2[14][31:24] = buffer_data_2[3199:3192];
        layer2[14][39:32] = buffer_data_2[3207:3200];
        layer3[14][7:0] = buffer_data_1[3175:3168];
        layer3[14][15:8] = buffer_data_1[3183:3176];
        layer3[14][23:16] = buffer_data_1[3191:3184];
        layer3[14][31:24] = buffer_data_1[3199:3192];
        layer3[14][39:32] = buffer_data_1[3207:3200];
        layer4[14][7:0] = buffer_data_0[3175:3168];
        layer4[14][15:8] = buffer_data_0[3183:3176];
        layer4[14][23:16] = buffer_data_0[3191:3184];
        layer4[14][31:24] = buffer_data_0[3199:3192];
        layer4[14][39:32] = buffer_data_0[3207:3200];
        layer0[15][7:0] = buffer_data_4[3183:3176];
        layer0[15][15:8] = buffer_data_4[3191:3184];
        layer0[15][23:16] = buffer_data_4[3199:3192];
        layer0[15][31:24] = buffer_data_4[3207:3200];
        layer0[15][39:32] = buffer_data_4[3215:3208];
        layer1[15][7:0] = buffer_data_3[3183:3176];
        layer1[15][15:8] = buffer_data_3[3191:3184];
        layer1[15][23:16] = buffer_data_3[3199:3192];
        layer1[15][31:24] = buffer_data_3[3207:3200];
        layer1[15][39:32] = buffer_data_3[3215:3208];
        layer2[15][7:0] = buffer_data_2[3183:3176];
        layer2[15][15:8] = buffer_data_2[3191:3184];
        layer2[15][23:16] = buffer_data_2[3199:3192];
        layer2[15][31:24] = buffer_data_2[3207:3200];
        layer2[15][39:32] = buffer_data_2[3215:3208];
        layer3[15][7:0] = buffer_data_1[3183:3176];
        layer3[15][15:8] = buffer_data_1[3191:3184];
        layer3[15][23:16] = buffer_data_1[3199:3192];
        layer3[15][31:24] = buffer_data_1[3207:3200];
        layer3[15][39:32] = buffer_data_1[3215:3208];
        layer4[15][7:0] = buffer_data_0[3183:3176];
        layer4[15][15:8] = buffer_data_0[3191:3184];
        layer4[15][23:16] = buffer_data_0[3199:3192];
        layer4[15][31:24] = buffer_data_0[3207:3200];
        layer4[15][39:32] = buffer_data_0[3215:3208];
        layer0[16][7:0] = buffer_data_4[3191:3184];
        layer0[16][15:8] = buffer_data_4[3199:3192];
        layer0[16][23:16] = buffer_data_4[3207:3200];
        layer0[16][31:24] = buffer_data_4[3215:3208];
        layer0[16][39:32] = buffer_data_4[3223:3216];
        layer1[16][7:0] = buffer_data_3[3191:3184];
        layer1[16][15:8] = buffer_data_3[3199:3192];
        layer1[16][23:16] = buffer_data_3[3207:3200];
        layer1[16][31:24] = buffer_data_3[3215:3208];
        layer1[16][39:32] = buffer_data_3[3223:3216];
        layer2[16][7:0] = buffer_data_2[3191:3184];
        layer2[16][15:8] = buffer_data_2[3199:3192];
        layer2[16][23:16] = buffer_data_2[3207:3200];
        layer2[16][31:24] = buffer_data_2[3215:3208];
        layer2[16][39:32] = buffer_data_2[3223:3216];
        layer3[16][7:0] = buffer_data_1[3191:3184];
        layer3[16][15:8] = buffer_data_1[3199:3192];
        layer3[16][23:16] = buffer_data_1[3207:3200];
        layer3[16][31:24] = buffer_data_1[3215:3208];
        layer3[16][39:32] = buffer_data_1[3223:3216];
        layer4[16][7:0] = buffer_data_0[3191:3184];
        layer4[16][15:8] = buffer_data_0[3199:3192];
        layer4[16][23:16] = buffer_data_0[3207:3200];
        layer4[16][31:24] = buffer_data_0[3215:3208];
        layer4[16][39:32] = buffer_data_0[3223:3216];
        layer0[17][7:0] = buffer_data_4[3199:3192];
        layer0[17][15:8] = buffer_data_4[3207:3200];
        layer0[17][23:16] = buffer_data_4[3215:3208];
        layer0[17][31:24] = buffer_data_4[3223:3216];
        layer0[17][39:32] = buffer_data_4[3231:3224];
        layer1[17][7:0] = buffer_data_3[3199:3192];
        layer1[17][15:8] = buffer_data_3[3207:3200];
        layer1[17][23:16] = buffer_data_3[3215:3208];
        layer1[17][31:24] = buffer_data_3[3223:3216];
        layer1[17][39:32] = buffer_data_3[3231:3224];
        layer2[17][7:0] = buffer_data_2[3199:3192];
        layer2[17][15:8] = buffer_data_2[3207:3200];
        layer2[17][23:16] = buffer_data_2[3215:3208];
        layer2[17][31:24] = buffer_data_2[3223:3216];
        layer2[17][39:32] = buffer_data_2[3231:3224];
        layer3[17][7:0] = buffer_data_1[3199:3192];
        layer3[17][15:8] = buffer_data_1[3207:3200];
        layer3[17][23:16] = buffer_data_1[3215:3208];
        layer3[17][31:24] = buffer_data_1[3223:3216];
        layer3[17][39:32] = buffer_data_1[3231:3224];
        layer4[17][7:0] = buffer_data_0[3199:3192];
        layer4[17][15:8] = buffer_data_0[3207:3200];
        layer4[17][23:16] = buffer_data_0[3215:3208];
        layer4[17][31:24] = buffer_data_0[3223:3216];
        layer4[17][39:32] = buffer_data_0[3231:3224];
        layer0[18][7:0] = buffer_data_4[3207:3200];
        layer0[18][15:8] = buffer_data_4[3215:3208];
        layer0[18][23:16] = buffer_data_4[3223:3216];
        layer0[18][31:24] = buffer_data_4[3231:3224];
        layer0[18][39:32] = buffer_data_4[3239:3232];
        layer1[18][7:0] = buffer_data_3[3207:3200];
        layer1[18][15:8] = buffer_data_3[3215:3208];
        layer1[18][23:16] = buffer_data_3[3223:3216];
        layer1[18][31:24] = buffer_data_3[3231:3224];
        layer1[18][39:32] = buffer_data_3[3239:3232];
        layer2[18][7:0] = buffer_data_2[3207:3200];
        layer2[18][15:8] = buffer_data_2[3215:3208];
        layer2[18][23:16] = buffer_data_2[3223:3216];
        layer2[18][31:24] = buffer_data_2[3231:3224];
        layer2[18][39:32] = buffer_data_2[3239:3232];
        layer3[18][7:0] = buffer_data_1[3207:3200];
        layer3[18][15:8] = buffer_data_1[3215:3208];
        layer3[18][23:16] = buffer_data_1[3223:3216];
        layer3[18][31:24] = buffer_data_1[3231:3224];
        layer3[18][39:32] = buffer_data_1[3239:3232];
        layer4[18][7:0] = buffer_data_0[3207:3200];
        layer4[18][15:8] = buffer_data_0[3215:3208];
        layer4[18][23:16] = buffer_data_0[3223:3216];
        layer4[18][31:24] = buffer_data_0[3231:3224];
        layer4[18][39:32] = buffer_data_0[3239:3232];
        layer0[19][7:0] = buffer_data_4[3215:3208];
        layer0[19][15:8] = buffer_data_4[3223:3216];
        layer0[19][23:16] = buffer_data_4[3231:3224];
        layer0[19][31:24] = buffer_data_4[3239:3232];
        layer0[19][39:32] = buffer_data_4[3247:3240];
        layer1[19][7:0] = buffer_data_3[3215:3208];
        layer1[19][15:8] = buffer_data_3[3223:3216];
        layer1[19][23:16] = buffer_data_3[3231:3224];
        layer1[19][31:24] = buffer_data_3[3239:3232];
        layer1[19][39:32] = buffer_data_3[3247:3240];
        layer2[19][7:0] = buffer_data_2[3215:3208];
        layer2[19][15:8] = buffer_data_2[3223:3216];
        layer2[19][23:16] = buffer_data_2[3231:3224];
        layer2[19][31:24] = buffer_data_2[3239:3232];
        layer2[19][39:32] = buffer_data_2[3247:3240];
        layer3[19][7:0] = buffer_data_1[3215:3208];
        layer3[19][15:8] = buffer_data_1[3223:3216];
        layer3[19][23:16] = buffer_data_1[3231:3224];
        layer3[19][31:24] = buffer_data_1[3239:3232];
        layer3[19][39:32] = buffer_data_1[3247:3240];
        layer4[19][7:0] = buffer_data_0[3215:3208];
        layer4[19][15:8] = buffer_data_0[3223:3216];
        layer4[19][23:16] = buffer_data_0[3231:3224];
        layer4[19][31:24] = buffer_data_0[3239:3232];
        layer4[19][39:32] = buffer_data_0[3247:3240];
        layer0[20][7:0] = buffer_data_4[3223:3216];
        layer0[20][15:8] = buffer_data_4[3231:3224];
        layer0[20][23:16] = buffer_data_4[3239:3232];
        layer0[20][31:24] = buffer_data_4[3247:3240];
        layer0[20][39:32] = buffer_data_4[3255:3248];
        layer1[20][7:0] = buffer_data_3[3223:3216];
        layer1[20][15:8] = buffer_data_3[3231:3224];
        layer1[20][23:16] = buffer_data_3[3239:3232];
        layer1[20][31:24] = buffer_data_3[3247:3240];
        layer1[20][39:32] = buffer_data_3[3255:3248];
        layer2[20][7:0] = buffer_data_2[3223:3216];
        layer2[20][15:8] = buffer_data_2[3231:3224];
        layer2[20][23:16] = buffer_data_2[3239:3232];
        layer2[20][31:24] = buffer_data_2[3247:3240];
        layer2[20][39:32] = buffer_data_2[3255:3248];
        layer3[20][7:0] = buffer_data_1[3223:3216];
        layer3[20][15:8] = buffer_data_1[3231:3224];
        layer3[20][23:16] = buffer_data_1[3239:3232];
        layer3[20][31:24] = buffer_data_1[3247:3240];
        layer3[20][39:32] = buffer_data_1[3255:3248];
        layer4[20][7:0] = buffer_data_0[3223:3216];
        layer4[20][15:8] = buffer_data_0[3231:3224];
        layer4[20][23:16] = buffer_data_0[3239:3232];
        layer4[20][31:24] = buffer_data_0[3247:3240];
        layer4[20][39:32] = buffer_data_0[3255:3248];
        layer0[21][7:0] = buffer_data_4[3231:3224];
        layer0[21][15:8] = buffer_data_4[3239:3232];
        layer0[21][23:16] = buffer_data_4[3247:3240];
        layer0[21][31:24] = buffer_data_4[3255:3248];
        layer0[21][39:32] = buffer_data_4[3263:3256];
        layer1[21][7:0] = buffer_data_3[3231:3224];
        layer1[21][15:8] = buffer_data_3[3239:3232];
        layer1[21][23:16] = buffer_data_3[3247:3240];
        layer1[21][31:24] = buffer_data_3[3255:3248];
        layer1[21][39:32] = buffer_data_3[3263:3256];
        layer2[21][7:0] = buffer_data_2[3231:3224];
        layer2[21][15:8] = buffer_data_2[3239:3232];
        layer2[21][23:16] = buffer_data_2[3247:3240];
        layer2[21][31:24] = buffer_data_2[3255:3248];
        layer2[21][39:32] = buffer_data_2[3263:3256];
        layer3[21][7:0] = buffer_data_1[3231:3224];
        layer3[21][15:8] = buffer_data_1[3239:3232];
        layer3[21][23:16] = buffer_data_1[3247:3240];
        layer3[21][31:24] = buffer_data_1[3255:3248];
        layer3[21][39:32] = buffer_data_1[3263:3256];
        layer4[21][7:0] = buffer_data_0[3231:3224];
        layer4[21][15:8] = buffer_data_0[3239:3232];
        layer4[21][23:16] = buffer_data_0[3247:3240];
        layer4[21][31:24] = buffer_data_0[3255:3248];
        layer4[21][39:32] = buffer_data_0[3263:3256];
        layer0[22][7:0] = buffer_data_4[3239:3232];
        layer0[22][15:8] = buffer_data_4[3247:3240];
        layer0[22][23:16] = buffer_data_4[3255:3248];
        layer0[22][31:24] = buffer_data_4[3263:3256];
        layer0[22][39:32] = buffer_data_4[3271:3264];
        layer1[22][7:0] = buffer_data_3[3239:3232];
        layer1[22][15:8] = buffer_data_3[3247:3240];
        layer1[22][23:16] = buffer_data_3[3255:3248];
        layer1[22][31:24] = buffer_data_3[3263:3256];
        layer1[22][39:32] = buffer_data_3[3271:3264];
        layer2[22][7:0] = buffer_data_2[3239:3232];
        layer2[22][15:8] = buffer_data_2[3247:3240];
        layer2[22][23:16] = buffer_data_2[3255:3248];
        layer2[22][31:24] = buffer_data_2[3263:3256];
        layer2[22][39:32] = buffer_data_2[3271:3264];
        layer3[22][7:0] = buffer_data_1[3239:3232];
        layer3[22][15:8] = buffer_data_1[3247:3240];
        layer3[22][23:16] = buffer_data_1[3255:3248];
        layer3[22][31:24] = buffer_data_1[3263:3256];
        layer3[22][39:32] = buffer_data_1[3271:3264];
        layer4[22][7:0] = buffer_data_0[3239:3232];
        layer4[22][15:8] = buffer_data_0[3247:3240];
        layer4[22][23:16] = buffer_data_0[3255:3248];
        layer4[22][31:24] = buffer_data_0[3263:3256];
        layer4[22][39:32] = buffer_data_0[3271:3264];
        layer0[23][7:0] = buffer_data_4[3247:3240];
        layer0[23][15:8] = buffer_data_4[3255:3248];
        layer0[23][23:16] = buffer_data_4[3263:3256];
        layer0[23][31:24] = buffer_data_4[3271:3264];
        layer0[23][39:32] = buffer_data_4[3279:3272];
        layer1[23][7:0] = buffer_data_3[3247:3240];
        layer1[23][15:8] = buffer_data_3[3255:3248];
        layer1[23][23:16] = buffer_data_3[3263:3256];
        layer1[23][31:24] = buffer_data_3[3271:3264];
        layer1[23][39:32] = buffer_data_3[3279:3272];
        layer2[23][7:0] = buffer_data_2[3247:3240];
        layer2[23][15:8] = buffer_data_2[3255:3248];
        layer2[23][23:16] = buffer_data_2[3263:3256];
        layer2[23][31:24] = buffer_data_2[3271:3264];
        layer2[23][39:32] = buffer_data_2[3279:3272];
        layer3[23][7:0] = buffer_data_1[3247:3240];
        layer3[23][15:8] = buffer_data_1[3255:3248];
        layer3[23][23:16] = buffer_data_1[3263:3256];
        layer3[23][31:24] = buffer_data_1[3271:3264];
        layer3[23][39:32] = buffer_data_1[3279:3272];
        layer4[23][7:0] = buffer_data_0[3247:3240];
        layer4[23][15:8] = buffer_data_0[3255:3248];
        layer4[23][23:16] = buffer_data_0[3263:3256];
        layer4[23][31:24] = buffer_data_0[3271:3264];
        layer4[23][39:32] = buffer_data_0[3279:3272];
        layer0[24][7:0] = buffer_data_4[3255:3248];
        layer0[24][15:8] = buffer_data_4[3263:3256];
        layer0[24][23:16] = buffer_data_4[3271:3264];
        layer0[24][31:24] = buffer_data_4[3279:3272];
        layer0[24][39:32] = buffer_data_4[3287:3280];
        layer1[24][7:0] = buffer_data_3[3255:3248];
        layer1[24][15:8] = buffer_data_3[3263:3256];
        layer1[24][23:16] = buffer_data_3[3271:3264];
        layer1[24][31:24] = buffer_data_3[3279:3272];
        layer1[24][39:32] = buffer_data_3[3287:3280];
        layer2[24][7:0] = buffer_data_2[3255:3248];
        layer2[24][15:8] = buffer_data_2[3263:3256];
        layer2[24][23:16] = buffer_data_2[3271:3264];
        layer2[24][31:24] = buffer_data_2[3279:3272];
        layer2[24][39:32] = buffer_data_2[3287:3280];
        layer3[24][7:0] = buffer_data_1[3255:3248];
        layer3[24][15:8] = buffer_data_1[3263:3256];
        layer3[24][23:16] = buffer_data_1[3271:3264];
        layer3[24][31:24] = buffer_data_1[3279:3272];
        layer3[24][39:32] = buffer_data_1[3287:3280];
        layer4[24][7:0] = buffer_data_0[3255:3248];
        layer4[24][15:8] = buffer_data_0[3263:3256];
        layer4[24][23:16] = buffer_data_0[3271:3264];
        layer4[24][31:24] = buffer_data_0[3279:3272];
        layer4[24][39:32] = buffer_data_0[3287:3280];
        layer0[25][7:0] = buffer_data_4[3263:3256];
        layer0[25][15:8] = buffer_data_4[3271:3264];
        layer0[25][23:16] = buffer_data_4[3279:3272];
        layer0[25][31:24] = buffer_data_4[3287:3280];
        layer0[25][39:32] = buffer_data_4[3295:3288];
        layer1[25][7:0] = buffer_data_3[3263:3256];
        layer1[25][15:8] = buffer_data_3[3271:3264];
        layer1[25][23:16] = buffer_data_3[3279:3272];
        layer1[25][31:24] = buffer_data_3[3287:3280];
        layer1[25][39:32] = buffer_data_3[3295:3288];
        layer2[25][7:0] = buffer_data_2[3263:3256];
        layer2[25][15:8] = buffer_data_2[3271:3264];
        layer2[25][23:16] = buffer_data_2[3279:3272];
        layer2[25][31:24] = buffer_data_2[3287:3280];
        layer2[25][39:32] = buffer_data_2[3295:3288];
        layer3[25][7:0] = buffer_data_1[3263:3256];
        layer3[25][15:8] = buffer_data_1[3271:3264];
        layer3[25][23:16] = buffer_data_1[3279:3272];
        layer3[25][31:24] = buffer_data_1[3287:3280];
        layer3[25][39:32] = buffer_data_1[3295:3288];
        layer4[25][7:0] = buffer_data_0[3263:3256];
        layer4[25][15:8] = buffer_data_0[3271:3264];
        layer4[25][23:16] = buffer_data_0[3279:3272];
        layer4[25][31:24] = buffer_data_0[3287:3280];
        layer4[25][39:32] = buffer_data_0[3295:3288];
        layer0[26][7:0] = buffer_data_4[3271:3264];
        layer0[26][15:8] = buffer_data_4[3279:3272];
        layer0[26][23:16] = buffer_data_4[3287:3280];
        layer0[26][31:24] = buffer_data_4[3295:3288];
        layer0[26][39:32] = buffer_data_4[3303:3296];
        layer1[26][7:0] = buffer_data_3[3271:3264];
        layer1[26][15:8] = buffer_data_3[3279:3272];
        layer1[26][23:16] = buffer_data_3[3287:3280];
        layer1[26][31:24] = buffer_data_3[3295:3288];
        layer1[26][39:32] = buffer_data_3[3303:3296];
        layer2[26][7:0] = buffer_data_2[3271:3264];
        layer2[26][15:8] = buffer_data_2[3279:3272];
        layer2[26][23:16] = buffer_data_2[3287:3280];
        layer2[26][31:24] = buffer_data_2[3295:3288];
        layer2[26][39:32] = buffer_data_2[3303:3296];
        layer3[26][7:0] = buffer_data_1[3271:3264];
        layer3[26][15:8] = buffer_data_1[3279:3272];
        layer3[26][23:16] = buffer_data_1[3287:3280];
        layer3[26][31:24] = buffer_data_1[3295:3288];
        layer3[26][39:32] = buffer_data_1[3303:3296];
        layer4[26][7:0] = buffer_data_0[3271:3264];
        layer4[26][15:8] = buffer_data_0[3279:3272];
        layer4[26][23:16] = buffer_data_0[3287:3280];
        layer4[26][31:24] = buffer_data_0[3295:3288];
        layer4[26][39:32] = buffer_data_0[3303:3296];
        layer0[27][7:0] = buffer_data_4[3279:3272];
        layer0[27][15:8] = buffer_data_4[3287:3280];
        layer0[27][23:16] = buffer_data_4[3295:3288];
        layer0[27][31:24] = buffer_data_4[3303:3296];
        layer0[27][39:32] = buffer_data_4[3311:3304];
        layer1[27][7:0] = buffer_data_3[3279:3272];
        layer1[27][15:8] = buffer_data_3[3287:3280];
        layer1[27][23:16] = buffer_data_3[3295:3288];
        layer1[27][31:24] = buffer_data_3[3303:3296];
        layer1[27][39:32] = buffer_data_3[3311:3304];
        layer2[27][7:0] = buffer_data_2[3279:3272];
        layer2[27][15:8] = buffer_data_2[3287:3280];
        layer2[27][23:16] = buffer_data_2[3295:3288];
        layer2[27][31:24] = buffer_data_2[3303:3296];
        layer2[27][39:32] = buffer_data_2[3311:3304];
        layer3[27][7:0] = buffer_data_1[3279:3272];
        layer3[27][15:8] = buffer_data_1[3287:3280];
        layer3[27][23:16] = buffer_data_1[3295:3288];
        layer3[27][31:24] = buffer_data_1[3303:3296];
        layer3[27][39:32] = buffer_data_1[3311:3304];
        layer4[27][7:0] = buffer_data_0[3279:3272];
        layer4[27][15:8] = buffer_data_0[3287:3280];
        layer4[27][23:16] = buffer_data_0[3295:3288];
        layer4[27][31:24] = buffer_data_0[3303:3296];
        layer4[27][39:32] = buffer_data_0[3311:3304];
        layer0[28][7:0] = buffer_data_4[3287:3280];
        layer0[28][15:8] = buffer_data_4[3295:3288];
        layer0[28][23:16] = buffer_data_4[3303:3296];
        layer0[28][31:24] = buffer_data_4[3311:3304];
        layer0[28][39:32] = buffer_data_4[3319:3312];
        layer1[28][7:0] = buffer_data_3[3287:3280];
        layer1[28][15:8] = buffer_data_3[3295:3288];
        layer1[28][23:16] = buffer_data_3[3303:3296];
        layer1[28][31:24] = buffer_data_3[3311:3304];
        layer1[28][39:32] = buffer_data_3[3319:3312];
        layer2[28][7:0] = buffer_data_2[3287:3280];
        layer2[28][15:8] = buffer_data_2[3295:3288];
        layer2[28][23:16] = buffer_data_2[3303:3296];
        layer2[28][31:24] = buffer_data_2[3311:3304];
        layer2[28][39:32] = buffer_data_2[3319:3312];
        layer3[28][7:0] = buffer_data_1[3287:3280];
        layer3[28][15:8] = buffer_data_1[3295:3288];
        layer3[28][23:16] = buffer_data_1[3303:3296];
        layer3[28][31:24] = buffer_data_1[3311:3304];
        layer3[28][39:32] = buffer_data_1[3319:3312];
        layer4[28][7:0] = buffer_data_0[3287:3280];
        layer4[28][15:8] = buffer_data_0[3295:3288];
        layer4[28][23:16] = buffer_data_0[3303:3296];
        layer4[28][31:24] = buffer_data_0[3311:3304];
        layer4[28][39:32] = buffer_data_0[3319:3312];
        layer0[29][7:0] = buffer_data_4[3295:3288];
        layer0[29][15:8] = buffer_data_4[3303:3296];
        layer0[29][23:16] = buffer_data_4[3311:3304];
        layer0[29][31:24] = buffer_data_4[3319:3312];
        layer0[29][39:32] = buffer_data_4[3327:3320];
        layer1[29][7:0] = buffer_data_3[3295:3288];
        layer1[29][15:8] = buffer_data_3[3303:3296];
        layer1[29][23:16] = buffer_data_3[3311:3304];
        layer1[29][31:24] = buffer_data_3[3319:3312];
        layer1[29][39:32] = buffer_data_3[3327:3320];
        layer2[29][7:0] = buffer_data_2[3295:3288];
        layer2[29][15:8] = buffer_data_2[3303:3296];
        layer2[29][23:16] = buffer_data_2[3311:3304];
        layer2[29][31:24] = buffer_data_2[3319:3312];
        layer2[29][39:32] = buffer_data_2[3327:3320];
        layer3[29][7:0] = buffer_data_1[3295:3288];
        layer3[29][15:8] = buffer_data_1[3303:3296];
        layer3[29][23:16] = buffer_data_1[3311:3304];
        layer3[29][31:24] = buffer_data_1[3319:3312];
        layer3[29][39:32] = buffer_data_1[3327:3320];
        layer4[29][7:0] = buffer_data_0[3295:3288];
        layer4[29][15:8] = buffer_data_0[3303:3296];
        layer4[29][23:16] = buffer_data_0[3311:3304];
        layer4[29][31:24] = buffer_data_0[3319:3312];
        layer4[29][39:32] = buffer_data_0[3327:3320];
        layer0[30][7:0] = buffer_data_4[3303:3296];
        layer0[30][15:8] = buffer_data_4[3311:3304];
        layer0[30][23:16] = buffer_data_4[3319:3312];
        layer0[30][31:24] = buffer_data_4[3327:3320];
        layer0[30][39:32] = buffer_data_4[3335:3328];
        layer1[30][7:0] = buffer_data_3[3303:3296];
        layer1[30][15:8] = buffer_data_3[3311:3304];
        layer1[30][23:16] = buffer_data_3[3319:3312];
        layer1[30][31:24] = buffer_data_3[3327:3320];
        layer1[30][39:32] = buffer_data_3[3335:3328];
        layer2[30][7:0] = buffer_data_2[3303:3296];
        layer2[30][15:8] = buffer_data_2[3311:3304];
        layer2[30][23:16] = buffer_data_2[3319:3312];
        layer2[30][31:24] = buffer_data_2[3327:3320];
        layer2[30][39:32] = buffer_data_2[3335:3328];
        layer3[30][7:0] = buffer_data_1[3303:3296];
        layer3[30][15:8] = buffer_data_1[3311:3304];
        layer3[30][23:16] = buffer_data_1[3319:3312];
        layer3[30][31:24] = buffer_data_1[3327:3320];
        layer3[30][39:32] = buffer_data_1[3335:3328];
        layer4[30][7:0] = buffer_data_0[3303:3296];
        layer4[30][15:8] = buffer_data_0[3311:3304];
        layer4[30][23:16] = buffer_data_0[3319:3312];
        layer4[30][31:24] = buffer_data_0[3327:3320];
        layer4[30][39:32] = buffer_data_0[3335:3328];
        layer0[31][7:0] = buffer_data_4[3311:3304];
        layer0[31][15:8] = buffer_data_4[3319:3312];
        layer0[31][23:16] = buffer_data_4[3327:3320];
        layer0[31][31:24] = buffer_data_4[3335:3328];
        layer0[31][39:32] = buffer_data_4[3343:3336];
        layer1[31][7:0] = buffer_data_3[3311:3304];
        layer1[31][15:8] = buffer_data_3[3319:3312];
        layer1[31][23:16] = buffer_data_3[3327:3320];
        layer1[31][31:24] = buffer_data_3[3335:3328];
        layer1[31][39:32] = buffer_data_3[3343:3336];
        layer2[31][7:0] = buffer_data_2[3311:3304];
        layer2[31][15:8] = buffer_data_2[3319:3312];
        layer2[31][23:16] = buffer_data_2[3327:3320];
        layer2[31][31:24] = buffer_data_2[3335:3328];
        layer2[31][39:32] = buffer_data_2[3343:3336];
        layer3[31][7:0] = buffer_data_1[3311:3304];
        layer3[31][15:8] = buffer_data_1[3319:3312];
        layer3[31][23:16] = buffer_data_1[3327:3320];
        layer3[31][31:24] = buffer_data_1[3335:3328];
        layer3[31][39:32] = buffer_data_1[3343:3336];
        layer4[31][7:0] = buffer_data_0[3311:3304];
        layer4[31][15:8] = buffer_data_0[3319:3312];
        layer4[31][23:16] = buffer_data_0[3327:3320];
        layer4[31][31:24] = buffer_data_0[3335:3328];
        layer4[31][39:32] = buffer_data_0[3343:3336];
        layer0[32][7:0] = buffer_data_4[3319:3312];
        layer0[32][15:8] = buffer_data_4[3327:3320];
        layer0[32][23:16] = buffer_data_4[3335:3328];
        layer0[32][31:24] = buffer_data_4[3343:3336];
        layer0[32][39:32] = buffer_data_4[3351:3344];
        layer1[32][7:0] = buffer_data_3[3319:3312];
        layer1[32][15:8] = buffer_data_3[3327:3320];
        layer1[32][23:16] = buffer_data_3[3335:3328];
        layer1[32][31:24] = buffer_data_3[3343:3336];
        layer1[32][39:32] = buffer_data_3[3351:3344];
        layer2[32][7:0] = buffer_data_2[3319:3312];
        layer2[32][15:8] = buffer_data_2[3327:3320];
        layer2[32][23:16] = buffer_data_2[3335:3328];
        layer2[32][31:24] = buffer_data_2[3343:3336];
        layer2[32][39:32] = buffer_data_2[3351:3344];
        layer3[32][7:0] = buffer_data_1[3319:3312];
        layer3[32][15:8] = buffer_data_1[3327:3320];
        layer3[32][23:16] = buffer_data_1[3335:3328];
        layer3[32][31:24] = buffer_data_1[3343:3336];
        layer3[32][39:32] = buffer_data_1[3351:3344];
        layer4[32][7:0] = buffer_data_0[3319:3312];
        layer4[32][15:8] = buffer_data_0[3327:3320];
        layer4[32][23:16] = buffer_data_0[3335:3328];
        layer4[32][31:24] = buffer_data_0[3343:3336];
        layer4[32][39:32] = buffer_data_0[3351:3344];
        layer0[33][7:0] = buffer_data_4[3327:3320];
        layer0[33][15:8] = buffer_data_4[3335:3328];
        layer0[33][23:16] = buffer_data_4[3343:3336];
        layer0[33][31:24] = buffer_data_4[3351:3344];
        layer0[33][39:32] = buffer_data_4[3359:3352];
        layer1[33][7:0] = buffer_data_3[3327:3320];
        layer1[33][15:8] = buffer_data_3[3335:3328];
        layer1[33][23:16] = buffer_data_3[3343:3336];
        layer1[33][31:24] = buffer_data_3[3351:3344];
        layer1[33][39:32] = buffer_data_3[3359:3352];
        layer2[33][7:0] = buffer_data_2[3327:3320];
        layer2[33][15:8] = buffer_data_2[3335:3328];
        layer2[33][23:16] = buffer_data_2[3343:3336];
        layer2[33][31:24] = buffer_data_2[3351:3344];
        layer2[33][39:32] = buffer_data_2[3359:3352];
        layer3[33][7:0] = buffer_data_1[3327:3320];
        layer3[33][15:8] = buffer_data_1[3335:3328];
        layer3[33][23:16] = buffer_data_1[3343:3336];
        layer3[33][31:24] = buffer_data_1[3351:3344];
        layer3[33][39:32] = buffer_data_1[3359:3352];
        layer4[33][7:0] = buffer_data_0[3327:3320];
        layer4[33][15:8] = buffer_data_0[3335:3328];
        layer4[33][23:16] = buffer_data_0[3343:3336];
        layer4[33][31:24] = buffer_data_0[3351:3344];
        layer4[33][39:32] = buffer_data_0[3359:3352];
        layer0[34][7:0] = buffer_data_4[3335:3328];
        layer0[34][15:8] = buffer_data_4[3343:3336];
        layer0[34][23:16] = buffer_data_4[3351:3344];
        layer0[34][31:24] = buffer_data_4[3359:3352];
        layer0[34][39:32] = buffer_data_4[3367:3360];
        layer1[34][7:0] = buffer_data_3[3335:3328];
        layer1[34][15:8] = buffer_data_3[3343:3336];
        layer1[34][23:16] = buffer_data_3[3351:3344];
        layer1[34][31:24] = buffer_data_3[3359:3352];
        layer1[34][39:32] = buffer_data_3[3367:3360];
        layer2[34][7:0] = buffer_data_2[3335:3328];
        layer2[34][15:8] = buffer_data_2[3343:3336];
        layer2[34][23:16] = buffer_data_2[3351:3344];
        layer2[34][31:24] = buffer_data_2[3359:3352];
        layer2[34][39:32] = buffer_data_2[3367:3360];
        layer3[34][7:0] = buffer_data_1[3335:3328];
        layer3[34][15:8] = buffer_data_1[3343:3336];
        layer3[34][23:16] = buffer_data_1[3351:3344];
        layer3[34][31:24] = buffer_data_1[3359:3352];
        layer3[34][39:32] = buffer_data_1[3367:3360];
        layer4[34][7:0] = buffer_data_0[3335:3328];
        layer4[34][15:8] = buffer_data_0[3343:3336];
        layer4[34][23:16] = buffer_data_0[3351:3344];
        layer4[34][31:24] = buffer_data_0[3359:3352];
        layer4[34][39:32] = buffer_data_0[3367:3360];
        layer0[35][7:0] = buffer_data_4[3343:3336];
        layer0[35][15:8] = buffer_data_4[3351:3344];
        layer0[35][23:16] = buffer_data_4[3359:3352];
        layer0[35][31:24] = buffer_data_4[3367:3360];
        layer0[35][39:32] = buffer_data_4[3375:3368];
        layer1[35][7:0] = buffer_data_3[3343:3336];
        layer1[35][15:8] = buffer_data_3[3351:3344];
        layer1[35][23:16] = buffer_data_3[3359:3352];
        layer1[35][31:24] = buffer_data_3[3367:3360];
        layer1[35][39:32] = buffer_data_3[3375:3368];
        layer2[35][7:0] = buffer_data_2[3343:3336];
        layer2[35][15:8] = buffer_data_2[3351:3344];
        layer2[35][23:16] = buffer_data_2[3359:3352];
        layer2[35][31:24] = buffer_data_2[3367:3360];
        layer2[35][39:32] = buffer_data_2[3375:3368];
        layer3[35][7:0] = buffer_data_1[3343:3336];
        layer3[35][15:8] = buffer_data_1[3351:3344];
        layer3[35][23:16] = buffer_data_1[3359:3352];
        layer3[35][31:24] = buffer_data_1[3367:3360];
        layer3[35][39:32] = buffer_data_1[3375:3368];
        layer4[35][7:0] = buffer_data_0[3343:3336];
        layer4[35][15:8] = buffer_data_0[3351:3344];
        layer4[35][23:16] = buffer_data_0[3359:3352];
        layer4[35][31:24] = buffer_data_0[3367:3360];
        layer4[35][39:32] = buffer_data_0[3375:3368];
        layer0[36][7:0] = buffer_data_4[3351:3344];
        layer0[36][15:8] = buffer_data_4[3359:3352];
        layer0[36][23:16] = buffer_data_4[3367:3360];
        layer0[36][31:24] = buffer_data_4[3375:3368];
        layer0[36][39:32] = buffer_data_4[3383:3376];
        layer1[36][7:0] = buffer_data_3[3351:3344];
        layer1[36][15:8] = buffer_data_3[3359:3352];
        layer1[36][23:16] = buffer_data_3[3367:3360];
        layer1[36][31:24] = buffer_data_3[3375:3368];
        layer1[36][39:32] = buffer_data_3[3383:3376];
        layer2[36][7:0] = buffer_data_2[3351:3344];
        layer2[36][15:8] = buffer_data_2[3359:3352];
        layer2[36][23:16] = buffer_data_2[3367:3360];
        layer2[36][31:24] = buffer_data_2[3375:3368];
        layer2[36][39:32] = buffer_data_2[3383:3376];
        layer3[36][7:0] = buffer_data_1[3351:3344];
        layer3[36][15:8] = buffer_data_1[3359:3352];
        layer3[36][23:16] = buffer_data_1[3367:3360];
        layer3[36][31:24] = buffer_data_1[3375:3368];
        layer3[36][39:32] = buffer_data_1[3383:3376];
        layer4[36][7:0] = buffer_data_0[3351:3344];
        layer4[36][15:8] = buffer_data_0[3359:3352];
        layer4[36][23:16] = buffer_data_0[3367:3360];
        layer4[36][31:24] = buffer_data_0[3375:3368];
        layer4[36][39:32] = buffer_data_0[3383:3376];
        layer0[37][7:0] = buffer_data_4[3359:3352];
        layer0[37][15:8] = buffer_data_4[3367:3360];
        layer0[37][23:16] = buffer_data_4[3375:3368];
        layer0[37][31:24] = buffer_data_4[3383:3376];
        layer0[37][39:32] = buffer_data_4[3391:3384];
        layer1[37][7:0] = buffer_data_3[3359:3352];
        layer1[37][15:8] = buffer_data_3[3367:3360];
        layer1[37][23:16] = buffer_data_3[3375:3368];
        layer1[37][31:24] = buffer_data_3[3383:3376];
        layer1[37][39:32] = buffer_data_3[3391:3384];
        layer2[37][7:0] = buffer_data_2[3359:3352];
        layer2[37][15:8] = buffer_data_2[3367:3360];
        layer2[37][23:16] = buffer_data_2[3375:3368];
        layer2[37][31:24] = buffer_data_2[3383:3376];
        layer2[37][39:32] = buffer_data_2[3391:3384];
        layer3[37][7:0] = buffer_data_1[3359:3352];
        layer3[37][15:8] = buffer_data_1[3367:3360];
        layer3[37][23:16] = buffer_data_1[3375:3368];
        layer3[37][31:24] = buffer_data_1[3383:3376];
        layer3[37][39:32] = buffer_data_1[3391:3384];
        layer4[37][7:0] = buffer_data_0[3359:3352];
        layer4[37][15:8] = buffer_data_0[3367:3360];
        layer4[37][23:16] = buffer_data_0[3375:3368];
        layer4[37][31:24] = buffer_data_0[3383:3376];
        layer4[37][39:32] = buffer_data_0[3391:3384];
        layer0[38][7:0] = buffer_data_4[3367:3360];
        layer0[38][15:8] = buffer_data_4[3375:3368];
        layer0[38][23:16] = buffer_data_4[3383:3376];
        layer0[38][31:24] = buffer_data_4[3391:3384];
        layer0[38][39:32] = buffer_data_4[3399:3392];
        layer1[38][7:0] = buffer_data_3[3367:3360];
        layer1[38][15:8] = buffer_data_3[3375:3368];
        layer1[38][23:16] = buffer_data_3[3383:3376];
        layer1[38][31:24] = buffer_data_3[3391:3384];
        layer1[38][39:32] = buffer_data_3[3399:3392];
        layer2[38][7:0] = buffer_data_2[3367:3360];
        layer2[38][15:8] = buffer_data_2[3375:3368];
        layer2[38][23:16] = buffer_data_2[3383:3376];
        layer2[38][31:24] = buffer_data_2[3391:3384];
        layer2[38][39:32] = buffer_data_2[3399:3392];
        layer3[38][7:0] = buffer_data_1[3367:3360];
        layer3[38][15:8] = buffer_data_1[3375:3368];
        layer3[38][23:16] = buffer_data_1[3383:3376];
        layer3[38][31:24] = buffer_data_1[3391:3384];
        layer3[38][39:32] = buffer_data_1[3399:3392];
        layer4[38][7:0] = buffer_data_0[3367:3360];
        layer4[38][15:8] = buffer_data_0[3375:3368];
        layer4[38][23:16] = buffer_data_0[3383:3376];
        layer4[38][31:24] = buffer_data_0[3391:3384];
        layer4[38][39:32] = buffer_data_0[3399:3392];
        layer0[39][7:0] = buffer_data_4[3375:3368];
        layer0[39][15:8] = buffer_data_4[3383:3376];
        layer0[39][23:16] = buffer_data_4[3391:3384];
        layer0[39][31:24] = buffer_data_4[3399:3392];
        layer0[39][39:32] = buffer_data_4[3407:3400];
        layer1[39][7:0] = buffer_data_3[3375:3368];
        layer1[39][15:8] = buffer_data_3[3383:3376];
        layer1[39][23:16] = buffer_data_3[3391:3384];
        layer1[39][31:24] = buffer_data_3[3399:3392];
        layer1[39][39:32] = buffer_data_3[3407:3400];
        layer2[39][7:0] = buffer_data_2[3375:3368];
        layer2[39][15:8] = buffer_data_2[3383:3376];
        layer2[39][23:16] = buffer_data_2[3391:3384];
        layer2[39][31:24] = buffer_data_2[3399:3392];
        layer2[39][39:32] = buffer_data_2[3407:3400];
        layer3[39][7:0] = buffer_data_1[3375:3368];
        layer3[39][15:8] = buffer_data_1[3383:3376];
        layer3[39][23:16] = buffer_data_1[3391:3384];
        layer3[39][31:24] = buffer_data_1[3399:3392];
        layer3[39][39:32] = buffer_data_1[3407:3400];
        layer4[39][7:0] = buffer_data_0[3375:3368];
        layer4[39][15:8] = buffer_data_0[3383:3376];
        layer4[39][23:16] = buffer_data_0[3391:3384];
        layer4[39][31:24] = buffer_data_0[3399:3392];
        layer4[39][39:32] = buffer_data_0[3407:3400];
        layer0[40][7:0] = buffer_data_4[3383:3376];
        layer0[40][15:8] = buffer_data_4[3391:3384];
        layer0[40][23:16] = buffer_data_4[3399:3392];
        layer0[40][31:24] = buffer_data_4[3407:3400];
        layer0[40][39:32] = buffer_data_4[3415:3408];
        layer1[40][7:0] = buffer_data_3[3383:3376];
        layer1[40][15:8] = buffer_data_3[3391:3384];
        layer1[40][23:16] = buffer_data_3[3399:3392];
        layer1[40][31:24] = buffer_data_3[3407:3400];
        layer1[40][39:32] = buffer_data_3[3415:3408];
        layer2[40][7:0] = buffer_data_2[3383:3376];
        layer2[40][15:8] = buffer_data_2[3391:3384];
        layer2[40][23:16] = buffer_data_2[3399:3392];
        layer2[40][31:24] = buffer_data_2[3407:3400];
        layer2[40][39:32] = buffer_data_2[3415:3408];
        layer3[40][7:0] = buffer_data_1[3383:3376];
        layer3[40][15:8] = buffer_data_1[3391:3384];
        layer3[40][23:16] = buffer_data_1[3399:3392];
        layer3[40][31:24] = buffer_data_1[3407:3400];
        layer3[40][39:32] = buffer_data_1[3415:3408];
        layer4[40][7:0] = buffer_data_0[3383:3376];
        layer4[40][15:8] = buffer_data_0[3391:3384];
        layer4[40][23:16] = buffer_data_0[3399:3392];
        layer4[40][31:24] = buffer_data_0[3407:3400];
        layer4[40][39:32] = buffer_data_0[3415:3408];
        layer0[41][7:0] = buffer_data_4[3391:3384];
        layer0[41][15:8] = buffer_data_4[3399:3392];
        layer0[41][23:16] = buffer_data_4[3407:3400];
        layer0[41][31:24] = buffer_data_4[3415:3408];
        layer0[41][39:32] = buffer_data_4[3423:3416];
        layer1[41][7:0] = buffer_data_3[3391:3384];
        layer1[41][15:8] = buffer_data_3[3399:3392];
        layer1[41][23:16] = buffer_data_3[3407:3400];
        layer1[41][31:24] = buffer_data_3[3415:3408];
        layer1[41][39:32] = buffer_data_3[3423:3416];
        layer2[41][7:0] = buffer_data_2[3391:3384];
        layer2[41][15:8] = buffer_data_2[3399:3392];
        layer2[41][23:16] = buffer_data_2[3407:3400];
        layer2[41][31:24] = buffer_data_2[3415:3408];
        layer2[41][39:32] = buffer_data_2[3423:3416];
        layer3[41][7:0] = buffer_data_1[3391:3384];
        layer3[41][15:8] = buffer_data_1[3399:3392];
        layer3[41][23:16] = buffer_data_1[3407:3400];
        layer3[41][31:24] = buffer_data_1[3415:3408];
        layer3[41][39:32] = buffer_data_1[3423:3416];
        layer4[41][7:0] = buffer_data_0[3391:3384];
        layer4[41][15:8] = buffer_data_0[3399:3392];
        layer4[41][23:16] = buffer_data_0[3407:3400];
        layer4[41][31:24] = buffer_data_0[3415:3408];
        layer4[41][39:32] = buffer_data_0[3423:3416];
        layer0[42][7:0] = buffer_data_4[3399:3392];
        layer0[42][15:8] = buffer_data_4[3407:3400];
        layer0[42][23:16] = buffer_data_4[3415:3408];
        layer0[42][31:24] = buffer_data_4[3423:3416];
        layer0[42][39:32] = buffer_data_4[3431:3424];
        layer1[42][7:0] = buffer_data_3[3399:3392];
        layer1[42][15:8] = buffer_data_3[3407:3400];
        layer1[42][23:16] = buffer_data_3[3415:3408];
        layer1[42][31:24] = buffer_data_3[3423:3416];
        layer1[42][39:32] = buffer_data_3[3431:3424];
        layer2[42][7:0] = buffer_data_2[3399:3392];
        layer2[42][15:8] = buffer_data_2[3407:3400];
        layer2[42][23:16] = buffer_data_2[3415:3408];
        layer2[42][31:24] = buffer_data_2[3423:3416];
        layer2[42][39:32] = buffer_data_2[3431:3424];
        layer3[42][7:0] = buffer_data_1[3399:3392];
        layer3[42][15:8] = buffer_data_1[3407:3400];
        layer3[42][23:16] = buffer_data_1[3415:3408];
        layer3[42][31:24] = buffer_data_1[3423:3416];
        layer3[42][39:32] = buffer_data_1[3431:3424];
        layer4[42][7:0] = buffer_data_0[3399:3392];
        layer4[42][15:8] = buffer_data_0[3407:3400];
        layer4[42][23:16] = buffer_data_0[3415:3408];
        layer4[42][31:24] = buffer_data_0[3423:3416];
        layer4[42][39:32] = buffer_data_0[3431:3424];
        layer0[43][7:0] = buffer_data_4[3407:3400];
        layer0[43][15:8] = buffer_data_4[3415:3408];
        layer0[43][23:16] = buffer_data_4[3423:3416];
        layer0[43][31:24] = buffer_data_4[3431:3424];
        layer0[43][39:32] = buffer_data_4[3439:3432];
        layer1[43][7:0] = buffer_data_3[3407:3400];
        layer1[43][15:8] = buffer_data_3[3415:3408];
        layer1[43][23:16] = buffer_data_3[3423:3416];
        layer1[43][31:24] = buffer_data_3[3431:3424];
        layer1[43][39:32] = buffer_data_3[3439:3432];
        layer2[43][7:0] = buffer_data_2[3407:3400];
        layer2[43][15:8] = buffer_data_2[3415:3408];
        layer2[43][23:16] = buffer_data_2[3423:3416];
        layer2[43][31:24] = buffer_data_2[3431:3424];
        layer2[43][39:32] = buffer_data_2[3439:3432];
        layer3[43][7:0] = buffer_data_1[3407:3400];
        layer3[43][15:8] = buffer_data_1[3415:3408];
        layer3[43][23:16] = buffer_data_1[3423:3416];
        layer3[43][31:24] = buffer_data_1[3431:3424];
        layer3[43][39:32] = buffer_data_1[3439:3432];
        layer4[43][7:0] = buffer_data_0[3407:3400];
        layer4[43][15:8] = buffer_data_0[3415:3408];
        layer4[43][23:16] = buffer_data_0[3423:3416];
        layer4[43][31:24] = buffer_data_0[3431:3424];
        layer4[43][39:32] = buffer_data_0[3439:3432];
        layer0[44][7:0] = buffer_data_4[3415:3408];
        layer0[44][15:8] = buffer_data_4[3423:3416];
        layer0[44][23:16] = buffer_data_4[3431:3424];
        layer0[44][31:24] = buffer_data_4[3439:3432];
        layer0[44][39:32] = buffer_data_4[3447:3440];
        layer1[44][7:0] = buffer_data_3[3415:3408];
        layer1[44][15:8] = buffer_data_3[3423:3416];
        layer1[44][23:16] = buffer_data_3[3431:3424];
        layer1[44][31:24] = buffer_data_3[3439:3432];
        layer1[44][39:32] = buffer_data_3[3447:3440];
        layer2[44][7:0] = buffer_data_2[3415:3408];
        layer2[44][15:8] = buffer_data_2[3423:3416];
        layer2[44][23:16] = buffer_data_2[3431:3424];
        layer2[44][31:24] = buffer_data_2[3439:3432];
        layer2[44][39:32] = buffer_data_2[3447:3440];
        layer3[44][7:0] = buffer_data_1[3415:3408];
        layer3[44][15:8] = buffer_data_1[3423:3416];
        layer3[44][23:16] = buffer_data_1[3431:3424];
        layer3[44][31:24] = buffer_data_1[3439:3432];
        layer3[44][39:32] = buffer_data_1[3447:3440];
        layer4[44][7:0] = buffer_data_0[3415:3408];
        layer4[44][15:8] = buffer_data_0[3423:3416];
        layer4[44][23:16] = buffer_data_0[3431:3424];
        layer4[44][31:24] = buffer_data_0[3439:3432];
        layer4[44][39:32] = buffer_data_0[3447:3440];
        layer0[45][7:0] = buffer_data_4[3423:3416];
        layer0[45][15:8] = buffer_data_4[3431:3424];
        layer0[45][23:16] = buffer_data_4[3439:3432];
        layer0[45][31:24] = buffer_data_4[3447:3440];
        layer0[45][39:32] = buffer_data_4[3455:3448];
        layer1[45][7:0] = buffer_data_3[3423:3416];
        layer1[45][15:8] = buffer_data_3[3431:3424];
        layer1[45][23:16] = buffer_data_3[3439:3432];
        layer1[45][31:24] = buffer_data_3[3447:3440];
        layer1[45][39:32] = buffer_data_3[3455:3448];
        layer2[45][7:0] = buffer_data_2[3423:3416];
        layer2[45][15:8] = buffer_data_2[3431:3424];
        layer2[45][23:16] = buffer_data_2[3439:3432];
        layer2[45][31:24] = buffer_data_2[3447:3440];
        layer2[45][39:32] = buffer_data_2[3455:3448];
        layer3[45][7:0] = buffer_data_1[3423:3416];
        layer3[45][15:8] = buffer_data_1[3431:3424];
        layer3[45][23:16] = buffer_data_1[3439:3432];
        layer3[45][31:24] = buffer_data_1[3447:3440];
        layer3[45][39:32] = buffer_data_1[3455:3448];
        layer4[45][7:0] = buffer_data_0[3423:3416];
        layer4[45][15:8] = buffer_data_0[3431:3424];
        layer4[45][23:16] = buffer_data_0[3439:3432];
        layer4[45][31:24] = buffer_data_0[3447:3440];
        layer4[45][39:32] = buffer_data_0[3455:3448];
        layer0[46][7:0] = buffer_data_4[3431:3424];
        layer0[46][15:8] = buffer_data_4[3439:3432];
        layer0[46][23:16] = buffer_data_4[3447:3440];
        layer0[46][31:24] = buffer_data_4[3455:3448];
        layer0[46][39:32] = buffer_data_4[3463:3456];
        layer1[46][7:0] = buffer_data_3[3431:3424];
        layer1[46][15:8] = buffer_data_3[3439:3432];
        layer1[46][23:16] = buffer_data_3[3447:3440];
        layer1[46][31:24] = buffer_data_3[3455:3448];
        layer1[46][39:32] = buffer_data_3[3463:3456];
        layer2[46][7:0] = buffer_data_2[3431:3424];
        layer2[46][15:8] = buffer_data_2[3439:3432];
        layer2[46][23:16] = buffer_data_2[3447:3440];
        layer2[46][31:24] = buffer_data_2[3455:3448];
        layer2[46][39:32] = buffer_data_2[3463:3456];
        layer3[46][7:0] = buffer_data_1[3431:3424];
        layer3[46][15:8] = buffer_data_1[3439:3432];
        layer3[46][23:16] = buffer_data_1[3447:3440];
        layer3[46][31:24] = buffer_data_1[3455:3448];
        layer3[46][39:32] = buffer_data_1[3463:3456];
        layer4[46][7:0] = buffer_data_0[3431:3424];
        layer4[46][15:8] = buffer_data_0[3439:3432];
        layer4[46][23:16] = buffer_data_0[3447:3440];
        layer4[46][31:24] = buffer_data_0[3455:3448];
        layer4[46][39:32] = buffer_data_0[3463:3456];
        layer0[47][7:0] = buffer_data_4[3439:3432];
        layer0[47][15:8] = buffer_data_4[3447:3440];
        layer0[47][23:16] = buffer_data_4[3455:3448];
        layer0[47][31:24] = buffer_data_4[3463:3456];
        layer0[47][39:32] = buffer_data_4[3471:3464];
        layer1[47][7:0] = buffer_data_3[3439:3432];
        layer1[47][15:8] = buffer_data_3[3447:3440];
        layer1[47][23:16] = buffer_data_3[3455:3448];
        layer1[47][31:24] = buffer_data_3[3463:3456];
        layer1[47][39:32] = buffer_data_3[3471:3464];
        layer2[47][7:0] = buffer_data_2[3439:3432];
        layer2[47][15:8] = buffer_data_2[3447:3440];
        layer2[47][23:16] = buffer_data_2[3455:3448];
        layer2[47][31:24] = buffer_data_2[3463:3456];
        layer2[47][39:32] = buffer_data_2[3471:3464];
        layer3[47][7:0] = buffer_data_1[3439:3432];
        layer3[47][15:8] = buffer_data_1[3447:3440];
        layer3[47][23:16] = buffer_data_1[3455:3448];
        layer3[47][31:24] = buffer_data_1[3463:3456];
        layer3[47][39:32] = buffer_data_1[3471:3464];
        layer4[47][7:0] = buffer_data_0[3439:3432];
        layer4[47][15:8] = buffer_data_0[3447:3440];
        layer4[47][23:16] = buffer_data_0[3455:3448];
        layer4[47][31:24] = buffer_data_0[3463:3456];
        layer4[47][39:32] = buffer_data_0[3471:3464];
        layer0[48][7:0] = buffer_data_4[3447:3440];
        layer0[48][15:8] = buffer_data_4[3455:3448];
        layer0[48][23:16] = buffer_data_4[3463:3456];
        layer0[48][31:24] = buffer_data_4[3471:3464];
        layer0[48][39:32] = buffer_data_4[3479:3472];
        layer1[48][7:0] = buffer_data_3[3447:3440];
        layer1[48][15:8] = buffer_data_3[3455:3448];
        layer1[48][23:16] = buffer_data_3[3463:3456];
        layer1[48][31:24] = buffer_data_3[3471:3464];
        layer1[48][39:32] = buffer_data_3[3479:3472];
        layer2[48][7:0] = buffer_data_2[3447:3440];
        layer2[48][15:8] = buffer_data_2[3455:3448];
        layer2[48][23:16] = buffer_data_2[3463:3456];
        layer2[48][31:24] = buffer_data_2[3471:3464];
        layer2[48][39:32] = buffer_data_2[3479:3472];
        layer3[48][7:0] = buffer_data_1[3447:3440];
        layer3[48][15:8] = buffer_data_1[3455:3448];
        layer3[48][23:16] = buffer_data_1[3463:3456];
        layer3[48][31:24] = buffer_data_1[3471:3464];
        layer3[48][39:32] = buffer_data_1[3479:3472];
        layer4[48][7:0] = buffer_data_0[3447:3440];
        layer4[48][15:8] = buffer_data_0[3455:3448];
        layer4[48][23:16] = buffer_data_0[3463:3456];
        layer4[48][31:24] = buffer_data_0[3471:3464];
        layer4[48][39:32] = buffer_data_0[3479:3472];
        layer0[49][7:0] = buffer_data_4[3455:3448];
        layer0[49][15:8] = buffer_data_4[3463:3456];
        layer0[49][23:16] = buffer_data_4[3471:3464];
        layer0[49][31:24] = buffer_data_4[3479:3472];
        layer0[49][39:32] = buffer_data_4[3487:3480];
        layer1[49][7:0] = buffer_data_3[3455:3448];
        layer1[49][15:8] = buffer_data_3[3463:3456];
        layer1[49][23:16] = buffer_data_3[3471:3464];
        layer1[49][31:24] = buffer_data_3[3479:3472];
        layer1[49][39:32] = buffer_data_3[3487:3480];
        layer2[49][7:0] = buffer_data_2[3455:3448];
        layer2[49][15:8] = buffer_data_2[3463:3456];
        layer2[49][23:16] = buffer_data_2[3471:3464];
        layer2[49][31:24] = buffer_data_2[3479:3472];
        layer2[49][39:32] = buffer_data_2[3487:3480];
        layer3[49][7:0] = buffer_data_1[3455:3448];
        layer3[49][15:8] = buffer_data_1[3463:3456];
        layer3[49][23:16] = buffer_data_1[3471:3464];
        layer3[49][31:24] = buffer_data_1[3479:3472];
        layer3[49][39:32] = buffer_data_1[3487:3480];
        layer4[49][7:0] = buffer_data_0[3455:3448];
        layer4[49][15:8] = buffer_data_0[3463:3456];
        layer4[49][23:16] = buffer_data_0[3471:3464];
        layer4[49][31:24] = buffer_data_0[3479:3472];
        layer4[49][39:32] = buffer_data_0[3487:3480];
        layer0[50][7:0] = buffer_data_4[3463:3456];
        layer0[50][15:8] = buffer_data_4[3471:3464];
        layer0[50][23:16] = buffer_data_4[3479:3472];
        layer0[50][31:24] = buffer_data_4[3487:3480];
        layer0[50][39:32] = buffer_data_4[3495:3488];
        layer1[50][7:0] = buffer_data_3[3463:3456];
        layer1[50][15:8] = buffer_data_3[3471:3464];
        layer1[50][23:16] = buffer_data_3[3479:3472];
        layer1[50][31:24] = buffer_data_3[3487:3480];
        layer1[50][39:32] = buffer_data_3[3495:3488];
        layer2[50][7:0] = buffer_data_2[3463:3456];
        layer2[50][15:8] = buffer_data_2[3471:3464];
        layer2[50][23:16] = buffer_data_2[3479:3472];
        layer2[50][31:24] = buffer_data_2[3487:3480];
        layer2[50][39:32] = buffer_data_2[3495:3488];
        layer3[50][7:0] = buffer_data_1[3463:3456];
        layer3[50][15:8] = buffer_data_1[3471:3464];
        layer3[50][23:16] = buffer_data_1[3479:3472];
        layer3[50][31:24] = buffer_data_1[3487:3480];
        layer3[50][39:32] = buffer_data_1[3495:3488];
        layer4[50][7:0] = buffer_data_0[3463:3456];
        layer4[50][15:8] = buffer_data_0[3471:3464];
        layer4[50][23:16] = buffer_data_0[3479:3472];
        layer4[50][31:24] = buffer_data_0[3487:3480];
        layer4[50][39:32] = buffer_data_0[3495:3488];
        layer0[51][7:0] = buffer_data_4[3471:3464];
        layer0[51][15:8] = buffer_data_4[3479:3472];
        layer0[51][23:16] = buffer_data_4[3487:3480];
        layer0[51][31:24] = buffer_data_4[3495:3488];
        layer0[51][39:32] = buffer_data_4[3503:3496];
        layer1[51][7:0] = buffer_data_3[3471:3464];
        layer1[51][15:8] = buffer_data_3[3479:3472];
        layer1[51][23:16] = buffer_data_3[3487:3480];
        layer1[51][31:24] = buffer_data_3[3495:3488];
        layer1[51][39:32] = buffer_data_3[3503:3496];
        layer2[51][7:0] = buffer_data_2[3471:3464];
        layer2[51][15:8] = buffer_data_2[3479:3472];
        layer2[51][23:16] = buffer_data_2[3487:3480];
        layer2[51][31:24] = buffer_data_2[3495:3488];
        layer2[51][39:32] = buffer_data_2[3503:3496];
        layer3[51][7:0] = buffer_data_1[3471:3464];
        layer3[51][15:8] = buffer_data_1[3479:3472];
        layer3[51][23:16] = buffer_data_1[3487:3480];
        layer3[51][31:24] = buffer_data_1[3495:3488];
        layer3[51][39:32] = buffer_data_1[3503:3496];
        layer4[51][7:0] = buffer_data_0[3471:3464];
        layer4[51][15:8] = buffer_data_0[3479:3472];
        layer4[51][23:16] = buffer_data_0[3487:3480];
        layer4[51][31:24] = buffer_data_0[3495:3488];
        layer4[51][39:32] = buffer_data_0[3503:3496];
        layer0[52][7:0] = buffer_data_4[3479:3472];
        layer0[52][15:8] = buffer_data_4[3487:3480];
        layer0[52][23:16] = buffer_data_4[3495:3488];
        layer0[52][31:24] = buffer_data_4[3503:3496];
        layer0[52][39:32] = buffer_data_4[3511:3504];
        layer1[52][7:0] = buffer_data_3[3479:3472];
        layer1[52][15:8] = buffer_data_3[3487:3480];
        layer1[52][23:16] = buffer_data_3[3495:3488];
        layer1[52][31:24] = buffer_data_3[3503:3496];
        layer1[52][39:32] = buffer_data_3[3511:3504];
        layer2[52][7:0] = buffer_data_2[3479:3472];
        layer2[52][15:8] = buffer_data_2[3487:3480];
        layer2[52][23:16] = buffer_data_2[3495:3488];
        layer2[52][31:24] = buffer_data_2[3503:3496];
        layer2[52][39:32] = buffer_data_2[3511:3504];
        layer3[52][7:0] = buffer_data_1[3479:3472];
        layer3[52][15:8] = buffer_data_1[3487:3480];
        layer3[52][23:16] = buffer_data_1[3495:3488];
        layer3[52][31:24] = buffer_data_1[3503:3496];
        layer3[52][39:32] = buffer_data_1[3511:3504];
        layer4[52][7:0] = buffer_data_0[3479:3472];
        layer4[52][15:8] = buffer_data_0[3487:3480];
        layer4[52][23:16] = buffer_data_0[3495:3488];
        layer4[52][31:24] = buffer_data_0[3503:3496];
        layer4[52][39:32] = buffer_data_0[3511:3504];
        layer0[53][7:0] = buffer_data_4[3487:3480];
        layer0[53][15:8] = buffer_data_4[3495:3488];
        layer0[53][23:16] = buffer_data_4[3503:3496];
        layer0[53][31:24] = buffer_data_4[3511:3504];
        layer0[53][39:32] = buffer_data_4[3519:3512];
        layer1[53][7:0] = buffer_data_3[3487:3480];
        layer1[53][15:8] = buffer_data_3[3495:3488];
        layer1[53][23:16] = buffer_data_3[3503:3496];
        layer1[53][31:24] = buffer_data_3[3511:3504];
        layer1[53][39:32] = buffer_data_3[3519:3512];
        layer2[53][7:0] = buffer_data_2[3487:3480];
        layer2[53][15:8] = buffer_data_2[3495:3488];
        layer2[53][23:16] = buffer_data_2[3503:3496];
        layer2[53][31:24] = buffer_data_2[3511:3504];
        layer2[53][39:32] = buffer_data_2[3519:3512];
        layer3[53][7:0] = buffer_data_1[3487:3480];
        layer3[53][15:8] = buffer_data_1[3495:3488];
        layer3[53][23:16] = buffer_data_1[3503:3496];
        layer3[53][31:24] = buffer_data_1[3511:3504];
        layer3[53][39:32] = buffer_data_1[3519:3512];
        layer4[53][7:0] = buffer_data_0[3487:3480];
        layer4[53][15:8] = buffer_data_0[3495:3488];
        layer4[53][23:16] = buffer_data_0[3503:3496];
        layer4[53][31:24] = buffer_data_0[3511:3504];
        layer4[53][39:32] = buffer_data_0[3519:3512];
        layer0[54][7:0] = buffer_data_4[3495:3488];
        layer0[54][15:8] = buffer_data_4[3503:3496];
        layer0[54][23:16] = buffer_data_4[3511:3504];
        layer0[54][31:24] = buffer_data_4[3519:3512];
        layer0[54][39:32] = buffer_data_4[3527:3520];
        layer1[54][7:0] = buffer_data_3[3495:3488];
        layer1[54][15:8] = buffer_data_3[3503:3496];
        layer1[54][23:16] = buffer_data_3[3511:3504];
        layer1[54][31:24] = buffer_data_3[3519:3512];
        layer1[54][39:32] = buffer_data_3[3527:3520];
        layer2[54][7:0] = buffer_data_2[3495:3488];
        layer2[54][15:8] = buffer_data_2[3503:3496];
        layer2[54][23:16] = buffer_data_2[3511:3504];
        layer2[54][31:24] = buffer_data_2[3519:3512];
        layer2[54][39:32] = buffer_data_2[3527:3520];
        layer3[54][7:0] = buffer_data_1[3495:3488];
        layer3[54][15:8] = buffer_data_1[3503:3496];
        layer3[54][23:16] = buffer_data_1[3511:3504];
        layer3[54][31:24] = buffer_data_1[3519:3512];
        layer3[54][39:32] = buffer_data_1[3527:3520];
        layer4[54][7:0] = buffer_data_0[3495:3488];
        layer4[54][15:8] = buffer_data_0[3503:3496];
        layer4[54][23:16] = buffer_data_0[3511:3504];
        layer4[54][31:24] = buffer_data_0[3519:3512];
        layer4[54][39:32] = buffer_data_0[3527:3520];
        layer0[55][7:0] = buffer_data_4[3503:3496];
        layer0[55][15:8] = buffer_data_4[3511:3504];
        layer0[55][23:16] = buffer_data_4[3519:3512];
        layer0[55][31:24] = buffer_data_4[3527:3520];
        layer0[55][39:32] = buffer_data_4[3535:3528];
        layer1[55][7:0] = buffer_data_3[3503:3496];
        layer1[55][15:8] = buffer_data_3[3511:3504];
        layer1[55][23:16] = buffer_data_3[3519:3512];
        layer1[55][31:24] = buffer_data_3[3527:3520];
        layer1[55][39:32] = buffer_data_3[3535:3528];
        layer2[55][7:0] = buffer_data_2[3503:3496];
        layer2[55][15:8] = buffer_data_2[3511:3504];
        layer2[55][23:16] = buffer_data_2[3519:3512];
        layer2[55][31:24] = buffer_data_2[3527:3520];
        layer2[55][39:32] = buffer_data_2[3535:3528];
        layer3[55][7:0] = buffer_data_1[3503:3496];
        layer3[55][15:8] = buffer_data_1[3511:3504];
        layer3[55][23:16] = buffer_data_1[3519:3512];
        layer3[55][31:24] = buffer_data_1[3527:3520];
        layer3[55][39:32] = buffer_data_1[3535:3528];
        layer4[55][7:0] = buffer_data_0[3503:3496];
        layer4[55][15:8] = buffer_data_0[3511:3504];
        layer4[55][23:16] = buffer_data_0[3519:3512];
        layer4[55][31:24] = buffer_data_0[3527:3520];
        layer4[55][39:32] = buffer_data_0[3535:3528];
        layer0[56][7:0] = buffer_data_4[3511:3504];
        layer0[56][15:8] = buffer_data_4[3519:3512];
        layer0[56][23:16] = buffer_data_4[3527:3520];
        layer0[56][31:24] = buffer_data_4[3535:3528];
        layer0[56][39:32] = buffer_data_4[3543:3536];
        layer1[56][7:0] = buffer_data_3[3511:3504];
        layer1[56][15:8] = buffer_data_3[3519:3512];
        layer1[56][23:16] = buffer_data_3[3527:3520];
        layer1[56][31:24] = buffer_data_3[3535:3528];
        layer1[56][39:32] = buffer_data_3[3543:3536];
        layer2[56][7:0] = buffer_data_2[3511:3504];
        layer2[56][15:8] = buffer_data_2[3519:3512];
        layer2[56][23:16] = buffer_data_2[3527:3520];
        layer2[56][31:24] = buffer_data_2[3535:3528];
        layer2[56][39:32] = buffer_data_2[3543:3536];
        layer3[56][7:0] = buffer_data_1[3511:3504];
        layer3[56][15:8] = buffer_data_1[3519:3512];
        layer3[56][23:16] = buffer_data_1[3527:3520];
        layer3[56][31:24] = buffer_data_1[3535:3528];
        layer3[56][39:32] = buffer_data_1[3543:3536];
        layer4[56][7:0] = buffer_data_0[3511:3504];
        layer4[56][15:8] = buffer_data_0[3519:3512];
        layer4[56][23:16] = buffer_data_0[3527:3520];
        layer4[56][31:24] = buffer_data_0[3535:3528];
        layer4[56][39:32] = buffer_data_0[3543:3536];
        layer0[57][7:0] = buffer_data_4[3519:3512];
        layer0[57][15:8] = buffer_data_4[3527:3520];
        layer0[57][23:16] = buffer_data_4[3535:3528];
        layer0[57][31:24] = buffer_data_4[3543:3536];
        layer0[57][39:32] = buffer_data_4[3551:3544];
        layer1[57][7:0] = buffer_data_3[3519:3512];
        layer1[57][15:8] = buffer_data_3[3527:3520];
        layer1[57][23:16] = buffer_data_3[3535:3528];
        layer1[57][31:24] = buffer_data_3[3543:3536];
        layer1[57][39:32] = buffer_data_3[3551:3544];
        layer2[57][7:0] = buffer_data_2[3519:3512];
        layer2[57][15:8] = buffer_data_2[3527:3520];
        layer2[57][23:16] = buffer_data_2[3535:3528];
        layer2[57][31:24] = buffer_data_2[3543:3536];
        layer2[57][39:32] = buffer_data_2[3551:3544];
        layer3[57][7:0] = buffer_data_1[3519:3512];
        layer3[57][15:8] = buffer_data_1[3527:3520];
        layer3[57][23:16] = buffer_data_1[3535:3528];
        layer3[57][31:24] = buffer_data_1[3543:3536];
        layer3[57][39:32] = buffer_data_1[3551:3544];
        layer4[57][7:0] = buffer_data_0[3519:3512];
        layer4[57][15:8] = buffer_data_0[3527:3520];
        layer4[57][23:16] = buffer_data_0[3535:3528];
        layer4[57][31:24] = buffer_data_0[3543:3536];
        layer4[57][39:32] = buffer_data_0[3551:3544];
        layer0[58][7:0] = buffer_data_4[3527:3520];
        layer0[58][15:8] = buffer_data_4[3535:3528];
        layer0[58][23:16] = buffer_data_4[3543:3536];
        layer0[58][31:24] = buffer_data_4[3551:3544];
        layer0[58][39:32] = buffer_data_4[3559:3552];
        layer1[58][7:0] = buffer_data_3[3527:3520];
        layer1[58][15:8] = buffer_data_3[3535:3528];
        layer1[58][23:16] = buffer_data_3[3543:3536];
        layer1[58][31:24] = buffer_data_3[3551:3544];
        layer1[58][39:32] = buffer_data_3[3559:3552];
        layer2[58][7:0] = buffer_data_2[3527:3520];
        layer2[58][15:8] = buffer_data_2[3535:3528];
        layer2[58][23:16] = buffer_data_2[3543:3536];
        layer2[58][31:24] = buffer_data_2[3551:3544];
        layer2[58][39:32] = buffer_data_2[3559:3552];
        layer3[58][7:0] = buffer_data_1[3527:3520];
        layer3[58][15:8] = buffer_data_1[3535:3528];
        layer3[58][23:16] = buffer_data_1[3543:3536];
        layer3[58][31:24] = buffer_data_1[3551:3544];
        layer3[58][39:32] = buffer_data_1[3559:3552];
        layer4[58][7:0] = buffer_data_0[3527:3520];
        layer4[58][15:8] = buffer_data_0[3535:3528];
        layer4[58][23:16] = buffer_data_0[3543:3536];
        layer4[58][31:24] = buffer_data_0[3551:3544];
        layer4[58][39:32] = buffer_data_0[3559:3552];
        layer0[59][7:0] = buffer_data_4[3535:3528];
        layer0[59][15:8] = buffer_data_4[3543:3536];
        layer0[59][23:16] = buffer_data_4[3551:3544];
        layer0[59][31:24] = buffer_data_4[3559:3552];
        layer0[59][39:32] = buffer_data_4[3567:3560];
        layer1[59][7:0] = buffer_data_3[3535:3528];
        layer1[59][15:8] = buffer_data_3[3543:3536];
        layer1[59][23:16] = buffer_data_3[3551:3544];
        layer1[59][31:24] = buffer_data_3[3559:3552];
        layer1[59][39:32] = buffer_data_3[3567:3560];
        layer2[59][7:0] = buffer_data_2[3535:3528];
        layer2[59][15:8] = buffer_data_2[3543:3536];
        layer2[59][23:16] = buffer_data_2[3551:3544];
        layer2[59][31:24] = buffer_data_2[3559:3552];
        layer2[59][39:32] = buffer_data_2[3567:3560];
        layer3[59][7:0] = buffer_data_1[3535:3528];
        layer3[59][15:8] = buffer_data_1[3543:3536];
        layer3[59][23:16] = buffer_data_1[3551:3544];
        layer3[59][31:24] = buffer_data_1[3559:3552];
        layer3[59][39:32] = buffer_data_1[3567:3560];
        layer4[59][7:0] = buffer_data_0[3535:3528];
        layer4[59][15:8] = buffer_data_0[3543:3536];
        layer4[59][23:16] = buffer_data_0[3551:3544];
        layer4[59][31:24] = buffer_data_0[3559:3552];
        layer4[59][39:32] = buffer_data_0[3567:3560];
        layer0[60][7:0] = buffer_data_4[3543:3536];
        layer0[60][15:8] = buffer_data_4[3551:3544];
        layer0[60][23:16] = buffer_data_4[3559:3552];
        layer0[60][31:24] = buffer_data_4[3567:3560];
        layer0[60][39:32] = buffer_data_4[3575:3568];
        layer1[60][7:0] = buffer_data_3[3543:3536];
        layer1[60][15:8] = buffer_data_3[3551:3544];
        layer1[60][23:16] = buffer_data_3[3559:3552];
        layer1[60][31:24] = buffer_data_3[3567:3560];
        layer1[60][39:32] = buffer_data_3[3575:3568];
        layer2[60][7:0] = buffer_data_2[3543:3536];
        layer2[60][15:8] = buffer_data_2[3551:3544];
        layer2[60][23:16] = buffer_data_2[3559:3552];
        layer2[60][31:24] = buffer_data_2[3567:3560];
        layer2[60][39:32] = buffer_data_2[3575:3568];
        layer3[60][7:0] = buffer_data_1[3543:3536];
        layer3[60][15:8] = buffer_data_1[3551:3544];
        layer3[60][23:16] = buffer_data_1[3559:3552];
        layer3[60][31:24] = buffer_data_1[3567:3560];
        layer3[60][39:32] = buffer_data_1[3575:3568];
        layer4[60][7:0] = buffer_data_0[3543:3536];
        layer4[60][15:8] = buffer_data_0[3551:3544];
        layer4[60][23:16] = buffer_data_0[3559:3552];
        layer4[60][31:24] = buffer_data_0[3567:3560];
        layer4[60][39:32] = buffer_data_0[3575:3568];
        layer0[61][7:0] = buffer_data_4[3551:3544];
        layer0[61][15:8] = buffer_data_4[3559:3552];
        layer0[61][23:16] = buffer_data_4[3567:3560];
        layer0[61][31:24] = buffer_data_4[3575:3568];
        layer0[61][39:32] = buffer_data_4[3583:3576];
        layer1[61][7:0] = buffer_data_3[3551:3544];
        layer1[61][15:8] = buffer_data_3[3559:3552];
        layer1[61][23:16] = buffer_data_3[3567:3560];
        layer1[61][31:24] = buffer_data_3[3575:3568];
        layer1[61][39:32] = buffer_data_3[3583:3576];
        layer2[61][7:0] = buffer_data_2[3551:3544];
        layer2[61][15:8] = buffer_data_2[3559:3552];
        layer2[61][23:16] = buffer_data_2[3567:3560];
        layer2[61][31:24] = buffer_data_2[3575:3568];
        layer2[61][39:32] = buffer_data_2[3583:3576];
        layer3[61][7:0] = buffer_data_1[3551:3544];
        layer3[61][15:8] = buffer_data_1[3559:3552];
        layer3[61][23:16] = buffer_data_1[3567:3560];
        layer3[61][31:24] = buffer_data_1[3575:3568];
        layer3[61][39:32] = buffer_data_1[3583:3576];
        layer4[61][7:0] = buffer_data_0[3551:3544];
        layer4[61][15:8] = buffer_data_0[3559:3552];
        layer4[61][23:16] = buffer_data_0[3567:3560];
        layer4[61][31:24] = buffer_data_0[3575:3568];
        layer4[61][39:32] = buffer_data_0[3583:3576];
        layer0[62][7:0] = buffer_data_4[3559:3552];
        layer0[62][15:8] = buffer_data_4[3567:3560];
        layer0[62][23:16] = buffer_data_4[3575:3568];
        layer0[62][31:24] = buffer_data_4[3583:3576];
        layer0[62][39:32] = buffer_data_4[3591:3584];
        layer1[62][7:0] = buffer_data_3[3559:3552];
        layer1[62][15:8] = buffer_data_3[3567:3560];
        layer1[62][23:16] = buffer_data_3[3575:3568];
        layer1[62][31:24] = buffer_data_3[3583:3576];
        layer1[62][39:32] = buffer_data_3[3591:3584];
        layer2[62][7:0] = buffer_data_2[3559:3552];
        layer2[62][15:8] = buffer_data_2[3567:3560];
        layer2[62][23:16] = buffer_data_2[3575:3568];
        layer2[62][31:24] = buffer_data_2[3583:3576];
        layer2[62][39:32] = buffer_data_2[3591:3584];
        layer3[62][7:0] = buffer_data_1[3559:3552];
        layer3[62][15:8] = buffer_data_1[3567:3560];
        layer3[62][23:16] = buffer_data_1[3575:3568];
        layer3[62][31:24] = buffer_data_1[3583:3576];
        layer3[62][39:32] = buffer_data_1[3591:3584];
        layer4[62][7:0] = buffer_data_0[3559:3552];
        layer4[62][15:8] = buffer_data_0[3567:3560];
        layer4[62][23:16] = buffer_data_0[3575:3568];
        layer4[62][31:24] = buffer_data_0[3583:3576];
        layer4[62][39:32] = buffer_data_0[3591:3584];
        layer0[63][7:0] = buffer_data_4[3567:3560];
        layer0[63][15:8] = buffer_data_4[3575:3568];
        layer0[63][23:16] = buffer_data_4[3583:3576];
        layer0[63][31:24] = buffer_data_4[3591:3584];
        layer0[63][39:32] = buffer_data_4[3599:3592];
        layer1[63][7:0] = buffer_data_3[3567:3560];
        layer1[63][15:8] = buffer_data_3[3575:3568];
        layer1[63][23:16] = buffer_data_3[3583:3576];
        layer1[63][31:24] = buffer_data_3[3591:3584];
        layer1[63][39:32] = buffer_data_3[3599:3592];
        layer2[63][7:0] = buffer_data_2[3567:3560];
        layer2[63][15:8] = buffer_data_2[3575:3568];
        layer2[63][23:16] = buffer_data_2[3583:3576];
        layer2[63][31:24] = buffer_data_2[3591:3584];
        layer2[63][39:32] = buffer_data_2[3599:3592];
        layer3[63][7:0] = buffer_data_1[3567:3560];
        layer3[63][15:8] = buffer_data_1[3575:3568];
        layer3[63][23:16] = buffer_data_1[3583:3576];
        layer3[63][31:24] = buffer_data_1[3591:3584];
        layer3[63][39:32] = buffer_data_1[3599:3592];
        layer4[63][7:0] = buffer_data_0[3567:3560];
        layer4[63][15:8] = buffer_data_0[3575:3568];
        layer4[63][23:16] = buffer_data_0[3583:3576];
        layer4[63][31:24] = buffer_data_0[3591:3584];
        layer4[63][39:32] = buffer_data_0[3599:3592];
    end
    ST_GAUSSIAN_7: begin
        layer0[0][7:0] = buffer_data_4[3575:3568];
        layer0[0][15:8] = buffer_data_4[3583:3576];
        layer0[0][23:16] = buffer_data_4[3591:3584];
        layer0[0][31:24] = buffer_data_4[3599:3592];
        layer0[0][39:32] = buffer_data_4[3607:3600];
        layer1[0][7:0] = buffer_data_3[3575:3568];
        layer1[0][15:8] = buffer_data_3[3583:3576];
        layer1[0][23:16] = buffer_data_3[3591:3584];
        layer1[0][31:24] = buffer_data_3[3599:3592];
        layer1[0][39:32] = buffer_data_3[3607:3600];
        layer2[0][7:0] = buffer_data_2[3575:3568];
        layer2[0][15:8] = buffer_data_2[3583:3576];
        layer2[0][23:16] = buffer_data_2[3591:3584];
        layer2[0][31:24] = buffer_data_2[3599:3592];
        layer2[0][39:32] = buffer_data_2[3607:3600];
        layer3[0][7:0] = buffer_data_1[3575:3568];
        layer3[0][15:8] = buffer_data_1[3583:3576];
        layer3[0][23:16] = buffer_data_1[3591:3584];
        layer3[0][31:24] = buffer_data_1[3599:3592];
        layer3[0][39:32] = buffer_data_1[3607:3600];
        layer4[0][7:0] = buffer_data_0[3575:3568];
        layer4[0][15:8] = buffer_data_0[3583:3576];
        layer4[0][23:16] = buffer_data_0[3591:3584];
        layer4[0][31:24] = buffer_data_0[3599:3592];
        layer4[0][39:32] = buffer_data_0[3607:3600];
        layer0[1][7:0] = buffer_data_4[3583:3576];
        layer0[1][15:8] = buffer_data_4[3591:3584];
        layer0[1][23:16] = buffer_data_4[3599:3592];
        layer0[1][31:24] = buffer_data_4[3607:3600];
        layer0[1][39:32] = buffer_data_4[3615:3608];
        layer1[1][7:0] = buffer_data_3[3583:3576];
        layer1[1][15:8] = buffer_data_3[3591:3584];
        layer1[1][23:16] = buffer_data_3[3599:3592];
        layer1[1][31:24] = buffer_data_3[3607:3600];
        layer1[1][39:32] = buffer_data_3[3615:3608];
        layer2[1][7:0] = buffer_data_2[3583:3576];
        layer2[1][15:8] = buffer_data_2[3591:3584];
        layer2[1][23:16] = buffer_data_2[3599:3592];
        layer2[1][31:24] = buffer_data_2[3607:3600];
        layer2[1][39:32] = buffer_data_2[3615:3608];
        layer3[1][7:0] = buffer_data_1[3583:3576];
        layer3[1][15:8] = buffer_data_1[3591:3584];
        layer3[1][23:16] = buffer_data_1[3599:3592];
        layer3[1][31:24] = buffer_data_1[3607:3600];
        layer3[1][39:32] = buffer_data_1[3615:3608];
        layer4[1][7:0] = buffer_data_0[3583:3576];
        layer4[1][15:8] = buffer_data_0[3591:3584];
        layer4[1][23:16] = buffer_data_0[3599:3592];
        layer4[1][31:24] = buffer_data_0[3607:3600];
        layer4[1][39:32] = buffer_data_0[3615:3608];
        layer0[2][7:0] = buffer_data_4[3591:3584];
        layer0[2][15:8] = buffer_data_4[3599:3592];
        layer0[2][23:16] = buffer_data_4[3607:3600];
        layer0[2][31:24] = buffer_data_4[3615:3608];
        layer0[2][39:32] = buffer_data_4[3623:3616];
        layer1[2][7:0] = buffer_data_3[3591:3584];
        layer1[2][15:8] = buffer_data_3[3599:3592];
        layer1[2][23:16] = buffer_data_3[3607:3600];
        layer1[2][31:24] = buffer_data_3[3615:3608];
        layer1[2][39:32] = buffer_data_3[3623:3616];
        layer2[2][7:0] = buffer_data_2[3591:3584];
        layer2[2][15:8] = buffer_data_2[3599:3592];
        layer2[2][23:16] = buffer_data_2[3607:3600];
        layer2[2][31:24] = buffer_data_2[3615:3608];
        layer2[2][39:32] = buffer_data_2[3623:3616];
        layer3[2][7:0] = buffer_data_1[3591:3584];
        layer3[2][15:8] = buffer_data_1[3599:3592];
        layer3[2][23:16] = buffer_data_1[3607:3600];
        layer3[2][31:24] = buffer_data_1[3615:3608];
        layer3[2][39:32] = buffer_data_1[3623:3616];
        layer4[2][7:0] = buffer_data_0[3591:3584];
        layer4[2][15:8] = buffer_data_0[3599:3592];
        layer4[2][23:16] = buffer_data_0[3607:3600];
        layer4[2][31:24] = buffer_data_0[3615:3608];
        layer4[2][39:32] = buffer_data_0[3623:3616];
        layer0[3][7:0] = buffer_data_4[3599:3592];
        layer0[3][15:8] = buffer_data_4[3607:3600];
        layer0[3][23:16] = buffer_data_4[3615:3608];
        layer0[3][31:24] = buffer_data_4[3623:3616];
        layer0[3][39:32] = buffer_data_4[3631:3624];
        layer1[3][7:0] = buffer_data_3[3599:3592];
        layer1[3][15:8] = buffer_data_3[3607:3600];
        layer1[3][23:16] = buffer_data_3[3615:3608];
        layer1[3][31:24] = buffer_data_3[3623:3616];
        layer1[3][39:32] = buffer_data_3[3631:3624];
        layer2[3][7:0] = buffer_data_2[3599:3592];
        layer2[3][15:8] = buffer_data_2[3607:3600];
        layer2[3][23:16] = buffer_data_2[3615:3608];
        layer2[3][31:24] = buffer_data_2[3623:3616];
        layer2[3][39:32] = buffer_data_2[3631:3624];
        layer3[3][7:0] = buffer_data_1[3599:3592];
        layer3[3][15:8] = buffer_data_1[3607:3600];
        layer3[3][23:16] = buffer_data_1[3615:3608];
        layer3[3][31:24] = buffer_data_1[3623:3616];
        layer3[3][39:32] = buffer_data_1[3631:3624];
        layer4[3][7:0] = buffer_data_0[3599:3592];
        layer4[3][15:8] = buffer_data_0[3607:3600];
        layer4[3][23:16] = buffer_data_0[3615:3608];
        layer4[3][31:24] = buffer_data_0[3623:3616];
        layer4[3][39:32] = buffer_data_0[3631:3624];
        layer0[4][7:0] = buffer_data_4[3607:3600];
        layer0[4][15:8] = buffer_data_4[3615:3608];
        layer0[4][23:16] = buffer_data_4[3623:3616];
        layer0[4][31:24] = buffer_data_4[3631:3624];
        layer0[4][39:32] = buffer_data_4[3639:3632];
        layer1[4][7:0] = buffer_data_3[3607:3600];
        layer1[4][15:8] = buffer_data_3[3615:3608];
        layer1[4][23:16] = buffer_data_3[3623:3616];
        layer1[4][31:24] = buffer_data_3[3631:3624];
        layer1[4][39:32] = buffer_data_3[3639:3632];
        layer2[4][7:0] = buffer_data_2[3607:3600];
        layer2[4][15:8] = buffer_data_2[3615:3608];
        layer2[4][23:16] = buffer_data_2[3623:3616];
        layer2[4][31:24] = buffer_data_2[3631:3624];
        layer2[4][39:32] = buffer_data_2[3639:3632];
        layer3[4][7:0] = buffer_data_1[3607:3600];
        layer3[4][15:8] = buffer_data_1[3615:3608];
        layer3[4][23:16] = buffer_data_1[3623:3616];
        layer3[4][31:24] = buffer_data_1[3631:3624];
        layer3[4][39:32] = buffer_data_1[3639:3632];
        layer4[4][7:0] = buffer_data_0[3607:3600];
        layer4[4][15:8] = buffer_data_0[3615:3608];
        layer4[4][23:16] = buffer_data_0[3623:3616];
        layer4[4][31:24] = buffer_data_0[3631:3624];
        layer4[4][39:32] = buffer_data_0[3639:3632];
        layer0[5][7:0] = buffer_data_4[3615:3608];
        layer0[5][15:8] = buffer_data_4[3623:3616];
        layer0[5][23:16] = buffer_data_4[3631:3624];
        layer0[5][31:24] = buffer_data_4[3639:3632];
        layer0[5][39:32] = buffer_data_4[3647:3640];
        layer1[5][7:0] = buffer_data_3[3615:3608];
        layer1[5][15:8] = buffer_data_3[3623:3616];
        layer1[5][23:16] = buffer_data_3[3631:3624];
        layer1[5][31:24] = buffer_data_3[3639:3632];
        layer1[5][39:32] = buffer_data_3[3647:3640];
        layer2[5][7:0] = buffer_data_2[3615:3608];
        layer2[5][15:8] = buffer_data_2[3623:3616];
        layer2[5][23:16] = buffer_data_2[3631:3624];
        layer2[5][31:24] = buffer_data_2[3639:3632];
        layer2[5][39:32] = buffer_data_2[3647:3640];
        layer3[5][7:0] = buffer_data_1[3615:3608];
        layer3[5][15:8] = buffer_data_1[3623:3616];
        layer3[5][23:16] = buffer_data_1[3631:3624];
        layer3[5][31:24] = buffer_data_1[3639:3632];
        layer3[5][39:32] = buffer_data_1[3647:3640];
        layer4[5][7:0] = buffer_data_0[3615:3608];
        layer4[5][15:8] = buffer_data_0[3623:3616];
        layer4[5][23:16] = buffer_data_0[3631:3624];
        layer4[5][31:24] = buffer_data_0[3639:3632];
        layer4[5][39:32] = buffer_data_0[3647:3640];
        layer0[6][7:0] = buffer_data_4[3623:3616];
        layer0[6][15:8] = buffer_data_4[3631:3624];
        layer0[6][23:16] = buffer_data_4[3639:3632];
        layer0[6][31:24] = buffer_data_4[3647:3640];
        layer0[6][39:32] = buffer_data_4[3655:3648];
        layer1[6][7:0] = buffer_data_3[3623:3616];
        layer1[6][15:8] = buffer_data_3[3631:3624];
        layer1[6][23:16] = buffer_data_3[3639:3632];
        layer1[6][31:24] = buffer_data_3[3647:3640];
        layer1[6][39:32] = buffer_data_3[3655:3648];
        layer2[6][7:0] = buffer_data_2[3623:3616];
        layer2[6][15:8] = buffer_data_2[3631:3624];
        layer2[6][23:16] = buffer_data_2[3639:3632];
        layer2[6][31:24] = buffer_data_2[3647:3640];
        layer2[6][39:32] = buffer_data_2[3655:3648];
        layer3[6][7:0] = buffer_data_1[3623:3616];
        layer3[6][15:8] = buffer_data_1[3631:3624];
        layer3[6][23:16] = buffer_data_1[3639:3632];
        layer3[6][31:24] = buffer_data_1[3647:3640];
        layer3[6][39:32] = buffer_data_1[3655:3648];
        layer4[6][7:0] = buffer_data_0[3623:3616];
        layer4[6][15:8] = buffer_data_0[3631:3624];
        layer4[6][23:16] = buffer_data_0[3639:3632];
        layer4[6][31:24] = buffer_data_0[3647:3640];
        layer4[6][39:32] = buffer_data_0[3655:3648];
        layer0[7][7:0] = buffer_data_4[3631:3624];
        layer0[7][15:8] = buffer_data_4[3639:3632];
        layer0[7][23:16] = buffer_data_4[3647:3640];
        layer0[7][31:24] = buffer_data_4[3655:3648];
        layer0[7][39:32] = buffer_data_4[3663:3656];
        layer1[7][7:0] = buffer_data_3[3631:3624];
        layer1[7][15:8] = buffer_data_3[3639:3632];
        layer1[7][23:16] = buffer_data_3[3647:3640];
        layer1[7][31:24] = buffer_data_3[3655:3648];
        layer1[7][39:32] = buffer_data_3[3663:3656];
        layer2[7][7:0] = buffer_data_2[3631:3624];
        layer2[7][15:8] = buffer_data_2[3639:3632];
        layer2[7][23:16] = buffer_data_2[3647:3640];
        layer2[7][31:24] = buffer_data_2[3655:3648];
        layer2[7][39:32] = buffer_data_2[3663:3656];
        layer3[7][7:0] = buffer_data_1[3631:3624];
        layer3[7][15:8] = buffer_data_1[3639:3632];
        layer3[7][23:16] = buffer_data_1[3647:3640];
        layer3[7][31:24] = buffer_data_1[3655:3648];
        layer3[7][39:32] = buffer_data_1[3663:3656];
        layer4[7][7:0] = buffer_data_0[3631:3624];
        layer4[7][15:8] = buffer_data_0[3639:3632];
        layer4[7][23:16] = buffer_data_0[3647:3640];
        layer4[7][31:24] = buffer_data_0[3655:3648];
        layer4[7][39:32] = buffer_data_0[3663:3656];
        layer0[8][7:0] = buffer_data_4[3639:3632];
        layer0[8][15:8] = buffer_data_4[3647:3640];
        layer0[8][23:16] = buffer_data_4[3655:3648];
        layer0[8][31:24] = buffer_data_4[3663:3656];
        layer0[8][39:32] = buffer_data_4[3671:3664];
        layer1[8][7:0] = buffer_data_3[3639:3632];
        layer1[8][15:8] = buffer_data_3[3647:3640];
        layer1[8][23:16] = buffer_data_3[3655:3648];
        layer1[8][31:24] = buffer_data_3[3663:3656];
        layer1[8][39:32] = buffer_data_3[3671:3664];
        layer2[8][7:0] = buffer_data_2[3639:3632];
        layer2[8][15:8] = buffer_data_2[3647:3640];
        layer2[8][23:16] = buffer_data_2[3655:3648];
        layer2[8][31:24] = buffer_data_2[3663:3656];
        layer2[8][39:32] = buffer_data_2[3671:3664];
        layer3[8][7:0] = buffer_data_1[3639:3632];
        layer3[8][15:8] = buffer_data_1[3647:3640];
        layer3[8][23:16] = buffer_data_1[3655:3648];
        layer3[8][31:24] = buffer_data_1[3663:3656];
        layer3[8][39:32] = buffer_data_1[3671:3664];
        layer4[8][7:0] = buffer_data_0[3639:3632];
        layer4[8][15:8] = buffer_data_0[3647:3640];
        layer4[8][23:16] = buffer_data_0[3655:3648];
        layer4[8][31:24] = buffer_data_0[3663:3656];
        layer4[8][39:32] = buffer_data_0[3671:3664];
        layer0[9][7:0] = buffer_data_4[3647:3640];
        layer0[9][15:8] = buffer_data_4[3655:3648];
        layer0[9][23:16] = buffer_data_4[3663:3656];
        layer0[9][31:24] = buffer_data_4[3671:3664];
        layer0[9][39:32] = buffer_data_4[3679:3672];
        layer1[9][7:0] = buffer_data_3[3647:3640];
        layer1[9][15:8] = buffer_data_3[3655:3648];
        layer1[9][23:16] = buffer_data_3[3663:3656];
        layer1[9][31:24] = buffer_data_3[3671:3664];
        layer1[9][39:32] = buffer_data_3[3679:3672];
        layer2[9][7:0] = buffer_data_2[3647:3640];
        layer2[9][15:8] = buffer_data_2[3655:3648];
        layer2[9][23:16] = buffer_data_2[3663:3656];
        layer2[9][31:24] = buffer_data_2[3671:3664];
        layer2[9][39:32] = buffer_data_2[3679:3672];
        layer3[9][7:0] = buffer_data_1[3647:3640];
        layer3[9][15:8] = buffer_data_1[3655:3648];
        layer3[9][23:16] = buffer_data_1[3663:3656];
        layer3[9][31:24] = buffer_data_1[3671:3664];
        layer3[9][39:32] = buffer_data_1[3679:3672];
        layer4[9][7:0] = buffer_data_0[3647:3640];
        layer4[9][15:8] = buffer_data_0[3655:3648];
        layer4[9][23:16] = buffer_data_0[3663:3656];
        layer4[9][31:24] = buffer_data_0[3671:3664];
        layer4[9][39:32] = buffer_data_0[3679:3672];
        layer0[10][7:0] = buffer_data_4[3655:3648];
        layer0[10][15:8] = buffer_data_4[3663:3656];
        layer0[10][23:16] = buffer_data_4[3671:3664];
        layer0[10][31:24] = buffer_data_4[3679:3672];
        layer0[10][39:32] = buffer_data_4[3687:3680];
        layer1[10][7:0] = buffer_data_3[3655:3648];
        layer1[10][15:8] = buffer_data_3[3663:3656];
        layer1[10][23:16] = buffer_data_3[3671:3664];
        layer1[10][31:24] = buffer_data_3[3679:3672];
        layer1[10][39:32] = buffer_data_3[3687:3680];
        layer2[10][7:0] = buffer_data_2[3655:3648];
        layer2[10][15:8] = buffer_data_2[3663:3656];
        layer2[10][23:16] = buffer_data_2[3671:3664];
        layer2[10][31:24] = buffer_data_2[3679:3672];
        layer2[10][39:32] = buffer_data_2[3687:3680];
        layer3[10][7:0] = buffer_data_1[3655:3648];
        layer3[10][15:8] = buffer_data_1[3663:3656];
        layer3[10][23:16] = buffer_data_1[3671:3664];
        layer3[10][31:24] = buffer_data_1[3679:3672];
        layer3[10][39:32] = buffer_data_1[3687:3680];
        layer4[10][7:0] = buffer_data_0[3655:3648];
        layer4[10][15:8] = buffer_data_0[3663:3656];
        layer4[10][23:16] = buffer_data_0[3671:3664];
        layer4[10][31:24] = buffer_data_0[3679:3672];
        layer4[10][39:32] = buffer_data_0[3687:3680];
        layer0[11][7:0] = buffer_data_4[3663:3656];
        layer0[11][15:8] = buffer_data_4[3671:3664];
        layer0[11][23:16] = buffer_data_4[3679:3672];
        layer0[11][31:24] = buffer_data_4[3687:3680];
        layer0[11][39:32] = buffer_data_4[3695:3688];
        layer1[11][7:0] = buffer_data_3[3663:3656];
        layer1[11][15:8] = buffer_data_3[3671:3664];
        layer1[11][23:16] = buffer_data_3[3679:3672];
        layer1[11][31:24] = buffer_data_3[3687:3680];
        layer1[11][39:32] = buffer_data_3[3695:3688];
        layer2[11][7:0] = buffer_data_2[3663:3656];
        layer2[11][15:8] = buffer_data_2[3671:3664];
        layer2[11][23:16] = buffer_data_2[3679:3672];
        layer2[11][31:24] = buffer_data_2[3687:3680];
        layer2[11][39:32] = buffer_data_2[3695:3688];
        layer3[11][7:0] = buffer_data_1[3663:3656];
        layer3[11][15:8] = buffer_data_1[3671:3664];
        layer3[11][23:16] = buffer_data_1[3679:3672];
        layer3[11][31:24] = buffer_data_1[3687:3680];
        layer3[11][39:32] = buffer_data_1[3695:3688];
        layer4[11][7:0] = buffer_data_0[3663:3656];
        layer4[11][15:8] = buffer_data_0[3671:3664];
        layer4[11][23:16] = buffer_data_0[3679:3672];
        layer4[11][31:24] = buffer_data_0[3687:3680];
        layer4[11][39:32] = buffer_data_0[3695:3688];
        layer0[12][7:0] = buffer_data_4[3671:3664];
        layer0[12][15:8] = buffer_data_4[3679:3672];
        layer0[12][23:16] = buffer_data_4[3687:3680];
        layer0[12][31:24] = buffer_data_4[3695:3688];
        layer0[12][39:32] = buffer_data_4[3703:3696];
        layer1[12][7:0] = buffer_data_3[3671:3664];
        layer1[12][15:8] = buffer_data_3[3679:3672];
        layer1[12][23:16] = buffer_data_3[3687:3680];
        layer1[12][31:24] = buffer_data_3[3695:3688];
        layer1[12][39:32] = buffer_data_3[3703:3696];
        layer2[12][7:0] = buffer_data_2[3671:3664];
        layer2[12][15:8] = buffer_data_2[3679:3672];
        layer2[12][23:16] = buffer_data_2[3687:3680];
        layer2[12][31:24] = buffer_data_2[3695:3688];
        layer2[12][39:32] = buffer_data_2[3703:3696];
        layer3[12][7:0] = buffer_data_1[3671:3664];
        layer3[12][15:8] = buffer_data_1[3679:3672];
        layer3[12][23:16] = buffer_data_1[3687:3680];
        layer3[12][31:24] = buffer_data_1[3695:3688];
        layer3[12][39:32] = buffer_data_1[3703:3696];
        layer4[12][7:0] = buffer_data_0[3671:3664];
        layer4[12][15:8] = buffer_data_0[3679:3672];
        layer4[12][23:16] = buffer_data_0[3687:3680];
        layer4[12][31:24] = buffer_data_0[3695:3688];
        layer4[12][39:32] = buffer_data_0[3703:3696];
        layer0[13][7:0] = buffer_data_4[3679:3672];
        layer0[13][15:8] = buffer_data_4[3687:3680];
        layer0[13][23:16] = buffer_data_4[3695:3688];
        layer0[13][31:24] = buffer_data_4[3703:3696];
        layer0[13][39:32] = buffer_data_4[3711:3704];
        layer1[13][7:0] = buffer_data_3[3679:3672];
        layer1[13][15:8] = buffer_data_3[3687:3680];
        layer1[13][23:16] = buffer_data_3[3695:3688];
        layer1[13][31:24] = buffer_data_3[3703:3696];
        layer1[13][39:32] = buffer_data_3[3711:3704];
        layer2[13][7:0] = buffer_data_2[3679:3672];
        layer2[13][15:8] = buffer_data_2[3687:3680];
        layer2[13][23:16] = buffer_data_2[3695:3688];
        layer2[13][31:24] = buffer_data_2[3703:3696];
        layer2[13][39:32] = buffer_data_2[3711:3704];
        layer3[13][7:0] = buffer_data_1[3679:3672];
        layer3[13][15:8] = buffer_data_1[3687:3680];
        layer3[13][23:16] = buffer_data_1[3695:3688];
        layer3[13][31:24] = buffer_data_1[3703:3696];
        layer3[13][39:32] = buffer_data_1[3711:3704];
        layer4[13][7:0] = buffer_data_0[3679:3672];
        layer4[13][15:8] = buffer_data_0[3687:3680];
        layer4[13][23:16] = buffer_data_0[3695:3688];
        layer4[13][31:24] = buffer_data_0[3703:3696];
        layer4[13][39:32] = buffer_data_0[3711:3704];
        layer0[14][7:0] = buffer_data_4[3687:3680];
        layer0[14][15:8] = buffer_data_4[3695:3688];
        layer0[14][23:16] = buffer_data_4[3703:3696];
        layer0[14][31:24] = buffer_data_4[3711:3704];
        layer0[14][39:32] = buffer_data_4[3719:3712];
        layer1[14][7:0] = buffer_data_3[3687:3680];
        layer1[14][15:8] = buffer_data_3[3695:3688];
        layer1[14][23:16] = buffer_data_3[3703:3696];
        layer1[14][31:24] = buffer_data_3[3711:3704];
        layer1[14][39:32] = buffer_data_3[3719:3712];
        layer2[14][7:0] = buffer_data_2[3687:3680];
        layer2[14][15:8] = buffer_data_2[3695:3688];
        layer2[14][23:16] = buffer_data_2[3703:3696];
        layer2[14][31:24] = buffer_data_2[3711:3704];
        layer2[14][39:32] = buffer_data_2[3719:3712];
        layer3[14][7:0] = buffer_data_1[3687:3680];
        layer3[14][15:8] = buffer_data_1[3695:3688];
        layer3[14][23:16] = buffer_data_1[3703:3696];
        layer3[14][31:24] = buffer_data_1[3711:3704];
        layer3[14][39:32] = buffer_data_1[3719:3712];
        layer4[14][7:0] = buffer_data_0[3687:3680];
        layer4[14][15:8] = buffer_data_0[3695:3688];
        layer4[14][23:16] = buffer_data_0[3703:3696];
        layer4[14][31:24] = buffer_data_0[3711:3704];
        layer4[14][39:32] = buffer_data_0[3719:3712];
        layer0[15][7:0] = buffer_data_4[3695:3688];
        layer0[15][15:8] = buffer_data_4[3703:3696];
        layer0[15][23:16] = buffer_data_4[3711:3704];
        layer0[15][31:24] = buffer_data_4[3719:3712];
        layer0[15][39:32] = buffer_data_4[3727:3720];
        layer1[15][7:0] = buffer_data_3[3695:3688];
        layer1[15][15:8] = buffer_data_3[3703:3696];
        layer1[15][23:16] = buffer_data_3[3711:3704];
        layer1[15][31:24] = buffer_data_3[3719:3712];
        layer1[15][39:32] = buffer_data_3[3727:3720];
        layer2[15][7:0] = buffer_data_2[3695:3688];
        layer2[15][15:8] = buffer_data_2[3703:3696];
        layer2[15][23:16] = buffer_data_2[3711:3704];
        layer2[15][31:24] = buffer_data_2[3719:3712];
        layer2[15][39:32] = buffer_data_2[3727:3720];
        layer3[15][7:0] = buffer_data_1[3695:3688];
        layer3[15][15:8] = buffer_data_1[3703:3696];
        layer3[15][23:16] = buffer_data_1[3711:3704];
        layer3[15][31:24] = buffer_data_1[3719:3712];
        layer3[15][39:32] = buffer_data_1[3727:3720];
        layer4[15][7:0] = buffer_data_0[3695:3688];
        layer4[15][15:8] = buffer_data_0[3703:3696];
        layer4[15][23:16] = buffer_data_0[3711:3704];
        layer4[15][31:24] = buffer_data_0[3719:3712];
        layer4[15][39:32] = buffer_data_0[3727:3720];
        layer0[16][7:0] = buffer_data_4[3703:3696];
        layer0[16][15:8] = buffer_data_4[3711:3704];
        layer0[16][23:16] = buffer_data_4[3719:3712];
        layer0[16][31:24] = buffer_data_4[3727:3720];
        layer0[16][39:32] = buffer_data_4[3735:3728];
        layer1[16][7:0] = buffer_data_3[3703:3696];
        layer1[16][15:8] = buffer_data_3[3711:3704];
        layer1[16][23:16] = buffer_data_3[3719:3712];
        layer1[16][31:24] = buffer_data_3[3727:3720];
        layer1[16][39:32] = buffer_data_3[3735:3728];
        layer2[16][7:0] = buffer_data_2[3703:3696];
        layer2[16][15:8] = buffer_data_2[3711:3704];
        layer2[16][23:16] = buffer_data_2[3719:3712];
        layer2[16][31:24] = buffer_data_2[3727:3720];
        layer2[16][39:32] = buffer_data_2[3735:3728];
        layer3[16][7:0] = buffer_data_1[3703:3696];
        layer3[16][15:8] = buffer_data_1[3711:3704];
        layer3[16][23:16] = buffer_data_1[3719:3712];
        layer3[16][31:24] = buffer_data_1[3727:3720];
        layer3[16][39:32] = buffer_data_1[3735:3728];
        layer4[16][7:0] = buffer_data_0[3703:3696];
        layer4[16][15:8] = buffer_data_0[3711:3704];
        layer4[16][23:16] = buffer_data_0[3719:3712];
        layer4[16][31:24] = buffer_data_0[3727:3720];
        layer4[16][39:32] = buffer_data_0[3735:3728];
        layer0[17][7:0] = buffer_data_4[3711:3704];
        layer0[17][15:8] = buffer_data_4[3719:3712];
        layer0[17][23:16] = buffer_data_4[3727:3720];
        layer0[17][31:24] = buffer_data_4[3735:3728];
        layer0[17][39:32] = buffer_data_4[3743:3736];
        layer1[17][7:0] = buffer_data_3[3711:3704];
        layer1[17][15:8] = buffer_data_3[3719:3712];
        layer1[17][23:16] = buffer_data_3[3727:3720];
        layer1[17][31:24] = buffer_data_3[3735:3728];
        layer1[17][39:32] = buffer_data_3[3743:3736];
        layer2[17][7:0] = buffer_data_2[3711:3704];
        layer2[17][15:8] = buffer_data_2[3719:3712];
        layer2[17][23:16] = buffer_data_2[3727:3720];
        layer2[17][31:24] = buffer_data_2[3735:3728];
        layer2[17][39:32] = buffer_data_2[3743:3736];
        layer3[17][7:0] = buffer_data_1[3711:3704];
        layer3[17][15:8] = buffer_data_1[3719:3712];
        layer3[17][23:16] = buffer_data_1[3727:3720];
        layer3[17][31:24] = buffer_data_1[3735:3728];
        layer3[17][39:32] = buffer_data_1[3743:3736];
        layer4[17][7:0] = buffer_data_0[3711:3704];
        layer4[17][15:8] = buffer_data_0[3719:3712];
        layer4[17][23:16] = buffer_data_0[3727:3720];
        layer4[17][31:24] = buffer_data_0[3735:3728];
        layer4[17][39:32] = buffer_data_0[3743:3736];
        layer0[18][7:0] = buffer_data_4[3719:3712];
        layer0[18][15:8] = buffer_data_4[3727:3720];
        layer0[18][23:16] = buffer_data_4[3735:3728];
        layer0[18][31:24] = buffer_data_4[3743:3736];
        layer0[18][39:32] = buffer_data_4[3751:3744];
        layer1[18][7:0] = buffer_data_3[3719:3712];
        layer1[18][15:8] = buffer_data_3[3727:3720];
        layer1[18][23:16] = buffer_data_3[3735:3728];
        layer1[18][31:24] = buffer_data_3[3743:3736];
        layer1[18][39:32] = buffer_data_3[3751:3744];
        layer2[18][7:0] = buffer_data_2[3719:3712];
        layer2[18][15:8] = buffer_data_2[3727:3720];
        layer2[18][23:16] = buffer_data_2[3735:3728];
        layer2[18][31:24] = buffer_data_2[3743:3736];
        layer2[18][39:32] = buffer_data_2[3751:3744];
        layer3[18][7:0] = buffer_data_1[3719:3712];
        layer3[18][15:8] = buffer_data_1[3727:3720];
        layer3[18][23:16] = buffer_data_1[3735:3728];
        layer3[18][31:24] = buffer_data_1[3743:3736];
        layer3[18][39:32] = buffer_data_1[3751:3744];
        layer4[18][7:0] = buffer_data_0[3719:3712];
        layer4[18][15:8] = buffer_data_0[3727:3720];
        layer4[18][23:16] = buffer_data_0[3735:3728];
        layer4[18][31:24] = buffer_data_0[3743:3736];
        layer4[18][39:32] = buffer_data_0[3751:3744];
        layer0[19][7:0] = buffer_data_4[3727:3720];
        layer0[19][15:8] = buffer_data_4[3735:3728];
        layer0[19][23:16] = buffer_data_4[3743:3736];
        layer0[19][31:24] = buffer_data_4[3751:3744];
        layer0[19][39:32] = buffer_data_4[3759:3752];
        layer1[19][7:0] = buffer_data_3[3727:3720];
        layer1[19][15:8] = buffer_data_3[3735:3728];
        layer1[19][23:16] = buffer_data_3[3743:3736];
        layer1[19][31:24] = buffer_data_3[3751:3744];
        layer1[19][39:32] = buffer_data_3[3759:3752];
        layer2[19][7:0] = buffer_data_2[3727:3720];
        layer2[19][15:8] = buffer_data_2[3735:3728];
        layer2[19][23:16] = buffer_data_2[3743:3736];
        layer2[19][31:24] = buffer_data_2[3751:3744];
        layer2[19][39:32] = buffer_data_2[3759:3752];
        layer3[19][7:0] = buffer_data_1[3727:3720];
        layer3[19][15:8] = buffer_data_1[3735:3728];
        layer3[19][23:16] = buffer_data_1[3743:3736];
        layer3[19][31:24] = buffer_data_1[3751:3744];
        layer3[19][39:32] = buffer_data_1[3759:3752];
        layer4[19][7:0] = buffer_data_0[3727:3720];
        layer4[19][15:8] = buffer_data_0[3735:3728];
        layer4[19][23:16] = buffer_data_0[3743:3736];
        layer4[19][31:24] = buffer_data_0[3751:3744];
        layer4[19][39:32] = buffer_data_0[3759:3752];
        layer0[20][7:0] = buffer_data_4[3735:3728];
        layer0[20][15:8] = buffer_data_4[3743:3736];
        layer0[20][23:16] = buffer_data_4[3751:3744];
        layer0[20][31:24] = buffer_data_4[3759:3752];
        layer0[20][39:32] = buffer_data_4[3767:3760];
        layer1[20][7:0] = buffer_data_3[3735:3728];
        layer1[20][15:8] = buffer_data_3[3743:3736];
        layer1[20][23:16] = buffer_data_3[3751:3744];
        layer1[20][31:24] = buffer_data_3[3759:3752];
        layer1[20][39:32] = buffer_data_3[3767:3760];
        layer2[20][7:0] = buffer_data_2[3735:3728];
        layer2[20][15:8] = buffer_data_2[3743:3736];
        layer2[20][23:16] = buffer_data_2[3751:3744];
        layer2[20][31:24] = buffer_data_2[3759:3752];
        layer2[20][39:32] = buffer_data_2[3767:3760];
        layer3[20][7:0] = buffer_data_1[3735:3728];
        layer3[20][15:8] = buffer_data_1[3743:3736];
        layer3[20][23:16] = buffer_data_1[3751:3744];
        layer3[20][31:24] = buffer_data_1[3759:3752];
        layer3[20][39:32] = buffer_data_1[3767:3760];
        layer4[20][7:0] = buffer_data_0[3735:3728];
        layer4[20][15:8] = buffer_data_0[3743:3736];
        layer4[20][23:16] = buffer_data_0[3751:3744];
        layer4[20][31:24] = buffer_data_0[3759:3752];
        layer4[20][39:32] = buffer_data_0[3767:3760];
        layer0[21][7:0] = buffer_data_4[3743:3736];
        layer0[21][15:8] = buffer_data_4[3751:3744];
        layer0[21][23:16] = buffer_data_4[3759:3752];
        layer0[21][31:24] = buffer_data_4[3767:3760];
        layer0[21][39:32] = buffer_data_4[3775:3768];
        layer1[21][7:0] = buffer_data_3[3743:3736];
        layer1[21][15:8] = buffer_data_3[3751:3744];
        layer1[21][23:16] = buffer_data_3[3759:3752];
        layer1[21][31:24] = buffer_data_3[3767:3760];
        layer1[21][39:32] = buffer_data_3[3775:3768];
        layer2[21][7:0] = buffer_data_2[3743:3736];
        layer2[21][15:8] = buffer_data_2[3751:3744];
        layer2[21][23:16] = buffer_data_2[3759:3752];
        layer2[21][31:24] = buffer_data_2[3767:3760];
        layer2[21][39:32] = buffer_data_2[3775:3768];
        layer3[21][7:0] = buffer_data_1[3743:3736];
        layer3[21][15:8] = buffer_data_1[3751:3744];
        layer3[21][23:16] = buffer_data_1[3759:3752];
        layer3[21][31:24] = buffer_data_1[3767:3760];
        layer3[21][39:32] = buffer_data_1[3775:3768];
        layer4[21][7:0] = buffer_data_0[3743:3736];
        layer4[21][15:8] = buffer_data_0[3751:3744];
        layer4[21][23:16] = buffer_data_0[3759:3752];
        layer4[21][31:24] = buffer_data_0[3767:3760];
        layer4[21][39:32] = buffer_data_0[3775:3768];
        layer0[22][7:0] = buffer_data_4[3751:3744];
        layer0[22][15:8] = buffer_data_4[3759:3752];
        layer0[22][23:16] = buffer_data_4[3767:3760];
        layer0[22][31:24] = buffer_data_4[3775:3768];
        layer0[22][39:32] = buffer_data_4[3783:3776];
        layer1[22][7:0] = buffer_data_3[3751:3744];
        layer1[22][15:8] = buffer_data_3[3759:3752];
        layer1[22][23:16] = buffer_data_3[3767:3760];
        layer1[22][31:24] = buffer_data_3[3775:3768];
        layer1[22][39:32] = buffer_data_3[3783:3776];
        layer2[22][7:0] = buffer_data_2[3751:3744];
        layer2[22][15:8] = buffer_data_2[3759:3752];
        layer2[22][23:16] = buffer_data_2[3767:3760];
        layer2[22][31:24] = buffer_data_2[3775:3768];
        layer2[22][39:32] = buffer_data_2[3783:3776];
        layer3[22][7:0] = buffer_data_1[3751:3744];
        layer3[22][15:8] = buffer_data_1[3759:3752];
        layer3[22][23:16] = buffer_data_1[3767:3760];
        layer3[22][31:24] = buffer_data_1[3775:3768];
        layer3[22][39:32] = buffer_data_1[3783:3776];
        layer4[22][7:0] = buffer_data_0[3751:3744];
        layer4[22][15:8] = buffer_data_0[3759:3752];
        layer4[22][23:16] = buffer_data_0[3767:3760];
        layer4[22][31:24] = buffer_data_0[3775:3768];
        layer4[22][39:32] = buffer_data_0[3783:3776];
        layer0[23][7:0] = buffer_data_4[3759:3752];
        layer0[23][15:8] = buffer_data_4[3767:3760];
        layer0[23][23:16] = buffer_data_4[3775:3768];
        layer0[23][31:24] = buffer_data_4[3783:3776];
        layer0[23][39:32] = buffer_data_4[3791:3784];
        layer1[23][7:0] = buffer_data_3[3759:3752];
        layer1[23][15:8] = buffer_data_3[3767:3760];
        layer1[23][23:16] = buffer_data_3[3775:3768];
        layer1[23][31:24] = buffer_data_3[3783:3776];
        layer1[23][39:32] = buffer_data_3[3791:3784];
        layer2[23][7:0] = buffer_data_2[3759:3752];
        layer2[23][15:8] = buffer_data_2[3767:3760];
        layer2[23][23:16] = buffer_data_2[3775:3768];
        layer2[23][31:24] = buffer_data_2[3783:3776];
        layer2[23][39:32] = buffer_data_2[3791:3784];
        layer3[23][7:0] = buffer_data_1[3759:3752];
        layer3[23][15:8] = buffer_data_1[3767:3760];
        layer3[23][23:16] = buffer_data_1[3775:3768];
        layer3[23][31:24] = buffer_data_1[3783:3776];
        layer3[23][39:32] = buffer_data_1[3791:3784];
        layer4[23][7:0] = buffer_data_0[3759:3752];
        layer4[23][15:8] = buffer_data_0[3767:3760];
        layer4[23][23:16] = buffer_data_0[3775:3768];
        layer4[23][31:24] = buffer_data_0[3783:3776];
        layer4[23][39:32] = buffer_data_0[3791:3784];
        layer0[24][7:0] = buffer_data_4[3767:3760];
        layer0[24][15:8] = buffer_data_4[3775:3768];
        layer0[24][23:16] = buffer_data_4[3783:3776];
        layer0[24][31:24] = buffer_data_4[3791:3784];
        layer0[24][39:32] = buffer_data_4[3799:3792];
        layer1[24][7:0] = buffer_data_3[3767:3760];
        layer1[24][15:8] = buffer_data_3[3775:3768];
        layer1[24][23:16] = buffer_data_3[3783:3776];
        layer1[24][31:24] = buffer_data_3[3791:3784];
        layer1[24][39:32] = buffer_data_3[3799:3792];
        layer2[24][7:0] = buffer_data_2[3767:3760];
        layer2[24][15:8] = buffer_data_2[3775:3768];
        layer2[24][23:16] = buffer_data_2[3783:3776];
        layer2[24][31:24] = buffer_data_2[3791:3784];
        layer2[24][39:32] = buffer_data_2[3799:3792];
        layer3[24][7:0] = buffer_data_1[3767:3760];
        layer3[24][15:8] = buffer_data_1[3775:3768];
        layer3[24][23:16] = buffer_data_1[3783:3776];
        layer3[24][31:24] = buffer_data_1[3791:3784];
        layer3[24][39:32] = buffer_data_1[3799:3792];
        layer4[24][7:0] = buffer_data_0[3767:3760];
        layer4[24][15:8] = buffer_data_0[3775:3768];
        layer4[24][23:16] = buffer_data_0[3783:3776];
        layer4[24][31:24] = buffer_data_0[3791:3784];
        layer4[24][39:32] = buffer_data_0[3799:3792];
        layer0[25][7:0] = buffer_data_4[3775:3768];
        layer0[25][15:8] = buffer_data_4[3783:3776];
        layer0[25][23:16] = buffer_data_4[3791:3784];
        layer0[25][31:24] = buffer_data_4[3799:3792];
        layer0[25][39:32] = buffer_data_4[3807:3800];
        layer1[25][7:0] = buffer_data_3[3775:3768];
        layer1[25][15:8] = buffer_data_3[3783:3776];
        layer1[25][23:16] = buffer_data_3[3791:3784];
        layer1[25][31:24] = buffer_data_3[3799:3792];
        layer1[25][39:32] = buffer_data_3[3807:3800];
        layer2[25][7:0] = buffer_data_2[3775:3768];
        layer2[25][15:8] = buffer_data_2[3783:3776];
        layer2[25][23:16] = buffer_data_2[3791:3784];
        layer2[25][31:24] = buffer_data_2[3799:3792];
        layer2[25][39:32] = buffer_data_2[3807:3800];
        layer3[25][7:0] = buffer_data_1[3775:3768];
        layer3[25][15:8] = buffer_data_1[3783:3776];
        layer3[25][23:16] = buffer_data_1[3791:3784];
        layer3[25][31:24] = buffer_data_1[3799:3792];
        layer3[25][39:32] = buffer_data_1[3807:3800];
        layer4[25][7:0] = buffer_data_0[3775:3768];
        layer4[25][15:8] = buffer_data_0[3783:3776];
        layer4[25][23:16] = buffer_data_0[3791:3784];
        layer4[25][31:24] = buffer_data_0[3799:3792];
        layer4[25][39:32] = buffer_data_0[3807:3800];
        layer0[26][7:0] = buffer_data_4[3783:3776];
        layer0[26][15:8] = buffer_data_4[3791:3784];
        layer0[26][23:16] = buffer_data_4[3799:3792];
        layer0[26][31:24] = buffer_data_4[3807:3800];
        layer0[26][39:32] = buffer_data_4[3815:3808];
        layer1[26][7:0] = buffer_data_3[3783:3776];
        layer1[26][15:8] = buffer_data_3[3791:3784];
        layer1[26][23:16] = buffer_data_3[3799:3792];
        layer1[26][31:24] = buffer_data_3[3807:3800];
        layer1[26][39:32] = buffer_data_3[3815:3808];
        layer2[26][7:0] = buffer_data_2[3783:3776];
        layer2[26][15:8] = buffer_data_2[3791:3784];
        layer2[26][23:16] = buffer_data_2[3799:3792];
        layer2[26][31:24] = buffer_data_2[3807:3800];
        layer2[26][39:32] = buffer_data_2[3815:3808];
        layer3[26][7:0] = buffer_data_1[3783:3776];
        layer3[26][15:8] = buffer_data_1[3791:3784];
        layer3[26][23:16] = buffer_data_1[3799:3792];
        layer3[26][31:24] = buffer_data_1[3807:3800];
        layer3[26][39:32] = buffer_data_1[3815:3808];
        layer4[26][7:0] = buffer_data_0[3783:3776];
        layer4[26][15:8] = buffer_data_0[3791:3784];
        layer4[26][23:16] = buffer_data_0[3799:3792];
        layer4[26][31:24] = buffer_data_0[3807:3800];
        layer4[26][39:32] = buffer_data_0[3815:3808];
        layer0[27][7:0] = buffer_data_4[3791:3784];
        layer0[27][15:8] = buffer_data_4[3799:3792];
        layer0[27][23:16] = buffer_data_4[3807:3800];
        layer0[27][31:24] = buffer_data_4[3815:3808];
        layer0[27][39:32] = buffer_data_4[3823:3816];
        layer1[27][7:0] = buffer_data_3[3791:3784];
        layer1[27][15:8] = buffer_data_3[3799:3792];
        layer1[27][23:16] = buffer_data_3[3807:3800];
        layer1[27][31:24] = buffer_data_3[3815:3808];
        layer1[27][39:32] = buffer_data_3[3823:3816];
        layer2[27][7:0] = buffer_data_2[3791:3784];
        layer2[27][15:8] = buffer_data_2[3799:3792];
        layer2[27][23:16] = buffer_data_2[3807:3800];
        layer2[27][31:24] = buffer_data_2[3815:3808];
        layer2[27][39:32] = buffer_data_2[3823:3816];
        layer3[27][7:0] = buffer_data_1[3791:3784];
        layer3[27][15:8] = buffer_data_1[3799:3792];
        layer3[27][23:16] = buffer_data_1[3807:3800];
        layer3[27][31:24] = buffer_data_1[3815:3808];
        layer3[27][39:32] = buffer_data_1[3823:3816];
        layer4[27][7:0] = buffer_data_0[3791:3784];
        layer4[27][15:8] = buffer_data_0[3799:3792];
        layer4[27][23:16] = buffer_data_0[3807:3800];
        layer4[27][31:24] = buffer_data_0[3815:3808];
        layer4[27][39:32] = buffer_data_0[3823:3816];
        layer0[28][7:0] = buffer_data_4[3799:3792];
        layer0[28][15:8] = buffer_data_4[3807:3800];
        layer0[28][23:16] = buffer_data_4[3815:3808];
        layer0[28][31:24] = buffer_data_4[3823:3816];
        layer0[28][39:32] = buffer_data_4[3831:3824];
        layer1[28][7:0] = buffer_data_3[3799:3792];
        layer1[28][15:8] = buffer_data_3[3807:3800];
        layer1[28][23:16] = buffer_data_3[3815:3808];
        layer1[28][31:24] = buffer_data_3[3823:3816];
        layer1[28][39:32] = buffer_data_3[3831:3824];
        layer2[28][7:0] = buffer_data_2[3799:3792];
        layer2[28][15:8] = buffer_data_2[3807:3800];
        layer2[28][23:16] = buffer_data_2[3815:3808];
        layer2[28][31:24] = buffer_data_2[3823:3816];
        layer2[28][39:32] = buffer_data_2[3831:3824];
        layer3[28][7:0] = buffer_data_1[3799:3792];
        layer3[28][15:8] = buffer_data_1[3807:3800];
        layer3[28][23:16] = buffer_data_1[3815:3808];
        layer3[28][31:24] = buffer_data_1[3823:3816];
        layer3[28][39:32] = buffer_data_1[3831:3824];
        layer4[28][7:0] = buffer_data_0[3799:3792];
        layer4[28][15:8] = buffer_data_0[3807:3800];
        layer4[28][23:16] = buffer_data_0[3815:3808];
        layer4[28][31:24] = buffer_data_0[3823:3816];
        layer4[28][39:32] = buffer_data_0[3831:3824];
        layer0[29][7:0] = buffer_data_4[3807:3800];
        layer0[29][15:8] = buffer_data_4[3815:3808];
        layer0[29][23:16] = buffer_data_4[3823:3816];
        layer0[29][31:24] = buffer_data_4[3831:3824];
        layer0[29][39:32] = buffer_data_4[3839:3832];
        layer1[29][7:0] = buffer_data_3[3807:3800];
        layer1[29][15:8] = buffer_data_3[3815:3808];
        layer1[29][23:16] = buffer_data_3[3823:3816];
        layer1[29][31:24] = buffer_data_3[3831:3824];
        layer1[29][39:32] = buffer_data_3[3839:3832];
        layer2[29][7:0] = buffer_data_2[3807:3800];
        layer2[29][15:8] = buffer_data_2[3815:3808];
        layer2[29][23:16] = buffer_data_2[3823:3816];
        layer2[29][31:24] = buffer_data_2[3831:3824];
        layer2[29][39:32] = buffer_data_2[3839:3832];
        layer3[29][7:0] = buffer_data_1[3807:3800];
        layer3[29][15:8] = buffer_data_1[3815:3808];
        layer3[29][23:16] = buffer_data_1[3823:3816];
        layer3[29][31:24] = buffer_data_1[3831:3824];
        layer3[29][39:32] = buffer_data_1[3839:3832];
        layer4[29][7:0] = buffer_data_0[3807:3800];
        layer4[29][15:8] = buffer_data_0[3815:3808];
        layer4[29][23:16] = buffer_data_0[3823:3816];
        layer4[29][31:24] = buffer_data_0[3831:3824];
        layer4[29][39:32] = buffer_data_0[3839:3832];
        layer0[30][7:0] = buffer_data_4[3815:3808];
        layer0[30][15:8] = buffer_data_4[3823:3816];
        layer0[30][23:16] = buffer_data_4[3831:3824];
        layer0[30][31:24] = buffer_data_4[3839:3832];
        layer0[30][39:32] = buffer_data_4[3847:3840];
        layer1[30][7:0] = buffer_data_3[3815:3808];
        layer1[30][15:8] = buffer_data_3[3823:3816];
        layer1[30][23:16] = buffer_data_3[3831:3824];
        layer1[30][31:24] = buffer_data_3[3839:3832];
        layer1[30][39:32] = buffer_data_3[3847:3840];
        layer2[30][7:0] = buffer_data_2[3815:3808];
        layer2[30][15:8] = buffer_data_2[3823:3816];
        layer2[30][23:16] = buffer_data_2[3831:3824];
        layer2[30][31:24] = buffer_data_2[3839:3832];
        layer2[30][39:32] = buffer_data_2[3847:3840];
        layer3[30][7:0] = buffer_data_1[3815:3808];
        layer3[30][15:8] = buffer_data_1[3823:3816];
        layer3[30][23:16] = buffer_data_1[3831:3824];
        layer3[30][31:24] = buffer_data_1[3839:3832];
        layer3[30][39:32] = buffer_data_1[3847:3840];
        layer4[30][7:0] = buffer_data_0[3815:3808];
        layer4[30][15:8] = buffer_data_0[3823:3816];
        layer4[30][23:16] = buffer_data_0[3831:3824];
        layer4[30][31:24] = buffer_data_0[3839:3832];
        layer4[30][39:32] = buffer_data_0[3847:3840];
        layer0[31][7:0] = buffer_data_4[3823:3816];
        layer0[31][15:8] = buffer_data_4[3831:3824];
        layer0[31][23:16] = buffer_data_4[3839:3832];
        layer0[31][31:24] = buffer_data_4[3847:3840];
        layer0[31][39:32] = buffer_data_4[3855:3848];
        layer1[31][7:0] = buffer_data_3[3823:3816];
        layer1[31][15:8] = buffer_data_3[3831:3824];
        layer1[31][23:16] = buffer_data_3[3839:3832];
        layer1[31][31:24] = buffer_data_3[3847:3840];
        layer1[31][39:32] = buffer_data_3[3855:3848];
        layer2[31][7:0] = buffer_data_2[3823:3816];
        layer2[31][15:8] = buffer_data_2[3831:3824];
        layer2[31][23:16] = buffer_data_2[3839:3832];
        layer2[31][31:24] = buffer_data_2[3847:3840];
        layer2[31][39:32] = buffer_data_2[3855:3848];
        layer3[31][7:0] = buffer_data_1[3823:3816];
        layer3[31][15:8] = buffer_data_1[3831:3824];
        layer3[31][23:16] = buffer_data_1[3839:3832];
        layer3[31][31:24] = buffer_data_1[3847:3840];
        layer3[31][39:32] = buffer_data_1[3855:3848];
        layer4[31][7:0] = buffer_data_0[3823:3816];
        layer4[31][15:8] = buffer_data_0[3831:3824];
        layer4[31][23:16] = buffer_data_0[3839:3832];
        layer4[31][31:24] = buffer_data_0[3847:3840];
        layer4[31][39:32] = buffer_data_0[3855:3848];
        layer0[32][7:0] = buffer_data_4[3831:3824];
        layer0[32][15:8] = buffer_data_4[3839:3832];
        layer0[32][23:16] = buffer_data_4[3847:3840];
        layer0[32][31:24] = buffer_data_4[3855:3848];
        layer0[32][39:32] = buffer_data_4[3863:3856];
        layer1[32][7:0] = buffer_data_3[3831:3824];
        layer1[32][15:8] = buffer_data_3[3839:3832];
        layer1[32][23:16] = buffer_data_3[3847:3840];
        layer1[32][31:24] = buffer_data_3[3855:3848];
        layer1[32][39:32] = buffer_data_3[3863:3856];
        layer2[32][7:0] = buffer_data_2[3831:3824];
        layer2[32][15:8] = buffer_data_2[3839:3832];
        layer2[32][23:16] = buffer_data_2[3847:3840];
        layer2[32][31:24] = buffer_data_2[3855:3848];
        layer2[32][39:32] = buffer_data_2[3863:3856];
        layer3[32][7:0] = buffer_data_1[3831:3824];
        layer3[32][15:8] = buffer_data_1[3839:3832];
        layer3[32][23:16] = buffer_data_1[3847:3840];
        layer3[32][31:24] = buffer_data_1[3855:3848];
        layer3[32][39:32] = buffer_data_1[3863:3856];
        layer4[32][7:0] = buffer_data_0[3831:3824];
        layer4[32][15:8] = buffer_data_0[3839:3832];
        layer4[32][23:16] = buffer_data_0[3847:3840];
        layer4[32][31:24] = buffer_data_0[3855:3848];
        layer4[32][39:32] = buffer_data_0[3863:3856];
        layer0[33][7:0] = buffer_data_4[3839:3832];
        layer0[33][15:8] = buffer_data_4[3847:3840];
        layer0[33][23:16] = buffer_data_4[3855:3848];
        layer0[33][31:24] = buffer_data_4[3863:3856];
        layer0[33][39:32] = buffer_data_4[3871:3864];
        layer1[33][7:0] = buffer_data_3[3839:3832];
        layer1[33][15:8] = buffer_data_3[3847:3840];
        layer1[33][23:16] = buffer_data_3[3855:3848];
        layer1[33][31:24] = buffer_data_3[3863:3856];
        layer1[33][39:32] = buffer_data_3[3871:3864];
        layer2[33][7:0] = buffer_data_2[3839:3832];
        layer2[33][15:8] = buffer_data_2[3847:3840];
        layer2[33][23:16] = buffer_data_2[3855:3848];
        layer2[33][31:24] = buffer_data_2[3863:3856];
        layer2[33][39:32] = buffer_data_2[3871:3864];
        layer3[33][7:0] = buffer_data_1[3839:3832];
        layer3[33][15:8] = buffer_data_1[3847:3840];
        layer3[33][23:16] = buffer_data_1[3855:3848];
        layer3[33][31:24] = buffer_data_1[3863:3856];
        layer3[33][39:32] = buffer_data_1[3871:3864];
        layer4[33][7:0] = buffer_data_0[3839:3832];
        layer4[33][15:8] = buffer_data_0[3847:3840];
        layer4[33][23:16] = buffer_data_0[3855:3848];
        layer4[33][31:24] = buffer_data_0[3863:3856];
        layer4[33][39:32] = buffer_data_0[3871:3864];
        layer0[34][7:0] = buffer_data_4[3847:3840];
        layer0[34][15:8] = buffer_data_4[3855:3848];
        layer0[34][23:16] = buffer_data_4[3863:3856];
        layer0[34][31:24] = buffer_data_4[3871:3864];
        layer0[34][39:32] = buffer_data_4[3879:3872];
        layer1[34][7:0] = buffer_data_3[3847:3840];
        layer1[34][15:8] = buffer_data_3[3855:3848];
        layer1[34][23:16] = buffer_data_3[3863:3856];
        layer1[34][31:24] = buffer_data_3[3871:3864];
        layer1[34][39:32] = buffer_data_3[3879:3872];
        layer2[34][7:0] = buffer_data_2[3847:3840];
        layer2[34][15:8] = buffer_data_2[3855:3848];
        layer2[34][23:16] = buffer_data_2[3863:3856];
        layer2[34][31:24] = buffer_data_2[3871:3864];
        layer2[34][39:32] = buffer_data_2[3879:3872];
        layer3[34][7:0] = buffer_data_1[3847:3840];
        layer3[34][15:8] = buffer_data_1[3855:3848];
        layer3[34][23:16] = buffer_data_1[3863:3856];
        layer3[34][31:24] = buffer_data_1[3871:3864];
        layer3[34][39:32] = buffer_data_1[3879:3872];
        layer4[34][7:0] = buffer_data_0[3847:3840];
        layer4[34][15:8] = buffer_data_0[3855:3848];
        layer4[34][23:16] = buffer_data_0[3863:3856];
        layer4[34][31:24] = buffer_data_0[3871:3864];
        layer4[34][39:32] = buffer_data_0[3879:3872];
        layer0[35][7:0] = buffer_data_4[3855:3848];
        layer0[35][15:8] = buffer_data_4[3863:3856];
        layer0[35][23:16] = buffer_data_4[3871:3864];
        layer0[35][31:24] = buffer_data_4[3879:3872];
        layer0[35][39:32] = buffer_data_4[3887:3880];
        layer1[35][7:0] = buffer_data_3[3855:3848];
        layer1[35][15:8] = buffer_data_3[3863:3856];
        layer1[35][23:16] = buffer_data_3[3871:3864];
        layer1[35][31:24] = buffer_data_3[3879:3872];
        layer1[35][39:32] = buffer_data_3[3887:3880];
        layer2[35][7:0] = buffer_data_2[3855:3848];
        layer2[35][15:8] = buffer_data_2[3863:3856];
        layer2[35][23:16] = buffer_data_2[3871:3864];
        layer2[35][31:24] = buffer_data_2[3879:3872];
        layer2[35][39:32] = buffer_data_2[3887:3880];
        layer3[35][7:0] = buffer_data_1[3855:3848];
        layer3[35][15:8] = buffer_data_1[3863:3856];
        layer3[35][23:16] = buffer_data_1[3871:3864];
        layer3[35][31:24] = buffer_data_1[3879:3872];
        layer3[35][39:32] = buffer_data_1[3887:3880];
        layer4[35][7:0] = buffer_data_0[3855:3848];
        layer4[35][15:8] = buffer_data_0[3863:3856];
        layer4[35][23:16] = buffer_data_0[3871:3864];
        layer4[35][31:24] = buffer_data_0[3879:3872];
        layer4[35][39:32] = buffer_data_0[3887:3880];
        layer0[36][7:0] = buffer_data_4[3863:3856];
        layer0[36][15:8] = buffer_data_4[3871:3864];
        layer0[36][23:16] = buffer_data_4[3879:3872];
        layer0[36][31:24] = buffer_data_4[3887:3880];
        layer0[36][39:32] = buffer_data_4[3895:3888];
        layer1[36][7:0] = buffer_data_3[3863:3856];
        layer1[36][15:8] = buffer_data_3[3871:3864];
        layer1[36][23:16] = buffer_data_3[3879:3872];
        layer1[36][31:24] = buffer_data_3[3887:3880];
        layer1[36][39:32] = buffer_data_3[3895:3888];
        layer2[36][7:0] = buffer_data_2[3863:3856];
        layer2[36][15:8] = buffer_data_2[3871:3864];
        layer2[36][23:16] = buffer_data_2[3879:3872];
        layer2[36][31:24] = buffer_data_2[3887:3880];
        layer2[36][39:32] = buffer_data_2[3895:3888];
        layer3[36][7:0] = buffer_data_1[3863:3856];
        layer3[36][15:8] = buffer_data_1[3871:3864];
        layer3[36][23:16] = buffer_data_1[3879:3872];
        layer3[36][31:24] = buffer_data_1[3887:3880];
        layer3[36][39:32] = buffer_data_1[3895:3888];
        layer4[36][7:0] = buffer_data_0[3863:3856];
        layer4[36][15:8] = buffer_data_0[3871:3864];
        layer4[36][23:16] = buffer_data_0[3879:3872];
        layer4[36][31:24] = buffer_data_0[3887:3880];
        layer4[36][39:32] = buffer_data_0[3895:3888];
        layer0[37][7:0] = buffer_data_4[3871:3864];
        layer0[37][15:8] = buffer_data_4[3879:3872];
        layer0[37][23:16] = buffer_data_4[3887:3880];
        layer0[37][31:24] = buffer_data_4[3895:3888];
        layer0[37][39:32] = buffer_data_4[3903:3896];
        layer1[37][7:0] = buffer_data_3[3871:3864];
        layer1[37][15:8] = buffer_data_3[3879:3872];
        layer1[37][23:16] = buffer_data_3[3887:3880];
        layer1[37][31:24] = buffer_data_3[3895:3888];
        layer1[37][39:32] = buffer_data_3[3903:3896];
        layer2[37][7:0] = buffer_data_2[3871:3864];
        layer2[37][15:8] = buffer_data_2[3879:3872];
        layer2[37][23:16] = buffer_data_2[3887:3880];
        layer2[37][31:24] = buffer_data_2[3895:3888];
        layer2[37][39:32] = buffer_data_2[3903:3896];
        layer3[37][7:0] = buffer_data_1[3871:3864];
        layer3[37][15:8] = buffer_data_1[3879:3872];
        layer3[37][23:16] = buffer_data_1[3887:3880];
        layer3[37][31:24] = buffer_data_1[3895:3888];
        layer3[37][39:32] = buffer_data_1[3903:3896];
        layer4[37][7:0] = buffer_data_0[3871:3864];
        layer4[37][15:8] = buffer_data_0[3879:3872];
        layer4[37][23:16] = buffer_data_0[3887:3880];
        layer4[37][31:24] = buffer_data_0[3895:3888];
        layer4[37][39:32] = buffer_data_0[3903:3896];
        layer0[38][7:0] = buffer_data_4[3879:3872];
        layer0[38][15:8] = buffer_data_4[3887:3880];
        layer0[38][23:16] = buffer_data_4[3895:3888];
        layer0[38][31:24] = buffer_data_4[3903:3896];
        layer0[38][39:32] = buffer_data_4[3911:3904];
        layer1[38][7:0] = buffer_data_3[3879:3872];
        layer1[38][15:8] = buffer_data_3[3887:3880];
        layer1[38][23:16] = buffer_data_3[3895:3888];
        layer1[38][31:24] = buffer_data_3[3903:3896];
        layer1[38][39:32] = buffer_data_3[3911:3904];
        layer2[38][7:0] = buffer_data_2[3879:3872];
        layer2[38][15:8] = buffer_data_2[3887:3880];
        layer2[38][23:16] = buffer_data_2[3895:3888];
        layer2[38][31:24] = buffer_data_2[3903:3896];
        layer2[38][39:32] = buffer_data_2[3911:3904];
        layer3[38][7:0] = buffer_data_1[3879:3872];
        layer3[38][15:8] = buffer_data_1[3887:3880];
        layer3[38][23:16] = buffer_data_1[3895:3888];
        layer3[38][31:24] = buffer_data_1[3903:3896];
        layer3[38][39:32] = buffer_data_1[3911:3904];
        layer4[38][7:0] = buffer_data_0[3879:3872];
        layer4[38][15:8] = buffer_data_0[3887:3880];
        layer4[38][23:16] = buffer_data_0[3895:3888];
        layer4[38][31:24] = buffer_data_0[3903:3896];
        layer4[38][39:32] = buffer_data_0[3911:3904];
        layer0[39][7:0] = buffer_data_4[3887:3880];
        layer0[39][15:8] = buffer_data_4[3895:3888];
        layer0[39][23:16] = buffer_data_4[3903:3896];
        layer0[39][31:24] = buffer_data_4[3911:3904];
        layer0[39][39:32] = buffer_data_4[3919:3912];
        layer1[39][7:0] = buffer_data_3[3887:3880];
        layer1[39][15:8] = buffer_data_3[3895:3888];
        layer1[39][23:16] = buffer_data_3[3903:3896];
        layer1[39][31:24] = buffer_data_3[3911:3904];
        layer1[39][39:32] = buffer_data_3[3919:3912];
        layer2[39][7:0] = buffer_data_2[3887:3880];
        layer2[39][15:8] = buffer_data_2[3895:3888];
        layer2[39][23:16] = buffer_data_2[3903:3896];
        layer2[39][31:24] = buffer_data_2[3911:3904];
        layer2[39][39:32] = buffer_data_2[3919:3912];
        layer3[39][7:0] = buffer_data_1[3887:3880];
        layer3[39][15:8] = buffer_data_1[3895:3888];
        layer3[39][23:16] = buffer_data_1[3903:3896];
        layer3[39][31:24] = buffer_data_1[3911:3904];
        layer3[39][39:32] = buffer_data_1[3919:3912];
        layer4[39][7:0] = buffer_data_0[3887:3880];
        layer4[39][15:8] = buffer_data_0[3895:3888];
        layer4[39][23:16] = buffer_data_0[3903:3896];
        layer4[39][31:24] = buffer_data_0[3911:3904];
        layer4[39][39:32] = buffer_data_0[3919:3912];
        layer0[40][7:0] = buffer_data_4[3895:3888];
        layer0[40][15:8] = buffer_data_4[3903:3896];
        layer0[40][23:16] = buffer_data_4[3911:3904];
        layer0[40][31:24] = buffer_data_4[3919:3912];
        layer0[40][39:32] = buffer_data_4[3927:3920];
        layer1[40][7:0] = buffer_data_3[3895:3888];
        layer1[40][15:8] = buffer_data_3[3903:3896];
        layer1[40][23:16] = buffer_data_3[3911:3904];
        layer1[40][31:24] = buffer_data_3[3919:3912];
        layer1[40][39:32] = buffer_data_3[3927:3920];
        layer2[40][7:0] = buffer_data_2[3895:3888];
        layer2[40][15:8] = buffer_data_2[3903:3896];
        layer2[40][23:16] = buffer_data_2[3911:3904];
        layer2[40][31:24] = buffer_data_2[3919:3912];
        layer2[40][39:32] = buffer_data_2[3927:3920];
        layer3[40][7:0] = buffer_data_1[3895:3888];
        layer3[40][15:8] = buffer_data_1[3903:3896];
        layer3[40][23:16] = buffer_data_1[3911:3904];
        layer3[40][31:24] = buffer_data_1[3919:3912];
        layer3[40][39:32] = buffer_data_1[3927:3920];
        layer4[40][7:0] = buffer_data_0[3895:3888];
        layer4[40][15:8] = buffer_data_0[3903:3896];
        layer4[40][23:16] = buffer_data_0[3911:3904];
        layer4[40][31:24] = buffer_data_0[3919:3912];
        layer4[40][39:32] = buffer_data_0[3927:3920];
        layer0[41][7:0] = buffer_data_4[3903:3896];
        layer0[41][15:8] = buffer_data_4[3911:3904];
        layer0[41][23:16] = buffer_data_4[3919:3912];
        layer0[41][31:24] = buffer_data_4[3927:3920];
        layer0[41][39:32] = buffer_data_4[3935:3928];
        layer1[41][7:0] = buffer_data_3[3903:3896];
        layer1[41][15:8] = buffer_data_3[3911:3904];
        layer1[41][23:16] = buffer_data_3[3919:3912];
        layer1[41][31:24] = buffer_data_3[3927:3920];
        layer1[41][39:32] = buffer_data_3[3935:3928];
        layer2[41][7:0] = buffer_data_2[3903:3896];
        layer2[41][15:8] = buffer_data_2[3911:3904];
        layer2[41][23:16] = buffer_data_2[3919:3912];
        layer2[41][31:24] = buffer_data_2[3927:3920];
        layer2[41][39:32] = buffer_data_2[3935:3928];
        layer3[41][7:0] = buffer_data_1[3903:3896];
        layer3[41][15:8] = buffer_data_1[3911:3904];
        layer3[41][23:16] = buffer_data_1[3919:3912];
        layer3[41][31:24] = buffer_data_1[3927:3920];
        layer3[41][39:32] = buffer_data_1[3935:3928];
        layer4[41][7:0] = buffer_data_0[3903:3896];
        layer4[41][15:8] = buffer_data_0[3911:3904];
        layer4[41][23:16] = buffer_data_0[3919:3912];
        layer4[41][31:24] = buffer_data_0[3927:3920];
        layer4[41][39:32] = buffer_data_0[3935:3928];
        layer0[42][7:0] = buffer_data_4[3911:3904];
        layer0[42][15:8] = buffer_data_4[3919:3912];
        layer0[42][23:16] = buffer_data_4[3927:3920];
        layer0[42][31:24] = buffer_data_4[3935:3928];
        layer0[42][39:32] = buffer_data_4[3943:3936];
        layer1[42][7:0] = buffer_data_3[3911:3904];
        layer1[42][15:8] = buffer_data_3[3919:3912];
        layer1[42][23:16] = buffer_data_3[3927:3920];
        layer1[42][31:24] = buffer_data_3[3935:3928];
        layer1[42][39:32] = buffer_data_3[3943:3936];
        layer2[42][7:0] = buffer_data_2[3911:3904];
        layer2[42][15:8] = buffer_data_2[3919:3912];
        layer2[42][23:16] = buffer_data_2[3927:3920];
        layer2[42][31:24] = buffer_data_2[3935:3928];
        layer2[42][39:32] = buffer_data_2[3943:3936];
        layer3[42][7:0] = buffer_data_1[3911:3904];
        layer3[42][15:8] = buffer_data_1[3919:3912];
        layer3[42][23:16] = buffer_data_1[3927:3920];
        layer3[42][31:24] = buffer_data_1[3935:3928];
        layer3[42][39:32] = buffer_data_1[3943:3936];
        layer4[42][7:0] = buffer_data_0[3911:3904];
        layer4[42][15:8] = buffer_data_0[3919:3912];
        layer4[42][23:16] = buffer_data_0[3927:3920];
        layer4[42][31:24] = buffer_data_0[3935:3928];
        layer4[42][39:32] = buffer_data_0[3943:3936];
        layer0[43][7:0] = buffer_data_4[3919:3912];
        layer0[43][15:8] = buffer_data_4[3927:3920];
        layer0[43][23:16] = buffer_data_4[3935:3928];
        layer0[43][31:24] = buffer_data_4[3943:3936];
        layer0[43][39:32] = buffer_data_4[3951:3944];
        layer1[43][7:0] = buffer_data_3[3919:3912];
        layer1[43][15:8] = buffer_data_3[3927:3920];
        layer1[43][23:16] = buffer_data_3[3935:3928];
        layer1[43][31:24] = buffer_data_3[3943:3936];
        layer1[43][39:32] = buffer_data_3[3951:3944];
        layer2[43][7:0] = buffer_data_2[3919:3912];
        layer2[43][15:8] = buffer_data_2[3927:3920];
        layer2[43][23:16] = buffer_data_2[3935:3928];
        layer2[43][31:24] = buffer_data_2[3943:3936];
        layer2[43][39:32] = buffer_data_2[3951:3944];
        layer3[43][7:0] = buffer_data_1[3919:3912];
        layer3[43][15:8] = buffer_data_1[3927:3920];
        layer3[43][23:16] = buffer_data_1[3935:3928];
        layer3[43][31:24] = buffer_data_1[3943:3936];
        layer3[43][39:32] = buffer_data_1[3951:3944];
        layer4[43][7:0] = buffer_data_0[3919:3912];
        layer4[43][15:8] = buffer_data_0[3927:3920];
        layer4[43][23:16] = buffer_data_0[3935:3928];
        layer4[43][31:24] = buffer_data_0[3943:3936];
        layer4[43][39:32] = buffer_data_0[3951:3944];
        layer0[44][7:0] = buffer_data_4[3927:3920];
        layer0[44][15:8] = buffer_data_4[3935:3928];
        layer0[44][23:16] = buffer_data_4[3943:3936];
        layer0[44][31:24] = buffer_data_4[3951:3944];
        layer0[44][39:32] = buffer_data_4[3959:3952];
        layer1[44][7:0] = buffer_data_3[3927:3920];
        layer1[44][15:8] = buffer_data_3[3935:3928];
        layer1[44][23:16] = buffer_data_3[3943:3936];
        layer1[44][31:24] = buffer_data_3[3951:3944];
        layer1[44][39:32] = buffer_data_3[3959:3952];
        layer2[44][7:0] = buffer_data_2[3927:3920];
        layer2[44][15:8] = buffer_data_2[3935:3928];
        layer2[44][23:16] = buffer_data_2[3943:3936];
        layer2[44][31:24] = buffer_data_2[3951:3944];
        layer2[44][39:32] = buffer_data_2[3959:3952];
        layer3[44][7:0] = buffer_data_1[3927:3920];
        layer3[44][15:8] = buffer_data_1[3935:3928];
        layer3[44][23:16] = buffer_data_1[3943:3936];
        layer3[44][31:24] = buffer_data_1[3951:3944];
        layer3[44][39:32] = buffer_data_1[3959:3952];
        layer4[44][7:0] = buffer_data_0[3927:3920];
        layer4[44][15:8] = buffer_data_0[3935:3928];
        layer4[44][23:16] = buffer_data_0[3943:3936];
        layer4[44][31:24] = buffer_data_0[3951:3944];
        layer4[44][39:32] = buffer_data_0[3959:3952];
        layer0[45][7:0] = buffer_data_4[3935:3928];
        layer0[45][15:8] = buffer_data_4[3943:3936];
        layer0[45][23:16] = buffer_data_4[3951:3944];
        layer0[45][31:24] = buffer_data_4[3959:3952];
        layer0[45][39:32] = buffer_data_4[3967:3960];
        layer1[45][7:0] = buffer_data_3[3935:3928];
        layer1[45][15:8] = buffer_data_3[3943:3936];
        layer1[45][23:16] = buffer_data_3[3951:3944];
        layer1[45][31:24] = buffer_data_3[3959:3952];
        layer1[45][39:32] = buffer_data_3[3967:3960];
        layer2[45][7:0] = buffer_data_2[3935:3928];
        layer2[45][15:8] = buffer_data_2[3943:3936];
        layer2[45][23:16] = buffer_data_2[3951:3944];
        layer2[45][31:24] = buffer_data_2[3959:3952];
        layer2[45][39:32] = buffer_data_2[3967:3960];
        layer3[45][7:0] = buffer_data_1[3935:3928];
        layer3[45][15:8] = buffer_data_1[3943:3936];
        layer3[45][23:16] = buffer_data_1[3951:3944];
        layer3[45][31:24] = buffer_data_1[3959:3952];
        layer3[45][39:32] = buffer_data_1[3967:3960];
        layer4[45][7:0] = buffer_data_0[3935:3928];
        layer4[45][15:8] = buffer_data_0[3943:3936];
        layer4[45][23:16] = buffer_data_0[3951:3944];
        layer4[45][31:24] = buffer_data_0[3959:3952];
        layer4[45][39:32] = buffer_data_0[3967:3960];
        layer0[46][7:0] = buffer_data_4[3943:3936];
        layer0[46][15:8] = buffer_data_4[3951:3944];
        layer0[46][23:16] = buffer_data_4[3959:3952];
        layer0[46][31:24] = buffer_data_4[3967:3960];
        layer0[46][39:32] = buffer_data_4[3975:3968];
        layer1[46][7:0] = buffer_data_3[3943:3936];
        layer1[46][15:8] = buffer_data_3[3951:3944];
        layer1[46][23:16] = buffer_data_3[3959:3952];
        layer1[46][31:24] = buffer_data_3[3967:3960];
        layer1[46][39:32] = buffer_data_3[3975:3968];
        layer2[46][7:0] = buffer_data_2[3943:3936];
        layer2[46][15:8] = buffer_data_2[3951:3944];
        layer2[46][23:16] = buffer_data_2[3959:3952];
        layer2[46][31:24] = buffer_data_2[3967:3960];
        layer2[46][39:32] = buffer_data_2[3975:3968];
        layer3[46][7:0] = buffer_data_1[3943:3936];
        layer3[46][15:8] = buffer_data_1[3951:3944];
        layer3[46][23:16] = buffer_data_1[3959:3952];
        layer3[46][31:24] = buffer_data_1[3967:3960];
        layer3[46][39:32] = buffer_data_1[3975:3968];
        layer4[46][7:0] = buffer_data_0[3943:3936];
        layer4[46][15:8] = buffer_data_0[3951:3944];
        layer4[46][23:16] = buffer_data_0[3959:3952];
        layer4[46][31:24] = buffer_data_0[3967:3960];
        layer4[46][39:32] = buffer_data_0[3975:3968];
        layer0[47][7:0] = buffer_data_4[3951:3944];
        layer0[47][15:8] = buffer_data_4[3959:3952];
        layer0[47][23:16] = buffer_data_4[3967:3960];
        layer0[47][31:24] = buffer_data_4[3975:3968];
        layer0[47][39:32] = buffer_data_4[3983:3976];
        layer1[47][7:0] = buffer_data_3[3951:3944];
        layer1[47][15:8] = buffer_data_3[3959:3952];
        layer1[47][23:16] = buffer_data_3[3967:3960];
        layer1[47][31:24] = buffer_data_3[3975:3968];
        layer1[47][39:32] = buffer_data_3[3983:3976];
        layer2[47][7:0] = buffer_data_2[3951:3944];
        layer2[47][15:8] = buffer_data_2[3959:3952];
        layer2[47][23:16] = buffer_data_2[3967:3960];
        layer2[47][31:24] = buffer_data_2[3975:3968];
        layer2[47][39:32] = buffer_data_2[3983:3976];
        layer3[47][7:0] = buffer_data_1[3951:3944];
        layer3[47][15:8] = buffer_data_1[3959:3952];
        layer3[47][23:16] = buffer_data_1[3967:3960];
        layer3[47][31:24] = buffer_data_1[3975:3968];
        layer3[47][39:32] = buffer_data_1[3983:3976];
        layer4[47][7:0] = buffer_data_0[3951:3944];
        layer4[47][15:8] = buffer_data_0[3959:3952];
        layer4[47][23:16] = buffer_data_0[3967:3960];
        layer4[47][31:24] = buffer_data_0[3975:3968];
        layer4[47][39:32] = buffer_data_0[3983:3976];
        layer0[48][7:0] = buffer_data_4[3959:3952];
        layer0[48][15:8] = buffer_data_4[3967:3960];
        layer0[48][23:16] = buffer_data_4[3975:3968];
        layer0[48][31:24] = buffer_data_4[3983:3976];
        layer0[48][39:32] = buffer_data_4[3991:3984];
        layer1[48][7:0] = buffer_data_3[3959:3952];
        layer1[48][15:8] = buffer_data_3[3967:3960];
        layer1[48][23:16] = buffer_data_3[3975:3968];
        layer1[48][31:24] = buffer_data_3[3983:3976];
        layer1[48][39:32] = buffer_data_3[3991:3984];
        layer2[48][7:0] = buffer_data_2[3959:3952];
        layer2[48][15:8] = buffer_data_2[3967:3960];
        layer2[48][23:16] = buffer_data_2[3975:3968];
        layer2[48][31:24] = buffer_data_2[3983:3976];
        layer2[48][39:32] = buffer_data_2[3991:3984];
        layer3[48][7:0] = buffer_data_1[3959:3952];
        layer3[48][15:8] = buffer_data_1[3967:3960];
        layer3[48][23:16] = buffer_data_1[3975:3968];
        layer3[48][31:24] = buffer_data_1[3983:3976];
        layer3[48][39:32] = buffer_data_1[3991:3984];
        layer4[48][7:0] = buffer_data_0[3959:3952];
        layer4[48][15:8] = buffer_data_0[3967:3960];
        layer4[48][23:16] = buffer_data_0[3975:3968];
        layer4[48][31:24] = buffer_data_0[3983:3976];
        layer4[48][39:32] = buffer_data_0[3991:3984];
        layer0[49][7:0] = buffer_data_4[3967:3960];
        layer0[49][15:8] = buffer_data_4[3975:3968];
        layer0[49][23:16] = buffer_data_4[3983:3976];
        layer0[49][31:24] = buffer_data_4[3991:3984];
        layer0[49][39:32] = buffer_data_4[3999:3992];
        layer1[49][7:0] = buffer_data_3[3967:3960];
        layer1[49][15:8] = buffer_data_3[3975:3968];
        layer1[49][23:16] = buffer_data_3[3983:3976];
        layer1[49][31:24] = buffer_data_3[3991:3984];
        layer1[49][39:32] = buffer_data_3[3999:3992];
        layer2[49][7:0] = buffer_data_2[3967:3960];
        layer2[49][15:8] = buffer_data_2[3975:3968];
        layer2[49][23:16] = buffer_data_2[3983:3976];
        layer2[49][31:24] = buffer_data_2[3991:3984];
        layer2[49][39:32] = buffer_data_2[3999:3992];
        layer3[49][7:0] = buffer_data_1[3967:3960];
        layer3[49][15:8] = buffer_data_1[3975:3968];
        layer3[49][23:16] = buffer_data_1[3983:3976];
        layer3[49][31:24] = buffer_data_1[3991:3984];
        layer3[49][39:32] = buffer_data_1[3999:3992];
        layer4[49][7:0] = buffer_data_0[3967:3960];
        layer4[49][15:8] = buffer_data_0[3975:3968];
        layer4[49][23:16] = buffer_data_0[3983:3976];
        layer4[49][31:24] = buffer_data_0[3991:3984];
        layer4[49][39:32] = buffer_data_0[3999:3992];
        layer0[50][7:0] = buffer_data_4[3975:3968];
        layer0[50][15:8] = buffer_data_4[3983:3976];
        layer0[50][23:16] = buffer_data_4[3991:3984];
        layer0[50][31:24] = buffer_data_4[3999:3992];
        layer0[50][39:32] = buffer_data_4[4007:4000];
        layer1[50][7:0] = buffer_data_3[3975:3968];
        layer1[50][15:8] = buffer_data_3[3983:3976];
        layer1[50][23:16] = buffer_data_3[3991:3984];
        layer1[50][31:24] = buffer_data_3[3999:3992];
        layer1[50][39:32] = buffer_data_3[4007:4000];
        layer2[50][7:0] = buffer_data_2[3975:3968];
        layer2[50][15:8] = buffer_data_2[3983:3976];
        layer2[50][23:16] = buffer_data_2[3991:3984];
        layer2[50][31:24] = buffer_data_2[3999:3992];
        layer2[50][39:32] = buffer_data_2[4007:4000];
        layer3[50][7:0] = buffer_data_1[3975:3968];
        layer3[50][15:8] = buffer_data_1[3983:3976];
        layer3[50][23:16] = buffer_data_1[3991:3984];
        layer3[50][31:24] = buffer_data_1[3999:3992];
        layer3[50][39:32] = buffer_data_1[4007:4000];
        layer4[50][7:0] = buffer_data_0[3975:3968];
        layer4[50][15:8] = buffer_data_0[3983:3976];
        layer4[50][23:16] = buffer_data_0[3991:3984];
        layer4[50][31:24] = buffer_data_0[3999:3992];
        layer4[50][39:32] = buffer_data_0[4007:4000];
        layer0[51][7:0] = buffer_data_4[3983:3976];
        layer0[51][15:8] = buffer_data_4[3991:3984];
        layer0[51][23:16] = buffer_data_4[3999:3992];
        layer0[51][31:24] = buffer_data_4[4007:4000];
        layer0[51][39:32] = buffer_data_4[4015:4008];
        layer1[51][7:0] = buffer_data_3[3983:3976];
        layer1[51][15:8] = buffer_data_3[3991:3984];
        layer1[51][23:16] = buffer_data_3[3999:3992];
        layer1[51][31:24] = buffer_data_3[4007:4000];
        layer1[51][39:32] = buffer_data_3[4015:4008];
        layer2[51][7:0] = buffer_data_2[3983:3976];
        layer2[51][15:8] = buffer_data_2[3991:3984];
        layer2[51][23:16] = buffer_data_2[3999:3992];
        layer2[51][31:24] = buffer_data_2[4007:4000];
        layer2[51][39:32] = buffer_data_2[4015:4008];
        layer3[51][7:0] = buffer_data_1[3983:3976];
        layer3[51][15:8] = buffer_data_1[3991:3984];
        layer3[51][23:16] = buffer_data_1[3999:3992];
        layer3[51][31:24] = buffer_data_1[4007:4000];
        layer3[51][39:32] = buffer_data_1[4015:4008];
        layer4[51][7:0] = buffer_data_0[3983:3976];
        layer4[51][15:8] = buffer_data_0[3991:3984];
        layer4[51][23:16] = buffer_data_0[3999:3992];
        layer4[51][31:24] = buffer_data_0[4007:4000];
        layer4[51][39:32] = buffer_data_0[4015:4008];
        layer0[52][7:0] = buffer_data_4[3991:3984];
        layer0[52][15:8] = buffer_data_4[3999:3992];
        layer0[52][23:16] = buffer_data_4[4007:4000];
        layer0[52][31:24] = buffer_data_4[4015:4008];
        layer0[52][39:32] = buffer_data_4[4023:4016];
        layer1[52][7:0] = buffer_data_3[3991:3984];
        layer1[52][15:8] = buffer_data_3[3999:3992];
        layer1[52][23:16] = buffer_data_3[4007:4000];
        layer1[52][31:24] = buffer_data_3[4015:4008];
        layer1[52][39:32] = buffer_data_3[4023:4016];
        layer2[52][7:0] = buffer_data_2[3991:3984];
        layer2[52][15:8] = buffer_data_2[3999:3992];
        layer2[52][23:16] = buffer_data_2[4007:4000];
        layer2[52][31:24] = buffer_data_2[4015:4008];
        layer2[52][39:32] = buffer_data_2[4023:4016];
        layer3[52][7:0] = buffer_data_1[3991:3984];
        layer3[52][15:8] = buffer_data_1[3999:3992];
        layer3[52][23:16] = buffer_data_1[4007:4000];
        layer3[52][31:24] = buffer_data_1[4015:4008];
        layer3[52][39:32] = buffer_data_1[4023:4016];
        layer4[52][7:0] = buffer_data_0[3991:3984];
        layer4[52][15:8] = buffer_data_0[3999:3992];
        layer4[52][23:16] = buffer_data_0[4007:4000];
        layer4[52][31:24] = buffer_data_0[4015:4008];
        layer4[52][39:32] = buffer_data_0[4023:4016];
        layer0[53][7:0] = buffer_data_4[3999:3992];
        layer0[53][15:8] = buffer_data_4[4007:4000];
        layer0[53][23:16] = buffer_data_4[4015:4008];
        layer0[53][31:24] = buffer_data_4[4023:4016];
        layer0[53][39:32] = buffer_data_4[4031:4024];
        layer1[53][7:0] = buffer_data_3[3999:3992];
        layer1[53][15:8] = buffer_data_3[4007:4000];
        layer1[53][23:16] = buffer_data_3[4015:4008];
        layer1[53][31:24] = buffer_data_3[4023:4016];
        layer1[53][39:32] = buffer_data_3[4031:4024];
        layer2[53][7:0] = buffer_data_2[3999:3992];
        layer2[53][15:8] = buffer_data_2[4007:4000];
        layer2[53][23:16] = buffer_data_2[4015:4008];
        layer2[53][31:24] = buffer_data_2[4023:4016];
        layer2[53][39:32] = buffer_data_2[4031:4024];
        layer3[53][7:0] = buffer_data_1[3999:3992];
        layer3[53][15:8] = buffer_data_1[4007:4000];
        layer3[53][23:16] = buffer_data_1[4015:4008];
        layer3[53][31:24] = buffer_data_1[4023:4016];
        layer3[53][39:32] = buffer_data_1[4031:4024];
        layer4[53][7:0] = buffer_data_0[3999:3992];
        layer4[53][15:8] = buffer_data_0[4007:4000];
        layer4[53][23:16] = buffer_data_0[4015:4008];
        layer4[53][31:24] = buffer_data_0[4023:4016];
        layer4[53][39:32] = buffer_data_0[4031:4024];
        layer0[54][7:0] = buffer_data_4[4007:4000];
        layer0[54][15:8] = buffer_data_4[4015:4008];
        layer0[54][23:16] = buffer_data_4[4023:4016];
        layer0[54][31:24] = buffer_data_4[4031:4024];
        layer0[54][39:32] = buffer_data_4[4039:4032];
        layer1[54][7:0] = buffer_data_3[4007:4000];
        layer1[54][15:8] = buffer_data_3[4015:4008];
        layer1[54][23:16] = buffer_data_3[4023:4016];
        layer1[54][31:24] = buffer_data_3[4031:4024];
        layer1[54][39:32] = buffer_data_3[4039:4032];
        layer2[54][7:0] = buffer_data_2[4007:4000];
        layer2[54][15:8] = buffer_data_2[4015:4008];
        layer2[54][23:16] = buffer_data_2[4023:4016];
        layer2[54][31:24] = buffer_data_2[4031:4024];
        layer2[54][39:32] = buffer_data_2[4039:4032];
        layer3[54][7:0] = buffer_data_1[4007:4000];
        layer3[54][15:8] = buffer_data_1[4015:4008];
        layer3[54][23:16] = buffer_data_1[4023:4016];
        layer3[54][31:24] = buffer_data_1[4031:4024];
        layer3[54][39:32] = buffer_data_1[4039:4032];
        layer4[54][7:0] = buffer_data_0[4007:4000];
        layer4[54][15:8] = buffer_data_0[4015:4008];
        layer4[54][23:16] = buffer_data_0[4023:4016];
        layer4[54][31:24] = buffer_data_0[4031:4024];
        layer4[54][39:32] = buffer_data_0[4039:4032];
        layer0[55][7:0] = buffer_data_4[4015:4008];
        layer0[55][15:8] = buffer_data_4[4023:4016];
        layer0[55][23:16] = buffer_data_4[4031:4024];
        layer0[55][31:24] = buffer_data_4[4039:4032];
        layer0[55][39:32] = buffer_data_4[4047:4040];
        layer1[55][7:0] = buffer_data_3[4015:4008];
        layer1[55][15:8] = buffer_data_3[4023:4016];
        layer1[55][23:16] = buffer_data_3[4031:4024];
        layer1[55][31:24] = buffer_data_3[4039:4032];
        layer1[55][39:32] = buffer_data_3[4047:4040];
        layer2[55][7:0] = buffer_data_2[4015:4008];
        layer2[55][15:8] = buffer_data_2[4023:4016];
        layer2[55][23:16] = buffer_data_2[4031:4024];
        layer2[55][31:24] = buffer_data_2[4039:4032];
        layer2[55][39:32] = buffer_data_2[4047:4040];
        layer3[55][7:0] = buffer_data_1[4015:4008];
        layer3[55][15:8] = buffer_data_1[4023:4016];
        layer3[55][23:16] = buffer_data_1[4031:4024];
        layer3[55][31:24] = buffer_data_1[4039:4032];
        layer3[55][39:32] = buffer_data_1[4047:4040];
        layer4[55][7:0] = buffer_data_0[4015:4008];
        layer4[55][15:8] = buffer_data_0[4023:4016];
        layer4[55][23:16] = buffer_data_0[4031:4024];
        layer4[55][31:24] = buffer_data_0[4039:4032];
        layer4[55][39:32] = buffer_data_0[4047:4040];
        layer0[56][7:0] = buffer_data_4[4023:4016];
        layer0[56][15:8] = buffer_data_4[4031:4024];
        layer0[56][23:16] = buffer_data_4[4039:4032];
        layer0[56][31:24] = buffer_data_4[4047:4040];
        layer0[56][39:32] = buffer_data_4[4055:4048];
        layer1[56][7:0] = buffer_data_3[4023:4016];
        layer1[56][15:8] = buffer_data_3[4031:4024];
        layer1[56][23:16] = buffer_data_3[4039:4032];
        layer1[56][31:24] = buffer_data_3[4047:4040];
        layer1[56][39:32] = buffer_data_3[4055:4048];
        layer2[56][7:0] = buffer_data_2[4023:4016];
        layer2[56][15:8] = buffer_data_2[4031:4024];
        layer2[56][23:16] = buffer_data_2[4039:4032];
        layer2[56][31:24] = buffer_data_2[4047:4040];
        layer2[56][39:32] = buffer_data_2[4055:4048];
        layer3[56][7:0] = buffer_data_1[4023:4016];
        layer3[56][15:8] = buffer_data_1[4031:4024];
        layer3[56][23:16] = buffer_data_1[4039:4032];
        layer3[56][31:24] = buffer_data_1[4047:4040];
        layer3[56][39:32] = buffer_data_1[4055:4048];
        layer4[56][7:0] = buffer_data_0[4023:4016];
        layer4[56][15:8] = buffer_data_0[4031:4024];
        layer4[56][23:16] = buffer_data_0[4039:4032];
        layer4[56][31:24] = buffer_data_0[4047:4040];
        layer4[56][39:32] = buffer_data_0[4055:4048];
        layer0[57][7:0] = buffer_data_4[4031:4024];
        layer0[57][15:8] = buffer_data_4[4039:4032];
        layer0[57][23:16] = buffer_data_4[4047:4040];
        layer0[57][31:24] = buffer_data_4[4055:4048];
        layer0[57][39:32] = buffer_data_4[4063:4056];
        layer1[57][7:0] = buffer_data_3[4031:4024];
        layer1[57][15:8] = buffer_data_3[4039:4032];
        layer1[57][23:16] = buffer_data_3[4047:4040];
        layer1[57][31:24] = buffer_data_3[4055:4048];
        layer1[57][39:32] = buffer_data_3[4063:4056];
        layer2[57][7:0] = buffer_data_2[4031:4024];
        layer2[57][15:8] = buffer_data_2[4039:4032];
        layer2[57][23:16] = buffer_data_2[4047:4040];
        layer2[57][31:24] = buffer_data_2[4055:4048];
        layer2[57][39:32] = buffer_data_2[4063:4056];
        layer3[57][7:0] = buffer_data_1[4031:4024];
        layer3[57][15:8] = buffer_data_1[4039:4032];
        layer3[57][23:16] = buffer_data_1[4047:4040];
        layer3[57][31:24] = buffer_data_1[4055:4048];
        layer3[57][39:32] = buffer_data_1[4063:4056];
        layer4[57][7:0] = buffer_data_0[4031:4024];
        layer4[57][15:8] = buffer_data_0[4039:4032];
        layer4[57][23:16] = buffer_data_0[4047:4040];
        layer4[57][31:24] = buffer_data_0[4055:4048];
        layer4[57][39:32] = buffer_data_0[4063:4056];
        layer0[58][7:0] = buffer_data_4[4039:4032];
        layer0[58][15:8] = buffer_data_4[4047:4040];
        layer0[58][23:16] = buffer_data_4[4055:4048];
        layer0[58][31:24] = buffer_data_4[4063:4056];
        layer0[58][39:32] = buffer_data_4[4071:4064];
        layer1[58][7:0] = buffer_data_3[4039:4032];
        layer1[58][15:8] = buffer_data_3[4047:4040];
        layer1[58][23:16] = buffer_data_3[4055:4048];
        layer1[58][31:24] = buffer_data_3[4063:4056];
        layer1[58][39:32] = buffer_data_3[4071:4064];
        layer2[58][7:0] = buffer_data_2[4039:4032];
        layer2[58][15:8] = buffer_data_2[4047:4040];
        layer2[58][23:16] = buffer_data_2[4055:4048];
        layer2[58][31:24] = buffer_data_2[4063:4056];
        layer2[58][39:32] = buffer_data_2[4071:4064];
        layer3[58][7:0] = buffer_data_1[4039:4032];
        layer3[58][15:8] = buffer_data_1[4047:4040];
        layer3[58][23:16] = buffer_data_1[4055:4048];
        layer3[58][31:24] = buffer_data_1[4063:4056];
        layer3[58][39:32] = buffer_data_1[4071:4064];
        layer4[58][7:0] = buffer_data_0[4039:4032];
        layer4[58][15:8] = buffer_data_0[4047:4040];
        layer4[58][23:16] = buffer_data_0[4055:4048];
        layer4[58][31:24] = buffer_data_0[4063:4056];
        layer4[58][39:32] = buffer_data_0[4071:4064];
        layer0[59][7:0] = buffer_data_4[4047:4040];
        layer0[59][15:8] = buffer_data_4[4055:4048];
        layer0[59][23:16] = buffer_data_4[4063:4056];
        layer0[59][31:24] = buffer_data_4[4071:4064];
        layer0[59][39:32] = buffer_data_4[4079:4072];
        layer1[59][7:0] = buffer_data_3[4047:4040];
        layer1[59][15:8] = buffer_data_3[4055:4048];
        layer1[59][23:16] = buffer_data_3[4063:4056];
        layer1[59][31:24] = buffer_data_3[4071:4064];
        layer1[59][39:32] = buffer_data_3[4079:4072];
        layer2[59][7:0] = buffer_data_2[4047:4040];
        layer2[59][15:8] = buffer_data_2[4055:4048];
        layer2[59][23:16] = buffer_data_2[4063:4056];
        layer2[59][31:24] = buffer_data_2[4071:4064];
        layer2[59][39:32] = buffer_data_2[4079:4072];
        layer3[59][7:0] = buffer_data_1[4047:4040];
        layer3[59][15:8] = buffer_data_1[4055:4048];
        layer3[59][23:16] = buffer_data_1[4063:4056];
        layer3[59][31:24] = buffer_data_1[4071:4064];
        layer3[59][39:32] = buffer_data_1[4079:4072];
        layer4[59][7:0] = buffer_data_0[4047:4040];
        layer4[59][15:8] = buffer_data_0[4055:4048];
        layer4[59][23:16] = buffer_data_0[4063:4056];
        layer4[59][31:24] = buffer_data_0[4071:4064];
        layer4[59][39:32] = buffer_data_0[4079:4072];
        layer0[60][7:0] = buffer_data_4[4055:4048];
        layer0[60][15:8] = buffer_data_4[4063:4056];
        layer0[60][23:16] = buffer_data_4[4071:4064];
        layer0[60][31:24] = buffer_data_4[4079:4072];
        layer0[60][39:32] = buffer_data_4[4087:4080];
        layer1[60][7:0] = buffer_data_3[4055:4048];
        layer1[60][15:8] = buffer_data_3[4063:4056];
        layer1[60][23:16] = buffer_data_3[4071:4064];
        layer1[60][31:24] = buffer_data_3[4079:4072];
        layer1[60][39:32] = buffer_data_3[4087:4080];
        layer2[60][7:0] = buffer_data_2[4055:4048];
        layer2[60][15:8] = buffer_data_2[4063:4056];
        layer2[60][23:16] = buffer_data_2[4071:4064];
        layer2[60][31:24] = buffer_data_2[4079:4072];
        layer2[60][39:32] = buffer_data_2[4087:4080];
        layer3[60][7:0] = buffer_data_1[4055:4048];
        layer3[60][15:8] = buffer_data_1[4063:4056];
        layer3[60][23:16] = buffer_data_1[4071:4064];
        layer3[60][31:24] = buffer_data_1[4079:4072];
        layer3[60][39:32] = buffer_data_1[4087:4080];
        layer4[60][7:0] = buffer_data_0[4055:4048];
        layer4[60][15:8] = buffer_data_0[4063:4056];
        layer4[60][23:16] = buffer_data_0[4071:4064];
        layer4[60][31:24] = buffer_data_0[4079:4072];
        layer4[60][39:32] = buffer_data_0[4087:4080];
        layer0[61][7:0] = buffer_data_4[4063:4056];
        layer0[61][15:8] = buffer_data_4[4071:4064];
        layer0[61][23:16] = buffer_data_4[4079:4072];
        layer0[61][31:24] = buffer_data_4[4087:4080];
        layer0[61][39:32] = buffer_data_4[4095:4088];
        layer1[61][7:0] = buffer_data_3[4063:4056];
        layer1[61][15:8] = buffer_data_3[4071:4064];
        layer1[61][23:16] = buffer_data_3[4079:4072];
        layer1[61][31:24] = buffer_data_3[4087:4080];
        layer1[61][39:32] = buffer_data_3[4095:4088];
        layer2[61][7:0] = buffer_data_2[4063:4056];
        layer2[61][15:8] = buffer_data_2[4071:4064];
        layer2[61][23:16] = buffer_data_2[4079:4072];
        layer2[61][31:24] = buffer_data_2[4087:4080];
        layer2[61][39:32] = buffer_data_2[4095:4088];
        layer3[61][7:0] = buffer_data_1[4063:4056];
        layer3[61][15:8] = buffer_data_1[4071:4064];
        layer3[61][23:16] = buffer_data_1[4079:4072];
        layer3[61][31:24] = buffer_data_1[4087:4080];
        layer3[61][39:32] = buffer_data_1[4095:4088];
        layer4[61][7:0] = buffer_data_0[4063:4056];
        layer4[61][15:8] = buffer_data_0[4071:4064];
        layer4[61][23:16] = buffer_data_0[4079:4072];
        layer4[61][31:24] = buffer_data_0[4087:4080];
        layer4[61][39:32] = buffer_data_0[4095:4088];
        layer0[62][7:0] = buffer_data_4[4071:4064];
        layer0[62][15:8] = buffer_data_4[4079:4072];
        layer0[62][23:16] = buffer_data_4[4087:4080];
        layer0[62][31:24] = buffer_data_4[4095:4088];
        layer0[62][39:32] = buffer_data_4[4103:4096];
        layer1[62][7:0] = buffer_data_3[4071:4064];
        layer1[62][15:8] = buffer_data_3[4079:4072];
        layer1[62][23:16] = buffer_data_3[4087:4080];
        layer1[62][31:24] = buffer_data_3[4095:4088];
        layer1[62][39:32] = buffer_data_3[4103:4096];
        layer2[62][7:0] = buffer_data_2[4071:4064];
        layer2[62][15:8] = buffer_data_2[4079:4072];
        layer2[62][23:16] = buffer_data_2[4087:4080];
        layer2[62][31:24] = buffer_data_2[4095:4088];
        layer2[62][39:32] = buffer_data_2[4103:4096];
        layer3[62][7:0] = buffer_data_1[4071:4064];
        layer3[62][15:8] = buffer_data_1[4079:4072];
        layer3[62][23:16] = buffer_data_1[4087:4080];
        layer3[62][31:24] = buffer_data_1[4095:4088];
        layer3[62][39:32] = buffer_data_1[4103:4096];
        layer4[62][7:0] = buffer_data_0[4071:4064];
        layer4[62][15:8] = buffer_data_0[4079:4072];
        layer4[62][23:16] = buffer_data_0[4087:4080];
        layer4[62][31:24] = buffer_data_0[4095:4088];
        layer4[62][39:32] = buffer_data_0[4103:4096];
        layer0[63][7:0] = buffer_data_4[4079:4072];
        layer0[63][15:8] = buffer_data_4[4087:4080];
        layer0[63][23:16] = buffer_data_4[4095:4088];
        layer0[63][31:24] = buffer_data_4[4103:4096];
        layer0[63][39:32] = buffer_data_4[4111:4104];
        layer1[63][7:0] = buffer_data_3[4079:4072];
        layer1[63][15:8] = buffer_data_3[4087:4080];
        layer1[63][23:16] = buffer_data_3[4095:4088];
        layer1[63][31:24] = buffer_data_3[4103:4096];
        layer1[63][39:32] = buffer_data_3[4111:4104];
        layer2[63][7:0] = buffer_data_2[4079:4072];
        layer2[63][15:8] = buffer_data_2[4087:4080];
        layer2[63][23:16] = buffer_data_2[4095:4088];
        layer2[63][31:24] = buffer_data_2[4103:4096];
        layer2[63][39:32] = buffer_data_2[4111:4104];
        layer3[63][7:0] = buffer_data_1[4079:4072];
        layer3[63][15:8] = buffer_data_1[4087:4080];
        layer3[63][23:16] = buffer_data_1[4095:4088];
        layer3[63][31:24] = buffer_data_1[4103:4096];
        layer3[63][39:32] = buffer_data_1[4111:4104];
        layer4[63][7:0] = buffer_data_0[4079:4072];
        layer4[63][15:8] = buffer_data_0[4087:4080];
        layer4[63][23:16] = buffer_data_0[4095:4088];
        layer4[63][31:24] = buffer_data_0[4103:4096];
        layer4[63][39:32] = buffer_data_0[4111:4104];
    end
    ST_GAUSSIAN_8: begin
        layer0[0][7:0] = buffer_data_4[4087:4080];
        layer0[0][15:8] = buffer_data_4[4095:4088];
        layer0[0][23:16] = buffer_data_4[4103:4096];
        layer0[0][31:24] = buffer_data_4[4111:4104];
        layer0[0][39:32] = buffer_data_4[4119:4112];
        layer1[0][7:0] = buffer_data_3[4087:4080];
        layer1[0][15:8] = buffer_data_3[4095:4088];
        layer1[0][23:16] = buffer_data_3[4103:4096];
        layer1[0][31:24] = buffer_data_3[4111:4104];
        layer1[0][39:32] = buffer_data_3[4119:4112];
        layer2[0][7:0] = buffer_data_2[4087:4080];
        layer2[0][15:8] = buffer_data_2[4095:4088];
        layer2[0][23:16] = buffer_data_2[4103:4096];
        layer2[0][31:24] = buffer_data_2[4111:4104];
        layer2[0][39:32] = buffer_data_2[4119:4112];
        layer3[0][7:0] = buffer_data_1[4087:4080];
        layer3[0][15:8] = buffer_data_1[4095:4088];
        layer3[0][23:16] = buffer_data_1[4103:4096];
        layer3[0][31:24] = buffer_data_1[4111:4104];
        layer3[0][39:32] = buffer_data_1[4119:4112];
        layer4[0][7:0] = buffer_data_0[4087:4080];
        layer4[0][15:8] = buffer_data_0[4095:4088];
        layer4[0][23:16] = buffer_data_0[4103:4096];
        layer4[0][31:24] = buffer_data_0[4111:4104];
        layer4[0][39:32] = buffer_data_0[4119:4112];
        layer0[1][7:0] = buffer_data_4[4095:4088];
        layer0[1][15:8] = buffer_data_4[4103:4096];
        layer0[1][23:16] = buffer_data_4[4111:4104];
        layer0[1][31:24] = buffer_data_4[4119:4112];
        layer0[1][39:32] = buffer_data_4[4127:4120];
        layer1[1][7:0] = buffer_data_3[4095:4088];
        layer1[1][15:8] = buffer_data_3[4103:4096];
        layer1[1][23:16] = buffer_data_3[4111:4104];
        layer1[1][31:24] = buffer_data_3[4119:4112];
        layer1[1][39:32] = buffer_data_3[4127:4120];
        layer2[1][7:0] = buffer_data_2[4095:4088];
        layer2[1][15:8] = buffer_data_2[4103:4096];
        layer2[1][23:16] = buffer_data_2[4111:4104];
        layer2[1][31:24] = buffer_data_2[4119:4112];
        layer2[1][39:32] = buffer_data_2[4127:4120];
        layer3[1][7:0] = buffer_data_1[4095:4088];
        layer3[1][15:8] = buffer_data_1[4103:4096];
        layer3[1][23:16] = buffer_data_1[4111:4104];
        layer3[1][31:24] = buffer_data_1[4119:4112];
        layer3[1][39:32] = buffer_data_1[4127:4120];
        layer4[1][7:0] = buffer_data_0[4095:4088];
        layer4[1][15:8] = buffer_data_0[4103:4096];
        layer4[1][23:16] = buffer_data_0[4111:4104];
        layer4[1][31:24] = buffer_data_0[4119:4112];
        layer4[1][39:32] = buffer_data_0[4127:4120];
        layer0[2][7:0] = buffer_data_4[4103:4096];
        layer0[2][15:8] = buffer_data_4[4111:4104];
        layer0[2][23:16] = buffer_data_4[4119:4112];
        layer0[2][31:24] = buffer_data_4[4127:4120];
        layer0[2][39:32] = buffer_data_4[4135:4128];
        layer1[2][7:0] = buffer_data_3[4103:4096];
        layer1[2][15:8] = buffer_data_3[4111:4104];
        layer1[2][23:16] = buffer_data_3[4119:4112];
        layer1[2][31:24] = buffer_data_3[4127:4120];
        layer1[2][39:32] = buffer_data_3[4135:4128];
        layer2[2][7:0] = buffer_data_2[4103:4096];
        layer2[2][15:8] = buffer_data_2[4111:4104];
        layer2[2][23:16] = buffer_data_2[4119:4112];
        layer2[2][31:24] = buffer_data_2[4127:4120];
        layer2[2][39:32] = buffer_data_2[4135:4128];
        layer3[2][7:0] = buffer_data_1[4103:4096];
        layer3[2][15:8] = buffer_data_1[4111:4104];
        layer3[2][23:16] = buffer_data_1[4119:4112];
        layer3[2][31:24] = buffer_data_1[4127:4120];
        layer3[2][39:32] = buffer_data_1[4135:4128];
        layer4[2][7:0] = buffer_data_0[4103:4096];
        layer4[2][15:8] = buffer_data_0[4111:4104];
        layer4[2][23:16] = buffer_data_0[4119:4112];
        layer4[2][31:24] = buffer_data_0[4127:4120];
        layer4[2][39:32] = buffer_data_0[4135:4128];
        layer0[3][7:0] = buffer_data_4[4111:4104];
        layer0[3][15:8] = buffer_data_4[4119:4112];
        layer0[3][23:16] = buffer_data_4[4127:4120];
        layer0[3][31:24] = buffer_data_4[4135:4128];
        layer0[3][39:32] = buffer_data_4[4143:4136];
        layer1[3][7:0] = buffer_data_3[4111:4104];
        layer1[3][15:8] = buffer_data_3[4119:4112];
        layer1[3][23:16] = buffer_data_3[4127:4120];
        layer1[3][31:24] = buffer_data_3[4135:4128];
        layer1[3][39:32] = buffer_data_3[4143:4136];
        layer2[3][7:0] = buffer_data_2[4111:4104];
        layer2[3][15:8] = buffer_data_2[4119:4112];
        layer2[3][23:16] = buffer_data_2[4127:4120];
        layer2[3][31:24] = buffer_data_2[4135:4128];
        layer2[3][39:32] = buffer_data_2[4143:4136];
        layer3[3][7:0] = buffer_data_1[4111:4104];
        layer3[3][15:8] = buffer_data_1[4119:4112];
        layer3[3][23:16] = buffer_data_1[4127:4120];
        layer3[3][31:24] = buffer_data_1[4135:4128];
        layer3[3][39:32] = buffer_data_1[4143:4136];
        layer4[3][7:0] = buffer_data_0[4111:4104];
        layer4[3][15:8] = buffer_data_0[4119:4112];
        layer4[3][23:16] = buffer_data_0[4127:4120];
        layer4[3][31:24] = buffer_data_0[4135:4128];
        layer4[3][39:32] = buffer_data_0[4143:4136];
        layer0[4][7:0] = buffer_data_4[4119:4112];
        layer0[4][15:8] = buffer_data_4[4127:4120];
        layer0[4][23:16] = buffer_data_4[4135:4128];
        layer0[4][31:24] = buffer_data_4[4143:4136];
        layer0[4][39:32] = buffer_data_4[4151:4144];
        layer1[4][7:0] = buffer_data_3[4119:4112];
        layer1[4][15:8] = buffer_data_3[4127:4120];
        layer1[4][23:16] = buffer_data_3[4135:4128];
        layer1[4][31:24] = buffer_data_3[4143:4136];
        layer1[4][39:32] = buffer_data_3[4151:4144];
        layer2[4][7:0] = buffer_data_2[4119:4112];
        layer2[4][15:8] = buffer_data_2[4127:4120];
        layer2[4][23:16] = buffer_data_2[4135:4128];
        layer2[4][31:24] = buffer_data_2[4143:4136];
        layer2[4][39:32] = buffer_data_2[4151:4144];
        layer3[4][7:0] = buffer_data_1[4119:4112];
        layer3[4][15:8] = buffer_data_1[4127:4120];
        layer3[4][23:16] = buffer_data_1[4135:4128];
        layer3[4][31:24] = buffer_data_1[4143:4136];
        layer3[4][39:32] = buffer_data_1[4151:4144];
        layer4[4][7:0] = buffer_data_0[4119:4112];
        layer4[4][15:8] = buffer_data_0[4127:4120];
        layer4[4][23:16] = buffer_data_0[4135:4128];
        layer4[4][31:24] = buffer_data_0[4143:4136];
        layer4[4][39:32] = buffer_data_0[4151:4144];
        layer0[5][7:0] = buffer_data_4[4127:4120];
        layer0[5][15:8] = buffer_data_4[4135:4128];
        layer0[5][23:16] = buffer_data_4[4143:4136];
        layer0[5][31:24] = buffer_data_4[4151:4144];
        layer0[5][39:32] = buffer_data_4[4159:4152];
        layer1[5][7:0] = buffer_data_3[4127:4120];
        layer1[5][15:8] = buffer_data_3[4135:4128];
        layer1[5][23:16] = buffer_data_3[4143:4136];
        layer1[5][31:24] = buffer_data_3[4151:4144];
        layer1[5][39:32] = buffer_data_3[4159:4152];
        layer2[5][7:0] = buffer_data_2[4127:4120];
        layer2[5][15:8] = buffer_data_2[4135:4128];
        layer2[5][23:16] = buffer_data_2[4143:4136];
        layer2[5][31:24] = buffer_data_2[4151:4144];
        layer2[5][39:32] = buffer_data_2[4159:4152];
        layer3[5][7:0] = buffer_data_1[4127:4120];
        layer3[5][15:8] = buffer_data_1[4135:4128];
        layer3[5][23:16] = buffer_data_1[4143:4136];
        layer3[5][31:24] = buffer_data_1[4151:4144];
        layer3[5][39:32] = buffer_data_1[4159:4152];
        layer4[5][7:0] = buffer_data_0[4127:4120];
        layer4[5][15:8] = buffer_data_0[4135:4128];
        layer4[5][23:16] = buffer_data_0[4143:4136];
        layer4[5][31:24] = buffer_data_0[4151:4144];
        layer4[5][39:32] = buffer_data_0[4159:4152];
        layer0[6][7:0] = buffer_data_4[4135:4128];
        layer0[6][15:8] = buffer_data_4[4143:4136];
        layer0[6][23:16] = buffer_data_4[4151:4144];
        layer0[6][31:24] = buffer_data_4[4159:4152];
        layer0[6][39:32] = buffer_data_4[4167:4160];
        layer1[6][7:0] = buffer_data_3[4135:4128];
        layer1[6][15:8] = buffer_data_3[4143:4136];
        layer1[6][23:16] = buffer_data_3[4151:4144];
        layer1[6][31:24] = buffer_data_3[4159:4152];
        layer1[6][39:32] = buffer_data_3[4167:4160];
        layer2[6][7:0] = buffer_data_2[4135:4128];
        layer2[6][15:8] = buffer_data_2[4143:4136];
        layer2[6][23:16] = buffer_data_2[4151:4144];
        layer2[6][31:24] = buffer_data_2[4159:4152];
        layer2[6][39:32] = buffer_data_2[4167:4160];
        layer3[6][7:0] = buffer_data_1[4135:4128];
        layer3[6][15:8] = buffer_data_1[4143:4136];
        layer3[6][23:16] = buffer_data_1[4151:4144];
        layer3[6][31:24] = buffer_data_1[4159:4152];
        layer3[6][39:32] = buffer_data_1[4167:4160];
        layer4[6][7:0] = buffer_data_0[4135:4128];
        layer4[6][15:8] = buffer_data_0[4143:4136];
        layer4[6][23:16] = buffer_data_0[4151:4144];
        layer4[6][31:24] = buffer_data_0[4159:4152];
        layer4[6][39:32] = buffer_data_0[4167:4160];
        layer0[7][7:0] = buffer_data_4[4143:4136];
        layer0[7][15:8] = buffer_data_4[4151:4144];
        layer0[7][23:16] = buffer_data_4[4159:4152];
        layer0[7][31:24] = buffer_data_4[4167:4160];
        layer0[7][39:32] = buffer_data_4[4175:4168];
        layer1[7][7:0] = buffer_data_3[4143:4136];
        layer1[7][15:8] = buffer_data_3[4151:4144];
        layer1[7][23:16] = buffer_data_3[4159:4152];
        layer1[7][31:24] = buffer_data_3[4167:4160];
        layer1[7][39:32] = buffer_data_3[4175:4168];
        layer2[7][7:0] = buffer_data_2[4143:4136];
        layer2[7][15:8] = buffer_data_2[4151:4144];
        layer2[7][23:16] = buffer_data_2[4159:4152];
        layer2[7][31:24] = buffer_data_2[4167:4160];
        layer2[7][39:32] = buffer_data_2[4175:4168];
        layer3[7][7:0] = buffer_data_1[4143:4136];
        layer3[7][15:8] = buffer_data_1[4151:4144];
        layer3[7][23:16] = buffer_data_1[4159:4152];
        layer3[7][31:24] = buffer_data_1[4167:4160];
        layer3[7][39:32] = buffer_data_1[4175:4168];
        layer4[7][7:0] = buffer_data_0[4143:4136];
        layer4[7][15:8] = buffer_data_0[4151:4144];
        layer4[7][23:16] = buffer_data_0[4159:4152];
        layer4[7][31:24] = buffer_data_0[4167:4160];
        layer4[7][39:32] = buffer_data_0[4175:4168];
        layer0[8][7:0] = buffer_data_4[4151:4144];
        layer0[8][15:8] = buffer_data_4[4159:4152];
        layer0[8][23:16] = buffer_data_4[4167:4160];
        layer0[8][31:24] = buffer_data_4[4175:4168];
        layer0[8][39:32] = buffer_data_4[4183:4176];
        layer1[8][7:0] = buffer_data_3[4151:4144];
        layer1[8][15:8] = buffer_data_3[4159:4152];
        layer1[8][23:16] = buffer_data_3[4167:4160];
        layer1[8][31:24] = buffer_data_3[4175:4168];
        layer1[8][39:32] = buffer_data_3[4183:4176];
        layer2[8][7:0] = buffer_data_2[4151:4144];
        layer2[8][15:8] = buffer_data_2[4159:4152];
        layer2[8][23:16] = buffer_data_2[4167:4160];
        layer2[8][31:24] = buffer_data_2[4175:4168];
        layer2[8][39:32] = buffer_data_2[4183:4176];
        layer3[8][7:0] = buffer_data_1[4151:4144];
        layer3[8][15:8] = buffer_data_1[4159:4152];
        layer3[8][23:16] = buffer_data_1[4167:4160];
        layer3[8][31:24] = buffer_data_1[4175:4168];
        layer3[8][39:32] = buffer_data_1[4183:4176];
        layer4[8][7:0] = buffer_data_0[4151:4144];
        layer4[8][15:8] = buffer_data_0[4159:4152];
        layer4[8][23:16] = buffer_data_0[4167:4160];
        layer4[8][31:24] = buffer_data_0[4175:4168];
        layer4[8][39:32] = buffer_data_0[4183:4176];
        layer0[9][7:0] = buffer_data_4[4159:4152];
        layer0[9][15:8] = buffer_data_4[4167:4160];
        layer0[9][23:16] = buffer_data_4[4175:4168];
        layer0[9][31:24] = buffer_data_4[4183:4176];
        layer0[9][39:32] = buffer_data_4[4191:4184];
        layer1[9][7:0] = buffer_data_3[4159:4152];
        layer1[9][15:8] = buffer_data_3[4167:4160];
        layer1[9][23:16] = buffer_data_3[4175:4168];
        layer1[9][31:24] = buffer_data_3[4183:4176];
        layer1[9][39:32] = buffer_data_3[4191:4184];
        layer2[9][7:0] = buffer_data_2[4159:4152];
        layer2[9][15:8] = buffer_data_2[4167:4160];
        layer2[9][23:16] = buffer_data_2[4175:4168];
        layer2[9][31:24] = buffer_data_2[4183:4176];
        layer2[9][39:32] = buffer_data_2[4191:4184];
        layer3[9][7:0] = buffer_data_1[4159:4152];
        layer3[9][15:8] = buffer_data_1[4167:4160];
        layer3[9][23:16] = buffer_data_1[4175:4168];
        layer3[9][31:24] = buffer_data_1[4183:4176];
        layer3[9][39:32] = buffer_data_1[4191:4184];
        layer4[9][7:0] = buffer_data_0[4159:4152];
        layer4[9][15:8] = buffer_data_0[4167:4160];
        layer4[9][23:16] = buffer_data_0[4175:4168];
        layer4[9][31:24] = buffer_data_0[4183:4176];
        layer4[9][39:32] = buffer_data_0[4191:4184];
        layer0[10][7:0] = buffer_data_4[4167:4160];
        layer0[10][15:8] = buffer_data_4[4175:4168];
        layer0[10][23:16] = buffer_data_4[4183:4176];
        layer0[10][31:24] = buffer_data_4[4191:4184];
        layer0[10][39:32] = buffer_data_4[4199:4192];
        layer1[10][7:0] = buffer_data_3[4167:4160];
        layer1[10][15:8] = buffer_data_3[4175:4168];
        layer1[10][23:16] = buffer_data_3[4183:4176];
        layer1[10][31:24] = buffer_data_3[4191:4184];
        layer1[10][39:32] = buffer_data_3[4199:4192];
        layer2[10][7:0] = buffer_data_2[4167:4160];
        layer2[10][15:8] = buffer_data_2[4175:4168];
        layer2[10][23:16] = buffer_data_2[4183:4176];
        layer2[10][31:24] = buffer_data_2[4191:4184];
        layer2[10][39:32] = buffer_data_2[4199:4192];
        layer3[10][7:0] = buffer_data_1[4167:4160];
        layer3[10][15:8] = buffer_data_1[4175:4168];
        layer3[10][23:16] = buffer_data_1[4183:4176];
        layer3[10][31:24] = buffer_data_1[4191:4184];
        layer3[10][39:32] = buffer_data_1[4199:4192];
        layer4[10][7:0] = buffer_data_0[4167:4160];
        layer4[10][15:8] = buffer_data_0[4175:4168];
        layer4[10][23:16] = buffer_data_0[4183:4176];
        layer4[10][31:24] = buffer_data_0[4191:4184];
        layer4[10][39:32] = buffer_data_0[4199:4192];
        layer0[11][7:0] = buffer_data_4[4175:4168];
        layer0[11][15:8] = buffer_data_4[4183:4176];
        layer0[11][23:16] = buffer_data_4[4191:4184];
        layer0[11][31:24] = buffer_data_4[4199:4192];
        layer0[11][39:32] = buffer_data_4[4207:4200];
        layer1[11][7:0] = buffer_data_3[4175:4168];
        layer1[11][15:8] = buffer_data_3[4183:4176];
        layer1[11][23:16] = buffer_data_3[4191:4184];
        layer1[11][31:24] = buffer_data_3[4199:4192];
        layer1[11][39:32] = buffer_data_3[4207:4200];
        layer2[11][7:0] = buffer_data_2[4175:4168];
        layer2[11][15:8] = buffer_data_2[4183:4176];
        layer2[11][23:16] = buffer_data_2[4191:4184];
        layer2[11][31:24] = buffer_data_2[4199:4192];
        layer2[11][39:32] = buffer_data_2[4207:4200];
        layer3[11][7:0] = buffer_data_1[4175:4168];
        layer3[11][15:8] = buffer_data_1[4183:4176];
        layer3[11][23:16] = buffer_data_1[4191:4184];
        layer3[11][31:24] = buffer_data_1[4199:4192];
        layer3[11][39:32] = buffer_data_1[4207:4200];
        layer4[11][7:0] = buffer_data_0[4175:4168];
        layer4[11][15:8] = buffer_data_0[4183:4176];
        layer4[11][23:16] = buffer_data_0[4191:4184];
        layer4[11][31:24] = buffer_data_0[4199:4192];
        layer4[11][39:32] = buffer_data_0[4207:4200];
        layer0[12][7:0] = buffer_data_4[4183:4176];
        layer0[12][15:8] = buffer_data_4[4191:4184];
        layer0[12][23:16] = buffer_data_4[4199:4192];
        layer0[12][31:24] = buffer_data_4[4207:4200];
        layer0[12][39:32] = buffer_data_4[4215:4208];
        layer1[12][7:0] = buffer_data_3[4183:4176];
        layer1[12][15:8] = buffer_data_3[4191:4184];
        layer1[12][23:16] = buffer_data_3[4199:4192];
        layer1[12][31:24] = buffer_data_3[4207:4200];
        layer1[12][39:32] = buffer_data_3[4215:4208];
        layer2[12][7:0] = buffer_data_2[4183:4176];
        layer2[12][15:8] = buffer_data_2[4191:4184];
        layer2[12][23:16] = buffer_data_2[4199:4192];
        layer2[12][31:24] = buffer_data_2[4207:4200];
        layer2[12][39:32] = buffer_data_2[4215:4208];
        layer3[12][7:0] = buffer_data_1[4183:4176];
        layer3[12][15:8] = buffer_data_1[4191:4184];
        layer3[12][23:16] = buffer_data_1[4199:4192];
        layer3[12][31:24] = buffer_data_1[4207:4200];
        layer3[12][39:32] = buffer_data_1[4215:4208];
        layer4[12][7:0] = buffer_data_0[4183:4176];
        layer4[12][15:8] = buffer_data_0[4191:4184];
        layer4[12][23:16] = buffer_data_0[4199:4192];
        layer4[12][31:24] = buffer_data_0[4207:4200];
        layer4[12][39:32] = buffer_data_0[4215:4208];
        layer0[13][7:0] = buffer_data_4[4191:4184];
        layer0[13][15:8] = buffer_data_4[4199:4192];
        layer0[13][23:16] = buffer_data_4[4207:4200];
        layer0[13][31:24] = buffer_data_4[4215:4208];
        layer0[13][39:32] = buffer_data_4[4223:4216];
        layer1[13][7:0] = buffer_data_3[4191:4184];
        layer1[13][15:8] = buffer_data_3[4199:4192];
        layer1[13][23:16] = buffer_data_3[4207:4200];
        layer1[13][31:24] = buffer_data_3[4215:4208];
        layer1[13][39:32] = buffer_data_3[4223:4216];
        layer2[13][7:0] = buffer_data_2[4191:4184];
        layer2[13][15:8] = buffer_data_2[4199:4192];
        layer2[13][23:16] = buffer_data_2[4207:4200];
        layer2[13][31:24] = buffer_data_2[4215:4208];
        layer2[13][39:32] = buffer_data_2[4223:4216];
        layer3[13][7:0] = buffer_data_1[4191:4184];
        layer3[13][15:8] = buffer_data_1[4199:4192];
        layer3[13][23:16] = buffer_data_1[4207:4200];
        layer3[13][31:24] = buffer_data_1[4215:4208];
        layer3[13][39:32] = buffer_data_1[4223:4216];
        layer4[13][7:0] = buffer_data_0[4191:4184];
        layer4[13][15:8] = buffer_data_0[4199:4192];
        layer4[13][23:16] = buffer_data_0[4207:4200];
        layer4[13][31:24] = buffer_data_0[4215:4208];
        layer4[13][39:32] = buffer_data_0[4223:4216];
        layer0[14][7:0] = buffer_data_4[4199:4192];
        layer0[14][15:8] = buffer_data_4[4207:4200];
        layer0[14][23:16] = buffer_data_4[4215:4208];
        layer0[14][31:24] = buffer_data_4[4223:4216];
        layer0[14][39:32] = buffer_data_4[4231:4224];
        layer1[14][7:0] = buffer_data_3[4199:4192];
        layer1[14][15:8] = buffer_data_3[4207:4200];
        layer1[14][23:16] = buffer_data_3[4215:4208];
        layer1[14][31:24] = buffer_data_3[4223:4216];
        layer1[14][39:32] = buffer_data_3[4231:4224];
        layer2[14][7:0] = buffer_data_2[4199:4192];
        layer2[14][15:8] = buffer_data_2[4207:4200];
        layer2[14][23:16] = buffer_data_2[4215:4208];
        layer2[14][31:24] = buffer_data_2[4223:4216];
        layer2[14][39:32] = buffer_data_2[4231:4224];
        layer3[14][7:0] = buffer_data_1[4199:4192];
        layer3[14][15:8] = buffer_data_1[4207:4200];
        layer3[14][23:16] = buffer_data_1[4215:4208];
        layer3[14][31:24] = buffer_data_1[4223:4216];
        layer3[14][39:32] = buffer_data_1[4231:4224];
        layer4[14][7:0] = buffer_data_0[4199:4192];
        layer4[14][15:8] = buffer_data_0[4207:4200];
        layer4[14][23:16] = buffer_data_0[4215:4208];
        layer4[14][31:24] = buffer_data_0[4223:4216];
        layer4[14][39:32] = buffer_data_0[4231:4224];
        layer0[15][7:0] = buffer_data_4[4207:4200];
        layer0[15][15:8] = buffer_data_4[4215:4208];
        layer0[15][23:16] = buffer_data_4[4223:4216];
        layer0[15][31:24] = buffer_data_4[4231:4224];
        layer0[15][39:32] = buffer_data_4[4239:4232];
        layer1[15][7:0] = buffer_data_3[4207:4200];
        layer1[15][15:8] = buffer_data_3[4215:4208];
        layer1[15][23:16] = buffer_data_3[4223:4216];
        layer1[15][31:24] = buffer_data_3[4231:4224];
        layer1[15][39:32] = buffer_data_3[4239:4232];
        layer2[15][7:0] = buffer_data_2[4207:4200];
        layer2[15][15:8] = buffer_data_2[4215:4208];
        layer2[15][23:16] = buffer_data_2[4223:4216];
        layer2[15][31:24] = buffer_data_2[4231:4224];
        layer2[15][39:32] = buffer_data_2[4239:4232];
        layer3[15][7:0] = buffer_data_1[4207:4200];
        layer3[15][15:8] = buffer_data_1[4215:4208];
        layer3[15][23:16] = buffer_data_1[4223:4216];
        layer3[15][31:24] = buffer_data_1[4231:4224];
        layer3[15][39:32] = buffer_data_1[4239:4232];
        layer4[15][7:0] = buffer_data_0[4207:4200];
        layer4[15][15:8] = buffer_data_0[4215:4208];
        layer4[15][23:16] = buffer_data_0[4223:4216];
        layer4[15][31:24] = buffer_data_0[4231:4224];
        layer4[15][39:32] = buffer_data_0[4239:4232];
        layer0[16][7:0] = buffer_data_4[4215:4208];
        layer0[16][15:8] = buffer_data_4[4223:4216];
        layer0[16][23:16] = buffer_data_4[4231:4224];
        layer0[16][31:24] = buffer_data_4[4239:4232];
        layer0[16][39:32] = buffer_data_4[4247:4240];
        layer1[16][7:0] = buffer_data_3[4215:4208];
        layer1[16][15:8] = buffer_data_3[4223:4216];
        layer1[16][23:16] = buffer_data_3[4231:4224];
        layer1[16][31:24] = buffer_data_3[4239:4232];
        layer1[16][39:32] = buffer_data_3[4247:4240];
        layer2[16][7:0] = buffer_data_2[4215:4208];
        layer2[16][15:8] = buffer_data_2[4223:4216];
        layer2[16][23:16] = buffer_data_2[4231:4224];
        layer2[16][31:24] = buffer_data_2[4239:4232];
        layer2[16][39:32] = buffer_data_2[4247:4240];
        layer3[16][7:0] = buffer_data_1[4215:4208];
        layer3[16][15:8] = buffer_data_1[4223:4216];
        layer3[16][23:16] = buffer_data_1[4231:4224];
        layer3[16][31:24] = buffer_data_1[4239:4232];
        layer3[16][39:32] = buffer_data_1[4247:4240];
        layer4[16][7:0] = buffer_data_0[4215:4208];
        layer4[16][15:8] = buffer_data_0[4223:4216];
        layer4[16][23:16] = buffer_data_0[4231:4224];
        layer4[16][31:24] = buffer_data_0[4239:4232];
        layer4[16][39:32] = buffer_data_0[4247:4240];
        layer0[17][7:0] = buffer_data_4[4223:4216];
        layer0[17][15:8] = buffer_data_4[4231:4224];
        layer0[17][23:16] = buffer_data_4[4239:4232];
        layer0[17][31:24] = buffer_data_4[4247:4240];
        layer0[17][39:32] = buffer_data_4[4255:4248];
        layer1[17][7:0] = buffer_data_3[4223:4216];
        layer1[17][15:8] = buffer_data_3[4231:4224];
        layer1[17][23:16] = buffer_data_3[4239:4232];
        layer1[17][31:24] = buffer_data_3[4247:4240];
        layer1[17][39:32] = buffer_data_3[4255:4248];
        layer2[17][7:0] = buffer_data_2[4223:4216];
        layer2[17][15:8] = buffer_data_2[4231:4224];
        layer2[17][23:16] = buffer_data_2[4239:4232];
        layer2[17][31:24] = buffer_data_2[4247:4240];
        layer2[17][39:32] = buffer_data_2[4255:4248];
        layer3[17][7:0] = buffer_data_1[4223:4216];
        layer3[17][15:8] = buffer_data_1[4231:4224];
        layer3[17][23:16] = buffer_data_1[4239:4232];
        layer3[17][31:24] = buffer_data_1[4247:4240];
        layer3[17][39:32] = buffer_data_1[4255:4248];
        layer4[17][7:0] = buffer_data_0[4223:4216];
        layer4[17][15:8] = buffer_data_0[4231:4224];
        layer4[17][23:16] = buffer_data_0[4239:4232];
        layer4[17][31:24] = buffer_data_0[4247:4240];
        layer4[17][39:32] = buffer_data_0[4255:4248];
        layer0[18][7:0] = buffer_data_4[4231:4224];
        layer0[18][15:8] = buffer_data_4[4239:4232];
        layer0[18][23:16] = buffer_data_4[4247:4240];
        layer0[18][31:24] = buffer_data_4[4255:4248];
        layer0[18][39:32] = buffer_data_4[4263:4256];
        layer1[18][7:0] = buffer_data_3[4231:4224];
        layer1[18][15:8] = buffer_data_3[4239:4232];
        layer1[18][23:16] = buffer_data_3[4247:4240];
        layer1[18][31:24] = buffer_data_3[4255:4248];
        layer1[18][39:32] = buffer_data_3[4263:4256];
        layer2[18][7:0] = buffer_data_2[4231:4224];
        layer2[18][15:8] = buffer_data_2[4239:4232];
        layer2[18][23:16] = buffer_data_2[4247:4240];
        layer2[18][31:24] = buffer_data_2[4255:4248];
        layer2[18][39:32] = buffer_data_2[4263:4256];
        layer3[18][7:0] = buffer_data_1[4231:4224];
        layer3[18][15:8] = buffer_data_1[4239:4232];
        layer3[18][23:16] = buffer_data_1[4247:4240];
        layer3[18][31:24] = buffer_data_1[4255:4248];
        layer3[18][39:32] = buffer_data_1[4263:4256];
        layer4[18][7:0] = buffer_data_0[4231:4224];
        layer4[18][15:8] = buffer_data_0[4239:4232];
        layer4[18][23:16] = buffer_data_0[4247:4240];
        layer4[18][31:24] = buffer_data_0[4255:4248];
        layer4[18][39:32] = buffer_data_0[4263:4256];
        layer0[19][7:0] = buffer_data_4[4239:4232];
        layer0[19][15:8] = buffer_data_4[4247:4240];
        layer0[19][23:16] = buffer_data_4[4255:4248];
        layer0[19][31:24] = buffer_data_4[4263:4256];
        layer0[19][39:32] = buffer_data_4[4271:4264];
        layer1[19][7:0] = buffer_data_3[4239:4232];
        layer1[19][15:8] = buffer_data_3[4247:4240];
        layer1[19][23:16] = buffer_data_3[4255:4248];
        layer1[19][31:24] = buffer_data_3[4263:4256];
        layer1[19][39:32] = buffer_data_3[4271:4264];
        layer2[19][7:0] = buffer_data_2[4239:4232];
        layer2[19][15:8] = buffer_data_2[4247:4240];
        layer2[19][23:16] = buffer_data_2[4255:4248];
        layer2[19][31:24] = buffer_data_2[4263:4256];
        layer2[19][39:32] = buffer_data_2[4271:4264];
        layer3[19][7:0] = buffer_data_1[4239:4232];
        layer3[19][15:8] = buffer_data_1[4247:4240];
        layer3[19][23:16] = buffer_data_1[4255:4248];
        layer3[19][31:24] = buffer_data_1[4263:4256];
        layer3[19][39:32] = buffer_data_1[4271:4264];
        layer4[19][7:0] = buffer_data_0[4239:4232];
        layer4[19][15:8] = buffer_data_0[4247:4240];
        layer4[19][23:16] = buffer_data_0[4255:4248];
        layer4[19][31:24] = buffer_data_0[4263:4256];
        layer4[19][39:32] = buffer_data_0[4271:4264];
        layer0[20][7:0] = buffer_data_4[4247:4240];
        layer0[20][15:8] = buffer_data_4[4255:4248];
        layer0[20][23:16] = buffer_data_4[4263:4256];
        layer0[20][31:24] = buffer_data_4[4271:4264];
        layer0[20][39:32] = buffer_data_4[4279:4272];
        layer1[20][7:0] = buffer_data_3[4247:4240];
        layer1[20][15:8] = buffer_data_3[4255:4248];
        layer1[20][23:16] = buffer_data_3[4263:4256];
        layer1[20][31:24] = buffer_data_3[4271:4264];
        layer1[20][39:32] = buffer_data_3[4279:4272];
        layer2[20][7:0] = buffer_data_2[4247:4240];
        layer2[20][15:8] = buffer_data_2[4255:4248];
        layer2[20][23:16] = buffer_data_2[4263:4256];
        layer2[20][31:24] = buffer_data_2[4271:4264];
        layer2[20][39:32] = buffer_data_2[4279:4272];
        layer3[20][7:0] = buffer_data_1[4247:4240];
        layer3[20][15:8] = buffer_data_1[4255:4248];
        layer3[20][23:16] = buffer_data_1[4263:4256];
        layer3[20][31:24] = buffer_data_1[4271:4264];
        layer3[20][39:32] = buffer_data_1[4279:4272];
        layer4[20][7:0] = buffer_data_0[4247:4240];
        layer4[20][15:8] = buffer_data_0[4255:4248];
        layer4[20][23:16] = buffer_data_0[4263:4256];
        layer4[20][31:24] = buffer_data_0[4271:4264];
        layer4[20][39:32] = buffer_data_0[4279:4272];
        layer0[21][7:0] = buffer_data_4[4255:4248];
        layer0[21][15:8] = buffer_data_4[4263:4256];
        layer0[21][23:16] = buffer_data_4[4271:4264];
        layer0[21][31:24] = buffer_data_4[4279:4272];
        layer0[21][39:32] = buffer_data_4[4287:4280];
        layer1[21][7:0] = buffer_data_3[4255:4248];
        layer1[21][15:8] = buffer_data_3[4263:4256];
        layer1[21][23:16] = buffer_data_3[4271:4264];
        layer1[21][31:24] = buffer_data_3[4279:4272];
        layer1[21][39:32] = buffer_data_3[4287:4280];
        layer2[21][7:0] = buffer_data_2[4255:4248];
        layer2[21][15:8] = buffer_data_2[4263:4256];
        layer2[21][23:16] = buffer_data_2[4271:4264];
        layer2[21][31:24] = buffer_data_2[4279:4272];
        layer2[21][39:32] = buffer_data_2[4287:4280];
        layer3[21][7:0] = buffer_data_1[4255:4248];
        layer3[21][15:8] = buffer_data_1[4263:4256];
        layer3[21][23:16] = buffer_data_1[4271:4264];
        layer3[21][31:24] = buffer_data_1[4279:4272];
        layer3[21][39:32] = buffer_data_1[4287:4280];
        layer4[21][7:0] = buffer_data_0[4255:4248];
        layer4[21][15:8] = buffer_data_0[4263:4256];
        layer4[21][23:16] = buffer_data_0[4271:4264];
        layer4[21][31:24] = buffer_data_0[4279:4272];
        layer4[21][39:32] = buffer_data_0[4287:4280];
        layer0[22][7:0] = buffer_data_4[4263:4256];
        layer0[22][15:8] = buffer_data_4[4271:4264];
        layer0[22][23:16] = buffer_data_4[4279:4272];
        layer0[22][31:24] = buffer_data_4[4287:4280];
        layer0[22][39:32] = buffer_data_4[4295:4288];
        layer1[22][7:0] = buffer_data_3[4263:4256];
        layer1[22][15:8] = buffer_data_3[4271:4264];
        layer1[22][23:16] = buffer_data_3[4279:4272];
        layer1[22][31:24] = buffer_data_3[4287:4280];
        layer1[22][39:32] = buffer_data_3[4295:4288];
        layer2[22][7:0] = buffer_data_2[4263:4256];
        layer2[22][15:8] = buffer_data_2[4271:4264];
        layer2[22][23:16] = buffer_data_2[4279:4272];
        layer2[22][31:24] = buffer_data_2[4287:4280];
        layer2[22][39:32] = buffer_data_2[4295:4288];
        layer3[22][7:0] = buffer_data_1[4263:4256];
        layer3[22][15:8] = buffer_data_1[4271:4264];
        layer3[22][23:16] = buffer_data_1[4279:4272];
        layer3[22][31:24] = buffer_data_1[4287:4280];
        layer3[22][39:32] = buffer_data_1[4295:4288];
        layer4[22][7:0] = buffer_data_0[4263:4256];
        layer4[22][15:8] = buffer_data_0[4271:4264];
        layer4[22][23:16] = buffer_data_0[4279:4272];
        layer4[22][31:24] = buffer_data_0[4287:4280];
        layer4[22][39:32] = buffer_data_0[4295:4288];
        layer0[23][7:0] = buffer_data_4[4271:4264];
        layer0[23][15:8] = buffer_data_4[4279:4272];
        layer0[23][23:16] = buffer_data_4[4287:4280];
        layer0[23][31:24] = buffer_data_4[4295:4288];
        layer0[23][39:32] = buffer_data_4[4303:4296];
        layer1[23][7:0] = buffer_data_3[4271:4264];
        layer1[23][15:8] = buffer_data_3[4279:4272];
        layer1[23][23:16] = buffer_data_3[4287:4280];
        layer1[23][31:24] = buffer_data_3[4295:4288];
        layer1[23][39:32] = buffer_data_3[4303:4296];
        layer2[23][7:0] = buffer_data_2[4271:4264];
        layer2[23][15:8] = buffer_data_2[4279:4272];
        layer2[23][23:16] = buffer_data_2[4287:4280];
        layer2[23][31:24] = buffer_data_2[4295:4288];
        layer2[23][39:32] = buffer_data_2[4303:4296];
        layer3[23][7:0] = buffer_data_1[4271:4264];
        layer3[23][15:8] = buffer_data_1[4279:4272];
        layer3[23][23:16] = buffer_data_1[4287:4280];
        layer3[23][31:24] = buffer_data_1[4295:4288];
        layer3[23][39:32] = buffer_data_1[4303:4296];
        layer4[23][7:0] = buffer_data_0[4271:4264];
        layer4[23][15:8] = buffer_data_0[4279:4272];
        layer4[23][23:16] = buffer_data_0[4287:4280];
        layer4[23][31:24] = buffer_data_0[4295:4288];
        layer4[23][39:32] = buffer_data_0[4303:4296];
        layer0[24][7:0] = buffer_data_4[4279:4272];
        layer0[24][15:8] = buffer_data_4[4287:4280];
        layer0[24][23:16] = buffer_data_4[4295:4288];
        layer0[24][31:24] = buffer_data_4[4303:4296];
        layer0[24][39:32] = buffer_data_4[4311:4304];
        layer1[24][7:0] = buffer_data_3[4279:4272];
        layer1[24][15:8] = buffer_data_3[4287:4280];
        layer1[24][23:16] = buffer_data_3[4295:4288];
        layer1[24][31:24] = buffer_data_3[4303:4296];
        layer1[24][39:32] = buffer_data_3[4311:4304];
        layer2[24][7:0] = buffer_data_2[4279:4272];
        layer2[24][15:8] = buffer_data_2[4287:4280];
        layer2[24][23:16] = buffer_data_2[4295:4288];
        layer2[24][31:24] = buffer_data_2[4303:4296];
        layer2[24][39:32] = buffer_data_2[4311:4304];
        layer3[24][7:0] = buffer_data_1[4279:4272];
        layer3[24][15:8] = buffer_data_1[4287:4280];
        layer3[24][23:16] = buffer_data_1[4295:4288];
        layer3[24][31:24] = buffer_data_1[4303:4296];
        layer3[24][39:32] = buffer_data_1[4311:4304];
        layer4[24][7:0] = buffer_data_0[4279:4272];
        layer4[24][15:8] = buffer_data_0[4287:4280];
        layer4[24][23:16] = buffer_data_0[4295:4288];
        layer4[24][31:24] = buffer_data_0[4303:4296];
        layer4[24][39:32] = buffer_data_0[4311:4304];
        layer0[25][7:0] = buffer_data_4[4287:4280];
        layer0[25][15:8] = buffer_data_4[4295:4288];
        layer0[25][23:16] = buffer_data_4[4303:4296];
        layer0[25][31:24] = buffer_data_4[4311:4304];
        layer0[25][39:32] = buffer_data_4[4319:4312];
        layer1[25][7:0] = buffer_data_3[4287:4280];
        layer1[25][15:8] = buffer_data_3[4295:4288];
        layer1[25][23:16] = buffer_data_3[4303:4296];
        layer1[25][31:24] = buffer_data_3[4311:4304];
        layer1[25][39:32] = buffer_data_3[4319:4312];
        layer2[25][7:0] = buffer_data_2[4287:4280];
        layer2[25][15:8] = buffer_data_2[4295:4288];
        layer2[25][23:16] = buffer_data_2[4303:4296];
        layer2[25][31:24] = buffer_data_2[4311:4304];
        layer2[25][39:32] = buffer_data_2[4319:4312];
        layer3[25][7:0] = buffer_data_1[4287:4280];
        layer3[25][15:8] = buffer_data_1[4295:4288];
        layer3[25][23:16] = buffer_data_1[4303:4296];
        layer3[25][31:24] = buffer_data_1[4311:4304];
        layer3[25][39:32] = buffer_data_1[4319:4312];
        layer4[25][7:0] = buffer_data_0[4287:4280];
        layer4[25][15:8] = buffer_data_0[4295:4288];
        layer4[25][23:16] = buffer_data_0[4303:4296];
        layer4[25][31:24] = buffer_data_0[4311:4304];
        layer4[25][39:32] = buffer_data_0[4319:4312];
        layer0[26][7:0] = buffer_data_4[4295:4288];
        layer0[26][15:8] = buffer_data_4[4303:4296];
        layer0[26][23:16] = buffer_data_4[4311:4304];
        layer0[26][31:24] = buffer_data_4[4319:4312];
        layer0[26][39:32] = buffer_data_4[4327:4320];
        layer1[26][7:0] = buffer_data_3[4295:4288];
        layer1[26][15:8] = buffer_data_3[4303:4296];
        layer1[26][23:16] = buffer_data_3[4311:4304];
        layer1[26][31:24] = buffer_data_3[4319:4312];
        layer1[26][39:32] = buffer_data_3[4327:4320];
        layer2[26][7:0] = buffer_data_2[4295:4288];
        layer2[26][15:8] = buffer_data_2[4303:4296];
        layer2[26][23:16] = buffer_data_2[4311:4304];
        layer2[26][31:24] = buffer_data_2[4319:4312];
        layer2[26][39:32] = buffer_data_2[4327:4320];
        layer3[26][7:0] = buffer_data_1[4295:4288];
        layer3[26][15:8] = buffer_data_1[4303:4296];
        layer3[26][23:16] = buffer_data_1[4311:4304];
        layer3[26][31:24] = buffer_data_1[4319:4312];
        layer3[26][39:32] = buffer_data_1[4327:4320];
        layer4[26][7:0] = buffer_data_0[4295:4288];
        layer4[26][15:8] = buffer_data_0[4303:4296];
        layer4[26][23:16] = buffer_data_0[4311:4304];
        layer4[26][31:24] = buffer_data_0[4319:4312];
        layer4[26][39:32] = buffer_data_0[4327:4320];
        layer0[27][7:0] = buffer_data_4[4303:4296];
        layer0[27][15:8] = buffer_data_4[4311:4304];
        layer0[27][23:16] = buffer_data_4[4319:4312];
        layer0[27][31:24] = buffer_data_4[4327:4320];
        layer0[27][39:32] = buffer_data_4[4335:4328];
        layer1[27][7:0] = buffer_data_3[4303:4296];
        layer1[27][15:8] = buffer_data_3[4311:4304];
        layer1[27][23:16] = buffer_data_3[4319:4312];
        layer1[27][31:24] = buffer_data_3[4327:4320];
        layer1[27][39:32] = buffer_data_3[4335:4328];
        layer2[27][7:0] = buffer_data_2[4303:4296];
        layer2[27][15:8] = buffer_data_2[4311:4304];
        layer2[27][23:16] = buffer_data_2[4319:4312];
        layer2[27][31:24] = buffer_data_2[4327:4320];
        layer2[27][39:32] = buffer_data_2[4335:4328];
        layer3[27][7:0] = buffer_data_1[4303:4296];
        layer3[27][15:8] = buffer_data_1[4311:4304];
        layer3[27][23:16] = buffer_data_1[4319:4312];
        layer3[27][31:24] = buffer_data_1[4327:4320];
        layer3[27][39:32] = buffer_data_1[4335:4328];
        layer4[27][7:0] = buffer_data_0[4303:4296];
        layer4[27][15:8] = buffer_data_0[4311:4304];
        layer4[27][23:16] = buffer_data_0[4319:4312];
        layer4[27][31:24] = buffer_data_0[4327:4320];
        layer4[27][39:32] = buffer_data_0[4335:4328];
        layer0[28][7:0] = buffer_data_4[4311:4304];
        layer0[28][15:8] = buffer_data_4[4319:4312];
        layer0[28][23:16] = buffer_data_4[4327:4320];
        layer0[28][31:24] = buffer_data_4[4335:4328];
        layer0[28][39:32] = buffer_data_4[4343:4336];
        layer1[28][7:0] = buffer_data_3[4311:4304];
        layer1[28][15:8] = buffer_data_3[4319:4312];
        layer1[28][23:16] = buffer_data_3[4327:4320];
        layer1[28][31:24] = buffer_data_3[4335:4328];
        layer1[28][39:32] = buffer_data_3[4343:4336];
        layer2[28][7:0] = buffer_data_2[4311:4304];
        layer2[28][15:8] = buffer_data_2[4319:4312];
        layer2[28][23:16] = buffer_data_2[4327:4320];
        layer2[28][31:24] = buffer_data_2[4335:4328];
        layer2[28][39:32] = buffer_data_2[4343:4336];
        layer3[28][7:0] = buffer_data_1[4311:4304];
        layer3[28][15:8] = buffer_data_1[4319:4312];
        layer3[28][23:16] = buffer_data_1[4327:4320];
        layer3[28][31:24] = buffer_data_1[4335:4328];
        layer3[28][39:32] = buffer_data_1[4343:4336];
        layer4[28][7:0] = buffer_data_0[4311:4304];
        layer4[28][15:8] = buffer_data_0[4319:4312];
        layer4[28][23:16] = buffer_data_0[4327:4320];
        layer4[28][31:24] = buffer_data_0[4335:4328];
        layer4[28][39:32] = buffer_data_0[4343:4336];
        layer0[29][7:0] = buffer_data_4[4319:4312];
        layer0[29][15:8] = buffer_data_4[4327:4320];
        layer0[29][23:16] = buffer_data_4[4335:4328];
        layer0[29][31:24] = buffer_data_4[4343:4336];
        layer0[29][39:32] = buffer_data_4[4351:4344];
        layer1[29][7:0] = buffer_data_3[4319:4312];
        layer1[29][15:8] = buffer_data_3[4327:4320];
        layer1[29][23:16] = buffer_data_3[4335:4328];
        layer1[29][31:24] = buffer_data_3[4343:4336];
        layer1[29][39:32] = buffer_data_3[4351:4344];
        layer2[29][7:0] = buffer_data_2[4319:4312];
        layer2[29][15:8] = buffer_data_2[4327:4320];
        layer2[29][23:16] = buffer_data_2[4335:4328];
        layer2[29][31:24] = buffer_data_2[4343:4336];
        layer2[29][39:32] = buffer_data_2[4351:4344];
        layer3[29][7:0] = buffer_data_1[4319:4312];
        layer3[29][15:8] = buffer_data_1[4327:4320];
        layer3[29][23:16] = buffer_data_1[4335:4328];
        layer3[29][31:24] = buffer_data_1[4343:4336];
        layer3[29][39:32] = buffer_data_1[4351:4344];
        layer4[29][7:0] = buffer_data_0[4319:4312];
        layer4[29][15:8] = buffer_data_0[4327:4320];
        layer4[29][23:16] = buffer_data_0[4335:4328];
        layer4[29][31:24] = buffer_data_0[4343:4336];
        layer4[29][39:32] = buffer_data_0[4351:4344];
        layer0[30][7:0] = buffer_data_4[4327:4320];
        layer0[30][15:8] = buffer_data_4[4335:4328];
        layer0[30][23:16] = buffer_data_4[4343:4336];
        layer0[30][31:24] = buffer_data_4[4351:4344];
        layer0[30][39:32] = buffer_data_4[4359:4352];
        layer1[30][7:0] = buffer_data_3[4327:4320];
        layer1[30][15:8] = buffer_data_3[4335:4328];
        layer1[30][23:16] = buffer_data_3[4343:4336];
        layer1[30][31:24] = buffer_data_3[4351:4344];
        layer1[30][39:32] = buffer_data_3[4359:4352];
        layer2[30][7:0] = buffer_data_2[4327:4320];
        layer2[30][15:8] = buffer_data_2[4335:4328];
        layer2[30][23:16] = buffer_data_2[4343:4336];
        layer2[30][31:24] = buffer_data_2[4351:4344];
        layer2[30][39:32] = buffer_data_2[4359:4352];
        layer3[30][7:0] = buffer_data_1[4327:4320];
        layer3[30][15:8] = buffer_data_1[4335:4328];
        layer3[30][23:16] = buffer_data_1[4343:4336];
        layer3[30][31:24] = buffer_data_1[4351:4344];
        layer3[30][39:32] = buffer_data_1[4359:4352];
        layer4[30][7:0] = buffer_data_0[4327:4320];
        layer4[30][15:8] = buffer_data_0[4335:4328];
        layer4[30][23:16] = buffer_data_0[4343:4336];
        layer4[30][31:24] = buffer_data_0[4351:4344];
        layer4[30][39:32] = buffer_data_0[4359:4352];
        layer0[31][7:0] = buffer_data_4[4335:4328];
        layer0[31][15:8] = buffer_data_4[4343:4336];
        layer0[31][23:16] = buffer_data_4[4351:4344];
        layer0[31][31:24] = buffer_data_4[4359:4352];
        layer0[31][39:32] = buffer_data_4[4367:4360];
        layer1[31][7:0] = buffer_data_3[4335:4328];
        layer1[31][15:8] = buffer_data_3[4343:4336];
        layer1[31][23:16] = buffer_data_3[4351:4344];
        layer1[31][31:24] = buffer_data_3[4359:4352];
        layer1[31][39:32] = buffer_data_3[4367:4360];
        layer2[31][7:0] = buffer_data_2[4335:4328];
        layer2[31][15:8] = buffer_data_2[4343:4336];
        layer2[31][23:16] = buffer_data_2[4351:4344];
        layer2[31][31:24] = buffer_data_2[4359:4352];
        layer2[31][39:32] = buffer_data_2[4367:4360];
        layer3[31][7:0] = buffer_data_1[4335:4328];
        layer3[31][15:8] = buffer_data_1[4343:4336];
        layer3[31][23:16] = buffer_data_1[4351:4344];
        layer3[31][31:24] = buffer_data_1[4359:4352];
        layer3[31][39:32] = buffer_data_1[4367:4360];
        layer4[31][7:0] = buffer_data_0[4335:4328];
        layer4[31][15:8] = buffer_data_0[4343:4336];
        layer4[31][23:16] = buffer_data_0[4351:4344];
        layer4[31][31:24] = buffer_data_0[4359:4352];
        layer4[31][39:32] = buffer_data_0[4367:4360];
        layer0[32][7:0] = buffer_data_4[4343:4336];
        layer0[32][15:8] = buffer_data_4[4351:4344];
        layer0[32][23:16] = buffer_data_4[4359:4352];
        layer0[32][31:24] = buffer_data_4[4367:4360];
        layer0[32][39:32] = buffer_data_4[4375:4368];
        layer1[32][7:0] = buffer_data_3[4343:4336];
        layer1[32][15:8] = buffer_data_3[4351:4344];
        layer1[32][23:16] = buffer_data_3[4359:4352];
        layer1[32][31:24] = buffer_data_3[4367:4360];
        layer1[32][39:32] = buffer_data_3[4375:4368];
        layer2[32][7:0] = buffer_data_2[4343:4336];
        layer2[32][15:8] = buffer_data_2[4351:4344];
        layer2[32][23:16] = buffer_data_2[4359:4352];
        layer2[32][31:24] = buffer_data_2[4367:4360];
        layer2[32][39:32] = buffer_data_2[4375:4368];
        layer3[32][7:0] = buffer_data_1[4343:4336];
        layer3[32][15:8] = buffer_data_1[4351:4344];
        layer3[32][23:16] = buffer_data_1[4359:4352];
        layer3[32][31:24] = buffer_data_1[4367:4360];
        layer3[32][39:32] = buffer_data_1[4375:4368];
        layer4[32][7:0] = buffer_data_0[4343:4336];
        layer4[32][15:8] = buffer_data_0[4351:4344];
        layer4[32][23:16] = buffer_data_0[4359:4352];
        layer4[32][31:24] = buffer_data_0[4367:4360];
        layer4[32][39:32] = buffer_data_0[4375:4368];
        layer0[33][7:0] = buffer_data_4[4351:4344];
        layer0[33][15:8] = buffer_data_4[4359:4352];
        layer0[33][23:16] = buffer_data_4[4367:4360];
        layer0[33][31:24] = buffer_data_4[4375:4368];
        layer0[33][39:32] = buffer_data_4[4383:4376];
        layer1[33][7:0] = buffer_data_3[4351:4344];
        layer1[33][15:8] = buffer_data_3[4359:4352];
        layer1[33][23:16] = buffer_data_3[4367:4360];
        layer1[33][31:24] = buffer_data_3[4375:4368];
        layer1[33][39:32] = buffer_data_3[4383:4376];
        layer2[33][7:0] = buffer_data_2[4351:4344];
        layer2[33][15:8] = buffer_data_2[4359:4352];
        layer2[33][23:16] = buffer_data_2[4367:4360];
        layer2[33][31:24] = buffer_data_2[4375:4368];
        layer2[33][39:32] = buffer_data_2[4383:4376];
        layer3[33][7:0] = buffer_data_1[4351:4344];
        layer3[33][15:8] = buffer_data_1[4359:4352];
        layer3[33][23:16] = buffer_data_1[4367:4360];
        layer3[33][31:24] = buffer_data_1[4375:4368];
        layer3[33][39:32] = buffer_data_1[4383:4376];
        layer4[33][7:0] = buffer_data_0[4351:4344];
        layer4[33][15:8] = buffer_data_0[4359:4352];
        layer4[33][23:16] = buffer_data_0[4367:4360];
        layer4[33][31:24] = buffer_data_0[4375:4368];
        layer4[33][39:32] = buffer_data_0[4383:4376];
        layer0[34][7:0] = buffer_data_4[4359:4352];
        layer0[34][15:8] = buffer_data_4[4367:4360];
        layer0[34][23:16] = buffer_data_4[4375:4368];
        layer0[34][31:24] = buffer_data_4[4383:4376];
        layer0[34][39:32] = buffer_data_4[4391:4384];
        layer1[34][7:0] = buffer_data_3[4359:4352];
        layer1[34][15:8] = buffer_data_3[4367:4360];
        layer1[34][23:16] = buffer_data_3[4375:4368];
        layer1[34][31:24] = buffer_data_3[4383:4376];
        layer1[34][39:32] = buffer_data_3[4391:4384];
        layer2[34][7:0] = buffer_data_2[4359:4352];
        layer2[34][15:8] = buffer_data_2[4367:4360];
        layer2[34][23:16] = buffer_data_2[4375:4368];
        layer2[34][31:24] = buffer_data_2[4383:4376];
        layer2[34][39:32] = buffer_data_2[4391:4384];
        layer3[34][7:0] = buffer_data_1[4359:4352];
        layer3[34][15:8] = buffer_data_1[4367:4360];
        layer3[34][23:16] = buffer_data_1[4375:4368];
        layer3[34][31:24] = buffer_data_1[4383:4376];
        layer3[34][39:32] = buffer_data_1[4391:4384];
        layer4[34][7:0] = buffer_data_0[4359:4352];
        layer4[34][15:8] = buffer_data_0[4367:4360];
        layer4[34][23:16] = buffer_data_0[4375:4368];
        layer4[34][31:24] = buffer_data_0[4383:4376];
        layer4[34][39:32] = buffer_data_0[4391:4384];
        layer0[35][7:0] = buffer_data_4[4367:4360];
        layer0[35][15:8] = buffer_data_4[4375:4368];
        layer0[35][23:16] = buffer_data_4[4383:4376];
        layer0[35][31:24] = buffer_data_4[4391:4384];
        layer0[35][39:32] = buffer_data_4[4399:4392];
        layer1[35][7:0] = buffer_data_3[4367:4360];
        layer1[35][15:8] = buffer_data_3[4375:4368];
        layer1[35][23:16] = buffer_data_3[4383:4376];
        layer1[35][31:24] = buffer_data_3[4391:4384];
        layer1[35][39:32] = buffer_data_3[4399:4392];
        layer2[35][7:0] = buffer_data_2[4367:4360];
        layer2[35][15:8] = buffer_data_2[4375:4368];
        layer2[35][23:16] = buffer_data_2[4383:4376];
        layer2[35][31:24] = buffer_data_2[4391:4384];
        layer2[35][39:32] = buffer_data_2[4399:4392];
        layer3[35][7:0] = buffer_data_1[4367:4360];
        layer3[35][15:8] = buffer_data_1[4375:4368];
        layer3[35][23:16] = buffer_data_1[4383:4376];
        layer3[35][31:24] = buffer_data_1[4391:4384];
        layer3[35][39:32] = buffer_data_1[4399:4392];
        layer4[35][7:0] = buffer_data_0[4367:4360];
        layer4[35][15:8] = buffer_data_0[4375:4368];
        layer4[35][23:16] = buffer_data_0[4383:4376];
        layer4[35][31:24] = buffer_data_0[4391:4384];
        layer4[35][39:32] = buffer_data_0[4399:4392];
        layer0[36][7:0] = buffer_data_4[4375:4368];
        layer0[36][15:8] = buffer_data_4[4383:4376];
        layer0[36][23:16] = buffer_data_4[4391:4384];
        layer0[36][31:24] = buffer_data_4[4399:4392];
        layer0[36][39:32] = buffer_data_4[4407:4400];
        layer1[36][7:0] = buffer_data_3[4375:4368];
        layer1[36][15:8] = buffer_data_3[4383:4376];
        layer1[36][23:16] = buffer_data_3[4391:4384];
        layer1[36][31:24] = buffer_data_3[4399:4392];
        layer1[36][39:32] = buffer_data_3[4407:4400];
        layer2[36][7:0] = buffer_data_2[4375:4368];
        layer2[36][15:8] = buffer_data_2[4383:4376];
        layer2[36][23:16] = buffer_data_2[4391:4384];
        layer2[36][31:24] = buffer_data_2[4399:4392];
        layer2[36][39:32] = buffer_data_2[4407:4400];
        layer3[36][7:0] = buffer_data_1[4375:4368];
        layer3[36][15:8] = buffer_data_1[4383:4376];
        layer3[36][23:16] = buffer_data_1[4391:4384];
        layer3[36][31:24] = buffer_data_1[4399:4392];
        layer3[36][39:32] = buffer_data_1[4407:4400];
        layer4[36][7:0] = buffer_data_0[4375:4368];
        layer4[36][15:8] = buffer_data_0[4383:4376];
        layer4[36][23:16] = buffer_data_0[4391:4384];
        layer4[36][31:24] = buffer_data_0[4399:4392];
        layer4[36][39:32] = buffer_data_0[4407:4400];
        layer0[37][7:0] = buffer_data_4[4383:4376];
        layer0[37][15:8] = buffer_data_4[4391:4384];
        layer0[37][23:16] = buffer_data_4[4399:4392];
        layer0[37][31:24] = buffer_data_4[4407:4400];
        layer0[37][39:32] = buffer_data_4[4415:4408];
        layer1[37][7:0] = buffer_data_3[4383:4376];
        layer1[37][15:8] = buffer_data_3[4391:4384];
        layer1[37][23:16] = buffer_data_3[4399:4392];
        layer1[37][31:24] = buffer_data_3[4407:4400];
        layer1[37][39:32] = buffer_data_3[4415:4408];
        layer2[37][7:0] = buffer_data_2[4383:4376];
        layer2[37][15:8] = buffer_data_2[4391:4384];
        layer2[37][23:16] = buffer_data_2[4399:4392];
        layer2[37][31:24] = buffer_data_2[4407:4400];
        layer2[37][39:32] = buffer_data_2[4415:4408];
        layer3[37][7:0] = buffer_data_1[4383:4376];
        layer3[37][15:8] = buffer_data_1[4391:4384];
        layer3[37][23:16] = buffer_data_1[4399:4392];
        layer3[37][31:24] = buffer_data_1[4407:4400];
        layer3[37][39:32] = buffer_data_1[4415:4408];
        layer4[37][7:0] = buffer_data_0[4383:4376];
        layer4[37][15:8] = buffer_data_0[4391:4384];
        layer4[37][23:16] = buffer_data_0[4399:4392];
        layer4[37][31:24] = buffer_data_0[4407:4400];
        layer4[37][39:32] = buffer_data_0[4415:4408];
        layer0[38][7:0] = buffer_data_4[4391:4384];
        layer0[38][15:8] = buffer_data_4[4399:4392];
        layer0[38][23:16] = buffer_data_4[4407:4400];
        layer0[38][31:24] = buffer_data_4[4415:4408];
        layer0[38][39:32] = buffer_data_4[4423:4416];
        layer1[38][7:0] = buffer_data_3[4391:4384];
        layer1[38][15:8] = buffer_data_3[4399:4392];
        layer1[38][23:16] = buffer_data_3[4407:4400];
        layer1[38][31:24] = buffer_data_3[4415:4408];
        layer1[38][39:32] = buffer_data_3[4423:4416];
        layer2[38][7:0] = buffer_data_2[4391:4384];
        layer2[38][15:8] = buffer_data_2[4399:4392];
        layer2[38][23:16] = buffer_data_2[4407:4400];
        layer2[38][31:24] = buffer_data_2[4415:4408];
        layer2[38][39:32] = buffer_data_2[4423:4416];
        layer3[38][7:0] = buffer_data_1[4391:4384];
        layer3[38][15:8] = buffer_data_1[4399:4392];
        layer3[38][23:16] = buffer_data_1[4407:4400];
        layer3[38][31:24] = buffer_data_1[4415:4408];
        layer3[38][39:32] = buffer_data_1[4423:4416];
        layer4[38][7:0] = buffer_data_0[4391:4384];
        layer4[38][15:8] = buffer_data_0[4399:4392];
        layer4[38][23:16] = buffer_data_0[4407:4400];
        layer4[38][31:24] = buffer_data_0[4415:4408];
        layer4[38][39:32] = buffer_data_0[4423:4416];
        layer0[39][7:0] = buffer_data_4[4399:4392];
        layer0[39][15:8] = buffer_data_4[4407:4400];
        layer0[39][23:16] = buffer_data_4[4415:4408];
        layer0[39][31:24] = buffer_data_4[4423:4416];
        layer0[39][39:32] = buffer_data_4[4431:4424];
        layer1[39][7:0] = buffer_data_3[4399:4392];
        layer1[39][15:8] = buffer_data_3[4407:4400];
        layer1[39][23:16] = buffer_data_3[4415:4408];
        layer1[39][31:24] = buffer_data_3[4423:4416];
        layer1[39][39:32] = buffer_data_3[4431:4424];
        layer2[39][7:0] = buffer_data_2[4399:4392];
        layer2[39][15:8] = buffer_data_2[4407:4400];
        layer2[39][23:16] = buffer_data_2[4415:4408];
        layer2[39][31:24] = buffer_data_2[4423:4416];
        layer2[39][39:32] = buffer_data_2[4431:4424];
        layer3[39][7:0] = buffer_data_1[4399:4392];
        layer3[39][15:8] = buffer_data_1[4407:4400];
        layer3[39][23:16] = buffer_data_1[4415:4408];
        layer3[39][31:24] = buffer_data_1[4423:4416];
        layer3[39][39:32] = buffer_data_1[4431:4424];
        layer4[39][7:0] = buffer_data_0[4399:4392];
        layer4[39][15:8] = buffer_data_0[4407:4400];
        layer4[39][23:16] = buffer_data_0[4415:4408];
        layer4[39][31:24] = buffer_data_0[4423:4416];
        layer4[39][39:32] = buffer_data_0[4431:4424];
        layer0[40][7:0] = buffer_data_4[4407:4400];
        layer0[40][15:8] = buffer_data_4[4415:4408];
        layer0[40][23:16] = buffer_data_4[4423:4416];
        layer0[40][31:24] = buffer_data_4[4431:4424];
        layer0[40][39:32] = buffer_data_4[4439:4432];
        layer1[40][7:0] = buffer_data_3[4407:4400];
        layer1[40][15:8] = buffer_data_3[4415:4408];
        layer1[40][23:16] = buffer_data_3[4423:4416];
        layer1[40][31:24] = buffer_data_3[4431:4424];
        layer1[40][39:32] = buffer_data_3[4439:4432];
        layer2[40][7:0] = buffer_data_2[4407:4400];
        layer2[40][15:8] = buffer_data_2[4415:4408];
        layer2[40][23:16] = buffer_data_2[4423:4416];
        layer2[40][31:24] = buffer_data_2[4431:4424];
        layer2[40][39:32] = buffer_data_2[4439:4432];
        layer3[40][7:0] = buffer_data_1[4407:4400];
        layer3[40][15:8] = buffer_data_1[4415:4408];
        layer3[40][23:16] = buffer_data_1[4423:4416];
        layer3[40][31:24] = buffer_data_1[4431:4424];
        layer3[40][39:32] = buffer_data_1[4439:4432];
        layer4[40][7:0] = buffer_data_0[4407:4400];
        layer4[40][15:8] = buffer_data_0[4415:4408];
        layer4[40][23:16] = buffer_data_0[4423:4416];
        layer4[40][31:24] = buffer_data_0[4431:4424];
        layer4[40][39:32] = buffer_data_0[4439:4432];
        layer0[41][7:0] = buffer_data_4[4415:4408];
        layer0[41][15:8] = buffer_data_4[4423:4416];
        layer0[41][23:16] = buffer_data_4[4431:4424];
        layer0[41][31:24] = buffer_data_4[4439:4432];
        layer0[41][39:32] = buffer_data_4[4447:4440];
        layer1[41][7:0] = buffer_data_3[4415:4408];
        layer1[41][15:8] = buffer_data_3[4423:4416];
        layer1[41][23:16] = buffer_data_3[4431:4424];
        layer1[41][31:24] = buffer_data_3[4439:4432];
        layer1[41][39:32] = buffer_data_3[4447:4440];
        layer2[41][7:0] = buffer_data_2[4415:4408];
        layer2[41][15:8] = buffer_data_2[4423:4416];
        layer2[41][23:16] = buffer_data_2[4431:4424];
        layer2[41][31:24] = buffer_data_2[4439:4432];
        layer2[41][39:32] = buffer_data_2[4447:4440];
        layer3[41][7:0] = buffer_data_1[4415:4408];
        layer3[41][15:8] = buffer_data_1[4423:4416];
        layer3[41][23:16] = buffer_data_1[4431:4424];
        layer3[41][31:24] = buffer_data_1[4439:4432];
        layer3[41][39:32] = buffer_data_1[4447:4440];
        layer4[41][7:0] = buffer_data_0[4415:4408];
        layer4[41][15:8] = buffer_data_0[4423:4416];
        layer4[41][23:16] = buffer_data_0[4431:4424];
        layer4[41][31:24] = buffer_data_0[4439:4432];
        layer4[41][39:32] = buffer_data_0[4447:4440];
        layer0[42][7:0] = buffer_data_4[4423:4416];
        layer0[42][15:8] = buffer_data_4[4431:4424];
        layer0[42][23:16] = buffer_data_4[4439:4432];
        layer0[42][31:24] = buffer_data_4[4447:4440];
        layer0[42][39:32] = buffer_data_4[4455:4448];
        layer1[42][7:0] = buffer_data_3[4423:4416];
        layer1[42][15:8] = buffer_data_3[4431:4424];
        layer1[42][23:16] = buffer_data_3[4439:4432];
        layer1[42][31:24] = buffer_data_3[4447:4440];
        layer1[42][39:32] = buffer_data_3[4455:4448];
        layer2[42][7:0] = buffer_data_2[4423:4416];
        layer2[42][15:8] = buffer_data_2[4431:4424];
        layer2[42][23:16] = buffer_data_2[4439:4432];
        layer2[42][31:24] = buffer_data_2[4447:4440];
        layer2[42][39:32] = buffer_data_2[4455:4448];
        layer3[42][7:0] = buffer_data_1[4423:4416];
        layer3[42][15:8] = buffer_data_1[4431:4424];
        layer3[42][23:16] = buffer_data_1[4439:4432];
        layer3[42][31:24] = buffer_data_1[4447:4440];
        layer3[42][39:32] = buffer_data_1[4455:4448];
        layer4[42][7:0] = buffer_data_0[4423:4416];
        layer4[42][15:8] = buffer_data_0[4431:4424];
        layer4[42][23:16] = buffer_data_0[4439:4432];
        layer4[42][31:24] = buffer_data_0[4447:4440];
        layer4[42][39:32] = buffer_data_0[4455:4448];
        layer0[43][7:0] = buffer_data_4[4431:4424];
        layer0[43][15:8] = buffer_data_4[4439:4432];
        layer0[43][23:16] = buffer_data_4[4447:4440];
        layer0[43][31:24] = buffer_data_4[4455:4448];
        layer0[43][39:32] = buffer_data_4[4463:4456];
        layer1[43][7:0] = buffer_data_3[4431:4424];
        layer1[43][15:8] = buffer_data_3[4439:4432];
        layer1[43][23:16] = buffer_data_3[4447:4440];
        layer1[43][31:24] = buffer_data_3[4455:4448];
        layer1[43][39:32] = buffer_data_3[4463:4456];
        layer2[43][7:0] = buffer_data_2[4431:4424];
        layer2[43][15:8] = buffer_data_2[4439:4432];
        layer2[43][23:16] = buffer_data_2[4447:4440];
        layer2[43][31:24] = buffer_data_2[4455:4448];
        layer2[43][39:32] = buffer_data_2[4463:4456];
        layer3[43][7:0] = buffer_data_1[4431:4424];
        layer3[43][15:8] = buffer_data_1[4439:4432];
        layer3[43][23:16] = buffer_data_1[4447:4440];
        layer3[43][31:24] = buffer_data_1[4455:4448];
        layer3[43][39:32] = buffer_data_1[4463:4456];
        layer4[43][7:0] = buffer_data_0[4431:4424];
        layer4[43][15:8] = buffer_data_0[4439:4432];
        layer4[43][23:16] = buffer_data_0[4447:4440];
        layer4[43][31:24] = buffer_data_0[4455:4448];
        layer4[43][39:32] = buffer_data_0[4463:4456];
        layer0[44][7:0] = buffer_data_4[4439:4432];
        layer0[44][15:8] = buffer_data_4[4447:4440];
        layer0[44][23:16] = buffer_data_4[4455:4448];
        layer0[44][31:24] = buffer_data_4[4463:4456];
        layer0[44][39:32] = buffer_data_4[4471:4464];
        layer1[44][7:0] = buffer_data_3[4439:4432];
        layer1[44][15:8] = buffer_data_3[4447:4440];
        layer1[44][23:16] = buffer_data_3[4455:4448];
        layer1[44][31:24] = buffer_data_3[4463:4456];
        layer1[44][39:32] = buffer_data_3[4471:4464];
        layer2[44][7:0] = buffer_data_2[4439:4432];
        layer2[44][15:8] = buffer_data_2[4447:4440];
        layer2[44][23:16] = buffer_data_2[4455:4448];
        layer2[44][31:24] = buffer_data_2[4463:4456];
        layer2[44][39:32] = buffer_data_2[4471:4464];
        layer3[44][7:0] = buffer_data_1[4439:4432];
        layer3[44][15:8] = buffer_data_1[4447:4440];
        layer3[44][23:16] = buffer_data_1[4455:4448];
        layer3[44][31:24] = buffer_data_1[4463:4456];
        layer3[44][39:32] = buffer_data_1[4471:4464];
        layer4[44][7:0] = buffer_data_0[4439:4432];
        layer4[44][15:8] = buffer_data_0[4447:4440];
        layer4[44][23:16] = buffer_data_0[4455:4448];
        layer4[44][31:24] = buffer_data_0[4463:4456];
        layer4[44][39:32] = buffer_data_0[4471:4464];
        layer0[45][7:0] = buffer_data_4[4447:4440];
        layer0[45][15:8] = buffer_data_4[4455:4448];
        layer0[45][23:16] = buffer_data_4[4463:4456];
        layer0[45][31:24] = buffer_data_4[4471:4464];
        layer0[45][39:32] = buffer_data_4[4479:4472];
        layer1[45][7:0] = buffer_data_3[4447:4440];
        layer1[45][15:8] = buffer_data_3[4455:4448];
        layer1[45][23:16] = buffer_data_3[4463:4456];
        layer1[45][31:24] = buffer_data_3[4471:4464];
        layer1[45][39:32] = buffer_data_3[4479:4472];
        layer2[45][7:0] = buffer_data_2[4447:4440];
        layer2[45][15:8] = buffer_data_2[4455:4448];
        layer2[45][23:16] = buffer_data_2[4463:4456];
        layer2[45][31:24] = buffer_data_2[4471:4464];
        layer2[45][39:32] = buffer_data_2[4479:4472];
        layer3[45][7:0] = buffer_data_1[4447:4440];
        layer3[45][15:8] = buffer_data_1[4455:4448];
        layer3[45][23:16] = buffer_data_1[4463:4456];
        layer3[45][31:24] = buffer_data_1[4471:4464];
        layer3[45][39:32] = buffer_data_1[4479:4472];
        layer4[45][7:0] = buffer_data_0[4447:4440];
        layer4[45][15:8] = buffer_data_0[4455:4448];
        layer4[45][23:16] = buffer_data_0[4463:4456];
        layer4[45][31:24] = buffer_data_0[4471:4464];
        layer4[45][39:32] = buffer_data_0[4479:4472];
        layer0[46][7:0] = buffer_data_4[4455:4448];
        layer0[46][15:8] = buffer_data_4[4463:4456];
        layer0[46][23:16] = buffer_data_4[4471:4464];
        layer0[46][31:24] = buffer_data_4[4479:4472];
        layer0[46][39:32] = buffer_data_4[4487:4480];
        layer1[46][7:0] = buffer_data_3[4455:4448];
        layer1[46][15:8] = buffer_data_3[4463:4456];
        layer1[46][23:16] = buffer_data_3[4471:4464];
        layer1[46][31:24] = buffer_data_3[4479:4472];
        layer1[46][39:32] = buffer_data_3[4487:4480];
        layer2[46][7:0] = buffer_data_2[4455:4448];
        layer2[46][15:8] = buffer_data_2[4463:4456];
        layer2[46][23:16] = buffer_data_2[4471:4464];
        layer2[46][31:24] = buffer_data_2[4479:4472];
        layer2[46][39:32] = buffer_data_2[4487:4480];
        layer3[46][7:0] = buffer_data_1[4455:4448];
        layer3[46][15:8] = buffer_data_1[4463:4456];
        layer3[46][23:16] = buffer_data_1[4471:4464];
        layer3[46][31:24] = buffer_data_1[4479:4472];
        layer3[46][39:32] = buffer_data_1[4487:4480];
        layer4[46][7:0] = buffer_data_0[4455:4448];
        layer4[46][15:8] = buffer_data_0[4463:4456];
        layer4[46][23:16] = buffer_data_0[4471:4464];
        layer4[46][31:24] = buffer_data_0[4479:4472];
        layer4[46][39:32] = buffer_data_0[4487:4480];
        layer0[47][7:0] = buffer_data_4[4463:4456];
        layer0[47][15:8] = buffer_data_4[4471:4464];
        layer0[47][23:16] = buffer_data_4[4479:4472];
        layer0[47][31:24] = buffer_data_4[4487:4480];
        layer0[47][39:32] = buffer_data_4[4495:4488];
        layer1[47][7:0] = buffer_data_3[4463:4456];
        layer1[47][15:8] = buffer_data_3[4471:4464];
        layer1[47][23:16] = buffer_data_3[4479:4472];
        layer1[47][31:24] = buffer_data_3[4487:4480];
        layer1[47][39:32] = buffer_data_3[4495:4488];
        layer2[47][7:0] = buffer_data_2[4463:4456];
        layer2[47][15:8] = buffer_data_2[4471:4464];
        layer2[47][23:16] = buffer_data_2[4479:4472];
        layer2[47][31:24] = buffer_data_2[4487:4480];
        layer2[47][39:32] = buffer_data_2[4495:4488];
        layer3[47][7:0] = buffer_data_1[4463:4456];
        layer3[47][15:8] = buffer_data_1[4471:4464];
        layer3[47][23:16] = buffer_data_1[4479:4472];
        layer3[47][31:24] = buffer_data_1[4487:4480];
        layer3[47][39:32] = buffer_data_1[4495:4488];
        layer4[47][7:0] = buffer_data_0[4463:4456];
        layer4[47][15:8] = buffer_data_0[4471:4464];
        layer4[47][23:16] = buffer_data_0[4479:4472];
        layer4[47][31:24] = buffer_data_0[4487:4480];
        layer4[47][39:32] = buffer_data_0[4495:4488];
        layer0[48][7:0] = buffer_data_4[4471:4464];
        layer0[48][15:8] = buffer_data_4[4479:4472];
        layer0[48][23:16] = buffer_data_4[4487:4480];
        layer0[48][31:24] = buffer_data_4[4495:4488];
        layer0[48][39:32] = buffer_data_4[4503:4496];
        layer1[48][7:0] = buffer_data_3[4471:4464];
        layer1[48][15:8] = buffer_data_3[4479:4472];
        layer1[48][23:16] = buffer_data_3[4487:4480];
        layer1[48][31:24] = buffer_data_3[4495:4488];
        layer1[48][39:32] = buffer_data_3[4503:4496];
        layer2[48][7:0] = buffer_data_2[4471:4464];
        layer2[48][15:8] = buffer_data_2[4479:4472];
        layer2[48][23:16] = buffer_data_2[4487:4480];
        layer2[48][31:24] = buffer_data_2[4495:4488];
        layer2[48][39:32] = buffer_data_2[4503:4496];
        layer3[48][7:0] = buffer_data_1[4471:4464];
        layer3[48][15:8] = buffer_data_1[4479:4472];
        layer3[48][23:16] = buffer_data_1[4487:4480];
        layer3[48][31:24] = buffer_data_1[4495:4488];
        layer3[48][39:32] = buffer_data_1[4503:4496];
        layer4[48][7:0] = buffer_data_0[4471:4464];
        layer4[48][15:8] = buffer_data_0[4479:4472];
        layer4[48][23:16] = buffer_data_0[4487:4480];
        layer4[48][31:24] = buffer_data_0[4495:4488];
        layer4[48][39:32] = buffer_data_0[4503:4496];
        layer0[49][7:0] = buffer_data_4[4479:4472];
        layer0[49][15:8] = buffer_data_4[4487:4480];
        layer0[49][23:16] = buffer_data_4[4495:4488];
        layer0[49][31:24] = buffer_data_4[4503:4496];
        layer0[49][39:32] = buffer_data_4[4511:4504];
        layer1[49][7:0] = buffer_data_3[4479:4472];
        layer1[49][15:8] = buffer_data_3[4487:4480];
        layer1[49][23:16] = buffer_data_3[4495:4488];
        layer1[49][31:24] = buffer_data_3[4503:4496];
        layer1[49][39:32] = buffer_data_3[4511:4504];
        layer2[49][7:0] = buffer_data_2[4479:4472];
        layer2[49][15:8] = buffer_data_2[4487:4480];
        layer2[49][23:16] = buffer_data_2[4495:4488];
        layer2[49][31:24] = buffer_data_2[4503:4496];
        layer2[49][39:32] = buffer_data_2[4511:4504];
        layer3[49][7:0] = buffer_data_1[4479:4472];
        layer3[49][15:8] = buffer_data_1[4487:4480];
        layer3[49][23:16] = buffer_data_1[4495:4488];
        layer3[49][31:24] = buffer_data_1[4503:4496];
        layer3[49][39:32] = buffer_data_1[4511:4504];
        layer4[49][7:0] = buffer_data_0[4479:4472];
        layer4[49][15:8] = buffer_data_0[4487:4480];
        layer4[49][23:16] = buffer_data_0[4495:4488];
        layer4[49][31:24] = buffer_data_0[4503:4496];
        layer4[49][39:32] = buffer_data_0[4511:4504];
        layer0[50][7:0] = buffer_data_4[4487:4480];
        layer0[50][15:8] = buffer_data_4[4495:4488];
        layer0[50][23:16] = buffer_data_4[4503:4496];
        layer0[50][31:24] = buffer_data_4[4511:4504];
        layer0[50][39:32] = buffer_data_4[4519:4512];
        layer1[50][7:0] = buffer_data_3[4487:4480];
        layer1[50][15:8] = buffer_data_3[4495:4488];
        layer1[50][23:16] = buffer_data_3[4503:4496];
        layer1[50][31:24] = buffer_data_3[4511:4504];
        layer1[50][39:32] = buffer_data_3[4519:4512];
        layer2[50][7:0] = buffer_data_2[4487:4480];
        layer2[50][15:8] = buffer_data_2[4495:4488];
        layer2[50][23:16] = buffer_data_2[4503:4496];
        layer2[50][31:24] = buffer_data_2[4511:4504];
        layer2[50][39:32] = buffer_data_2[4519:4512];
        layer3[50][7:0] = buffer_data_1[4487:4480];
        layer3[50][15:8] = buffer_data_1[4495:4488];
        layer3[50][23:16] = buffer_data_1[4503:4496];
        layer3[50][31:24] = buffer_data_1[4511:4504];
        layer3[50][39:32] = buffer_data_1[4519:4512];
        layer4[50][7:0] = buffer_data_0[4487:4480];
        layer4[50][15:8] = buffer_data_0[4495:4488];
        layer4[50][23:16] = buffer_data_0[4503:4496];
        layer4[50][31:24] = buffer_data_0[4511:4504];
        layer4[50][39:32] = buffer_data_0[4519:4512];
        layer0[51][7:0] = buffer_data_4[4495:4488];
        layer0[51][15:8] = buffer_data_4[4503:4496];
        layer0[51][23:16] = buffer_data_4[4511:4504];
        layer0[51][31:24] = buffer_data_4[4519:4512];
        layer0[51][39:32] = buffer_data_4[4527:4520];
        layer1[51][7:0] = buffer_data_3[4495:4488];
        layer1[51][15:8] = buffer_data_3[4503:4496];
        layer1[51][23:16] = buffer_data_3[4511:4504];
        layer1[51][31:24] = buffer_data_3[4519:4512];
        layer1[51][39:32] = buffer_data_3[4527:4520];
        layer2[51][7:0] = buffer_data_2[4495:4488];
        layer2[51][15:8] = buffer_data_2[4503:4496];
        layer2[51][23:16] = buffer_data_2[4511:4504];
        layer2[51][31:24] = buffer_data_2[4519:4512];
        layer2[51][39:32] = buffer_data_2[4527:4520];
        layer3[51][7:0] = buffer_data_1[4495:4488];
        layer3[51][15:8] = buffer_data_1[4503:4496];
        layer3[51][23:16] = buffer_data_1[4511:4504];
        layer3[51][31:24] = buffer_data_1[4519:4512];
        layer3[51][39:32] = buffer_data_1[4527:4520];
        layer4[51][7:0] = buffer_data_0[4495:4488];
        layer4[51][15:8] = buffer_data_0[4503:4496];
        layer4[51][23:16] = buffer_data_0[4511:4504];
        layer4[51][31:24] = buffer_data_0[4519:4512];
        layer4[51][39:32] = buffer_data_0[4527:4520];
        layer0[52][7:0] = buffer_data_4[4503:4496];
        layer0[52][15:8] = buffer_data_4[4511:4504];
        layer0[52][23:16] = buffer_data_4[4519:4512];
        layer0[52][31:24] = buffer_data_4[4527:4520];
        layer0[52][39:32] = buffer_data_4[4535:4528];
        layer1[52][7:0] = buffer_data_3[4503:4496];
        layer1[52][15:8] = buffer_data_3[4511:4504];
        layer1[52][23:16] = buffer_data_3[4519:4512];
        layer1[52][31:24] = buffer_data_3[4527:4520];
        layer1[52][39:32] = buffer_data_3[4535:4528];
        layer2[52][7:0] = buffer_data_2[4503:4496];
        layer2[52][15:8] = buffer_data_2[4511:4504];
        layer2[52][23:16] = buffer_data_2[4519:4512];
        layer2[52][31:24] = buffer_data_2[4527:4520];
        layer2[52][39:32] = buffer_data_2[4535:4528];
        layer3[52][7:0] = buffer_data_1[4503:4496];
        layer3[52][15:8] = buffer_data_1[4511:4504];
        layer3[52][23:16] = buffer_data_1[4519:4512];
        layer3[52][31:24] = buffer_data_1[4527:4520];
        layer3[52][39:32] = buffer_data_1[4535:4528];
        layer4[52][7:0] = buffer_data_0[4503:4496];
        layer4[52][15:8] = buffer_data_0[4511:4504];
        layer4[52][23:16] = buffer_data_0[4519:4512];
        layer4[52][31:24] = buffer_data_0[4527:4520];
        layer4[52][39:32] = buffer_data_0[4535:4528];
        layer0[53][7:0] = buffer_data_4[4511:4504];
        layer0[53][15:8] = buffer_data_4[4519:4512];
        layer0[53][23:16] = buffer_data_4[4527:4520];
        layer0[53][31:24] = buffer_data_4[4535:4528];
        layer0[53][39:32] = buffer_data_4[4543:4536];
        layer1[53][7:0] = buffer_data_3[4511:4504];
        layer1[53][15:8] = buffer_data_3[4519:4512];
        layer1[53][23:16] = buffer_data_3[4527:4520];
        layer1[53][31:24] = buffer_data_3[4535:4528];
        layer1[53][39:32] = buffer_data_3[4543:4536];
        layer2[53][7:0] = buffer_data_2[4511:4504];
        layer2[53][15:8] = buffer_data_2[4519:4512];
        layer2[53][23:16] = buffer_data_2[4527:4520];
        layer2[53][31:24] = buffer_data_2[4535:4528];
        layer2[53][39:32] = buffer_data_2[4543:4536];
        layer3[53][7:0] = buffer_data_1[4511:4504];
        layer3[53][15:8] = buffer_data_1[4519:4512];
        layer3[53][23:16] = buffer_data_1[4527:4520];
        layer3[53][31:24] = buffer_data_1[4535:4528];
        layer3[53][39:32] = buffer_data_1[4543:4536];
        layer4[53][7:0] = buffer_data_0[4511:4504];
        layer4[53][15:8] = buffer_data_0[4519:4512];
        layer4[53][23:16] = buffer_data_0[4527:4520];
        layer4[53][31:24] = buffer_data_0[4535:4528];
        layer4[53][39:32] = buffer_data_0[4543:4536];
        layer0[54][7:0] = buffer_data_4[4519:4512];
        layer0[54][15:8] = buffer_data_4[4527:4520];
        layer0[54][23:16] = buffer_data_4[4535:4528];
        layer0[54][31:24] = buffer_data_4[4543:4536];
        layer0[54][39:32] = buffer_data_4[4551:4544];
        layer1[54][7:0] = buffer_data_3[4519:4512];
        layer1[54][15:8] = buffer_data_3[4527:4520];
        layer1[54][23:16] = buffer_data_3[4535:4528];
        layer1[54][31:24] = buffer_data_3[4543:4536];
        layer1[54][39:32] = buffer_data_3[4551:4544];
        layer2[54][7:0] = buffer_data_2[4519:4512];
        layer2[54][15:8] = buffer_data_2[4527:4520];
        layer2[54][23:16] = buffer_data_2[4535:4528];
        layer2[54][31:24] = buffer_data_2[4543:4536];
        layer2[54][39:32] = buffer_data_2[4551:4544];
        layer3[54][7:0] = buffer_data_1[4519:4512];
        layer3[54][15:8] = buffer_data_1[4527:4520];
        layer3[54][23:16] = buffer_data_1[4535:4528];
        layer3[54][31:24] = buffer_data_1[4543:4536];
        layer3[54][39:32] = buffer_data_1[4551:4544];
        layer4[54][7:0] = buffer_data_0[4519:4512];
        layer4[54][15:8] = buffer_data_0[4527:4520];
        layer4[54][23:16] = buffer_data_0[4535:4528];
        layer4[54][31:24] = buffer_data_0[4543:4536];
        layer4[54][39:32] = buffer_data_0[4551:4544];
        layer0[55][7:0] = buffer_data_4[4527:4520];
        layer0[55][15:8] = buffer_data_4[4535:4528];
        layer0[55][23:16] = buffer_data_4[4543:4536];
        layer0[55][31:24] = buffer_data_4[4551:4544];
        layer0[55][39:32] = buffer_data_4[4559:4552];
        layer1[55][7:0] = buffer_data_3[4527:4520];
        layer1[55][15:8] = buffer_data_3[4535:4528];
        layer1[55][23:16] = buffer_data_3[4543:4536];
        layer1[55][31:24] = buffer_data_3[4551:4544];
        layer1[55][39:32] = buffer_data_3[4559:4552];
        layer2[55][7:0] = buffer_data_2[4527:4520];
        layer2[55][15:8] = buffer_data_2[4535:4528];
        layer2[55][23:16] = buffer_data_2[4543:4536];
        layer2[55][31:24] = buffer_data_2[4551:4544];
        layer2[55][39:32] = buffer_data_2[4559:4552];
        layer3[55][7:0] = buffer_data_1[4527:4520];
        layer3[55][15:8] = buffer_data_1[4535:4528];
        layer3[55][23:16] = buffer_data_1[4543:4536];
        layer3[55][31:24] = buffer_data_1[4551:4544];
        layer3[55][39:32] = buffer_data_1[4559:4552];
        layer4[55][7:0] = buffer_data_0[4527:4520];
        layer4[55][15:8] = buffer_data_0[4535:4528];
        layer4[55][23:16] = buffer_data_0[4543:4536];
        layer4[55][31:24] = buffer_data_0[4551:4544];
        layer4[55][39:32] = buffer_data_0[4559:4552];
        layer0[56][7:0] = buffer_data_4[4535:4528];
        layer0[56][15:8] = buffer_data_4[4543:4536];
        layer0[56][23:16] = buffer_data_4[4551:4544];
        layer0[56][31:24] = buffer_data_4[4559:4552];
        layer0[56][39:32] = buffer_data_4[4567:4560];
        layer1[56][7:0] = buffer_data_3[4535:4528];
        layer1[56][15:8] = buffer_data_3[4543:4536];
        layer1[56][23:16] = buffer_data_3[4551:4544];
        layer1[56][31:24] = buffer_data_3[4559:4552];
        layer1[56][39:32] = buffer_data_3[4567:4560];
        layer2[56][7:0] = buffer_data_2[4535:4528];
        layer2[56][15:8] = buffer_data_2[4543:4536];
        layer2[56][23:16] = buffer_data_2[4551:4544];
        layer2[56][31:24] = buffer_data_2[4559:4552];
        layer2[56][39:32] = buffer_data_2[4567:4560];
        layer3[56][7:0] = buffer_data_1[4535:4528];
        layer3[56][15:8] = buffer_data_1[4543:4536];
        layer3[56][23:16] = buffer_data_1[4551:4544];
        layer3[56][31:24] = buffer_data_1[4559:4552];
        layer3[56][39:32] = buffer_data_1[4567:4560];
        layer4[56][7:0] = buffer_data_0[4535:4528];
        layer4[56][15:8] = buffer_data_0[4543:4536];
        layer4[56][23:16] = buffer_data_0[4551:4544];
        layer4[56][31:24] = buffer_data_0[4559:4552];
        layer4[56][39:32] = buffer_data_0[4567:4560];
        layer0[57][7:0] = buffer_data_4[4543:4536];
        layer0[57][15:8] = buffer_data_4[4551:4544];
        layer0[57][23:16] = buffer_data_4[4559:4552];
        layer0[57][31:24] = buffer_data_4[4567:4560];
        layer0[57][39:32] = buffer_data_4[4575:4568];
        layer1[57][7:0] = buffer_data_3[4543:4536];
        layer1[57][15:8] = buffer_data_3[4551:4544];
        layer1[57][23:16] = buffer_data_3[4559:4552];
        layer1[57][31:24] = buffer_data_3[4567:4560];
        layer1[57][39:32] = buffer_data_3[4575:4568];
        layer2[57][7:0] = buffer_data_2[4543:4536];
        layer2[57][15:8] = buffer_data_2[4551:4544];
        layer2[57][23:16] = buffer_data_2[4559:4552];
        layer2[57][31:24] = buffer_data_2[4567:4560];
        layer2[57][39:32] = buffer_data_2[4575:4568];
        layer3[57][7:0] = buffer_data_1[4543:4536];
        layer3[57][15:8] = buffer_data_1[4551:4544];
        layer3[57][23:16] = buffer_data_1[4559:4552];
        layer3[57][31:24] = buffer_data_1[4567:4560];
        layer3[57][39:32] = buffer_data_1[4575:4568];
        layer4[57][7:0] = buffer_data_0[4543:4536];
        layer4[57][15:8] = buffer_data_0[4551:4544];
        layer4[57][23:16] = buffer_data_0[4559:4552];
        layer4[57][31:24] = buffer_data_0[4567:4560];
        layer4[57][39:32] = buffer_data_0[4575:4568];
        layer0[58][7:0] = buffer_data_4[4551:4544];
        layer0[58][15:8] = buffer_data_4[4559:4552];
        layer0[58][23:16] = buffer_data_4[4567:4560];
        layer0[58][31:24] = buffer_data_4[4575:4568];
        layer0[58][39:32] = buffer_data_4[4583:4576];
        layer1[58][7:0] = buffer_data_3[4551:4544];
        layer1[58][15:8] = buffer_data_3[4559:4552];
        layer1[58][23:16] = buffer_data_3[4567:4560];
        layer1[58][31:24] = buffer_data_3[4575:4568];
        layer1[58][39:32] = buffer_data_3[4583:4576];
        layer2[58][7:0] = buffer_data_2[4551:4544];
        layer2[58][15:8] = buffer_data_2[4559:4552];
        layer2[58][23:16] = buffer_data_2[4567:4560];
        layer2[58][31:24] = buffer_data_2[4575:4568];
        layer2[58][39:32] = buffer_data_2[4583:4576];
        layer3[58][7:0] = buffer_data_1[4551:4544];
        layer3[58][15:8] = buffer_data_1[4559:4552];
        layer3[58][23:16] = buffer_data_1[4567:4560];
        layer3[58][31:24] = buffer_data_1[4575:4568];
        layer3[58][39:32] = buffer_data_1[4583:4576];
        layer4[58][7:0] = buffer_data_0[4551:4544];
        layer4[58][15:8] = buffer_data_0[4559:4552];
        layer4[58][23:16] = buffer_data_0[4567:4560];
        layer4[58][31:24] = buffer_data_0[4575:4568];
        layer4[58][39:32] = buffer_data_0[4583:4576];
        layer0[59][7:0] = buffer_data_4[4559:4552];
        layer0[59][15:8] = buffer_data_4[4567:4560];
        layer0[59][23:16] = buffer_data_4[4575:4568];
        layer0[59][31:24] = buffer_data_4[4583:4576];
        layer0[59][39:32] = buffer_data_4[4591:4584];
        layer1[59][7:0] = buffer_data_3[4559:4552];
        layer1[59][15:8] = buffer_data_3[4567:4560];
        layer1[59][23:16] = buffer_data_3[4575:4568];
        layer1[59][31:24] = buffer_data_3[4583:4576];
        layer1[59][39:32] = buffer_data_3[4591:4584];
        layer2[59][7:0] = buffer_data_2[4559:4552];
        layer2[59][15:8] = buffer_data_2[4567:4560];
        layer2[59][23:16] = buffer_data_2[4575:4568];
        layer2[59][31:24] = buffer_data_2[4583:4576];
        layer2[59][39:32] = buffer_data_2[4591:4584];
        layer3[59][7:0] = buffer_data_1[4559:4552];
        layer3[59][15:8] = buffer_data_1[4567:4560];
        layer3[59][23:16] = buffer_data_1[4575:4568];
        layer3[59][31:24] = buffer_data_1[4583:4576];
        layer3[59][39:32] = buffer_data_1[4591:4584];
        layer4[59][7:0] = buffer_data_0[4559:4552];
        layer4[59][15:8] = buffer_data_0[4567:4560];
        layer4[59][23:16] = buffer_data_0[4575:4568];
        layer4[59][31:24] = buffer_data_0[4583:4576];
        layer4[59][39:32] = buffer_data_0[4591:4584];
        layer0[60][7:0] = buffer_data_4[4567:4560];
        layer0[60][15:8] = buffer_data_4[4575:4568];
        layer0[60][23:16] = buffer_data_4[4583:4576];
        layer0[60][31:24] = buffer_data_4[4591:4584];
        layer0[60][39:32] = buffer_data_4[4599:4592];
        layer1[60][7:0] = buffer_data_3[4567:4560];
        layer1[60][15:8] = buffer_data_3[4575:4568];
        layer1[60][23:16] = buffer_data_3[4583:4576];
        layer1[60][31:24] = buffer_data_3[4591:4584];
        layer1[60][39:32] = buffer_data_3[4599:4592];
        layer2[60][7:0] = buffer_data_2[4567:4560];
        layer2[60][15:8] = buffer_data_2[4575:4568];
        layer2[60][23:16] = buffer_data_2[4583:4576];
        layer2[60][31:24] = buffer_data_2[4591:4584];
        layer2[60][39:32] = buffer_data_2[4599:4592];
        layer3[60][7:0] = buffer_data_1[4567:4560];
        layer3[60][15:8] = buffer_data_1[4575:4568];
        layer3[60][23:16] = buffer_data_1[4583:4576];
        layer3[60][31:24] = buffer_data_1[4591:4584];
        layer3[60][39:32] = buffer_data_1[4599:4592];
        layer4[60][7:0] = buffer_data_0[4567:4560];
        layer4[60][15:8] = buffer_data_0[4575:4568];
        layer4[60][23:16] = buffer_data_0[4583:4576];
        layer4[60][31:24] = buffer_data_0[4591:4584];
        layer4[60][39:32] = buffer_data_0[4599:4592];
        layer0[61][7:0] = buffer_data_4[4575:4568];
        layer0[61][15:8] = buffer_data_4[4583:4576];
        layer0[61][23:16] = buffer_data_4[4591:4584];
        layer0[61][31:24] = buffer_data_4[4599:4592];
        layer0[61][39:32] = buffer_data_4[4607:4600];
        layer1[61][7:0] = buffer_data_3[4575:4568];
        layer1[61][15:8] = buffer_data_3[4583:4576];
        layer1[61][23:16] = buffer_data_3[4591:4584];
        layer1[61][31:24] = buffer_data_3[4599:4592];
        layer1[61][39:32] = buffer_data_3[4607:4600];
        layer2[61][7:0] = buffer_data_2[4575:4568];
        layer2[61][15:8] = buffer_data_2[4583:4576];
        layer2[61][23:16] = buffer_data_2[4591:4584];
        layer2[61][31:24] = buffer_data_2[4599:4592];
        layer2[61][39:32] = buffer_data_2[4607:4600];
        layer3[61][7:0] = buffer_data_1[4575:4568];
        layer3[61][15:8] = buffer_data_1[4583:4576];
        layer3[61][23:16] = buffer_data_1[4591:4584];
        layer3[61][31:24] = buffer_data_1[4599:4592];
        layer3[61][39:32] = buffer_data_1[4607:4600];
        layer4[61][7:0] = buffer_data_0[4575:4568];
        layer4[61][15:8] = buffer_data_0[4583:4576];
        layer4[61][23:16] = buffer_data_0[4591:4584];
        layer4[61][31:24] = buffer_data_0[4599:4592];
        layer4[61][39:32] = buffer_data_0[4607:4600];
        layer0[62][7:0] = buffer_data_4[4583:4576];
        layer0[62][15:8] = buffer_data_4[4591:4584];
        layer0[62][23:16] = buffer_data_4[4599:4592];
        layer0[62][31:24] = buffer_data_4[4607:4600];
        layer0[62][39:32] = buffer_data_4[4615:4608];
        layer1[62][7:0] = buffer_data_3[4583:4576];
        layer1[62][15:8] = buffer_data_3[4591:4584];
        layer1[62][23:16] = buffer_data_3[4599:4592];
        layer1[62][31:24] = buffer_data_3[4607:4600];
        layer1[62][39:32] = buffer_data_3[4615:4608];
        layer2[62][7:0] = buffer_data_2[4583:4576];
        layer2[62][15:8] = buffer_data_2[4591:4584];
        layer2[62][23:16] = buffer_data_2[4599:4592];
        layer2[62][31:24] = buffer_data_2[4607:4600];
        layer2[62][39:32] = buffer_data_2[4615:4608];
        layer3[62][7:0] = buffer_data_1[4583:4576];
        layer3[62][15:8] = buffer_data_1[4591:4584];
        layer3[62][23:16] = buffer_data_1[4599:4592];
        layer3[62][31:24] = buffer_data_1[4607:4600];
        layer3[62][39:32] = buffer_data_1[4615:4608];
        layer4[62][7:0] = buffer_data_0[4583:4576];
        layer4[62][15:8] = buffer_data_0[4591:4584];
        layer4[62][23:16] = buffer_data_0[4599:4592];
        layer4[62][31:24] = buffer_data_0[4607:4600];
        layer4[62][39:32] = buffer_data_0[4615:4608];
        layer0[63][7:0] = buffer_data_4[4591:4584];
        layer0[63][15:8] = buffer_data_4[4599:4592];
        layer0[63][23:16] = buffer_data_4[4607:4600];
        layer0[63][31:24] = buffer_data_4[4615:4608];
        layer0[63][39:32] = buffer_data_4[4623:4616];
        layer1[63][7:0] = buffer_data_3[4591:4584];
        layer1[63][15:8] = buffer_data_3[4599:4592];
        layer1[63][23:16] = buffer_data_3[4607:4600];
        layer1[63][31:24] = buffer_data_3[4615:4608];
        layer1[63][39:32] = buffer_data_3[4623:4616];
        layer2[63][7:0] = buffer_data_2[4591:4584];
        layer2[63][15:8] = buffer_data_2[4599:4592];
        layer2[63][23:16] = buffer_data_2[4607:4600];
        layer2[63][31:24] = buffer_data_2[4615:4608];
        layer2[63][39:32] = buffer_data_2[4623:4616];
        layer3[63][7:0] = buffer_data_1[4591:4584];
        layer3[63][15:8] = buffer_data_1[4599:4592];
        layer3[63][23:16] = buffer_data_1[4607:4600];
        layer3[63][31:24] = buffer_data_1[4615:4608];
        layer3[63][39:32] = buffer_data_1[4623:4616];
        layer4[63][7:0] = buffer_data_0[4591:4584];
        layer4[63][15:8] = buffer_data_0[4599:4592];
        layer4[63][23:16] = buffer_data_0[4607:4600];
        layer4[63][31:24] = buffer_data_0[4615:4608];
        layer4[63][39:32] = buffer_data_0[4623:4616];
    end
    ST_GAUSSIAN_9: begin
        layer0[0][7:0] = buffer_data_4[4599:4592];
        layer0[0][15:8] = buffer_data_4[4607:4600];
        layer0[0][23:16] = buffer_data_4[4615:4608];
        layer0[0][31:24] = buffer_data_4[4623:4616];
        layer0[0][39:32] = buffer_data_4[4631:4624];
        layer1[0][7:0] = buffer_data_3[4599:4592];
        layer1[0][15:8] = buffer_data_3[4607:4600];
        layer1[0][23:16] = buffer_data_3[4615:4608];
        layer1[0][31:24] = buffer_data_3[4623:4616];
        layer1[0][39:32] = buffer_data_3[4631:4624];
        layer2[0][7:0] = buffer_data_2[4599:4592];
        layer2[0][15:8] = buffer_data_2[4607:4600];
        layer2[0][23:16] = buffer_data_2[4615:4608];
        layer2[0][31:24] = buffer_data_2[4623:4616];
        layer2[0][39:32] = buffer_data_2[4631:4624];
        layer3[0][7:0] = buffer_data_1[4599:4592];
        layer3[0][15:8] = buffer_data_1[4607:4600];
        layer3[0][23:16] = buffer_data_1[4615:4608];
        layer3[0][31:24] = buffer_data_1[4623:4616];
        layer3[0][39:32] = buffer_data_1[4631:4624];
        layer4[0][7:0] = buffer_data_0[4599:4592];
        layer4[0][15:8] = buffer_data_0[4607:4600];
        layer4[0][23:16] = buffer_data_0[4615:4608];
        layer4[0][31:24] = buffer_data_0[4623:4616];
        layer4[0][39:32] = buffer_data_0[4631:4624];
        layer0[1][7:0] = buffer_data_4[4607:4600];
        layer0[1][15:8] = buffer_data_4[4615:4608];
        layer0[1][23:16] = buffer_data_4[4623:4616];
        layer0[1][31:24] = buffer_data_4[4631:4624];
        layer0[1][39:32] = buffer_data_4[4639:4632];
        layer1[1][7:0] = buffer_data_3[4607:4600];
        layer1[1][15:8] = buffer_data_3[4615:4608];
        layer1[1][23:16] = buffer_data_3[4623:4616];
        layer1[1][31:24] = buffer_data_3[4631:4624];
        layer1[1][39:32] = buffer_data_3[4639:4632];
        layer2[1][7:0] = buffer_data_2[4607:4600];
        layer2[1][15:8] = buffer_data_2[4615:4608];
        layer2[1][23:16] = buffer_data_2[4623:4616];
        layer2[1][31:24] = buffer_data_2[4631:4624];
        layer2[1][39:32] = buffer_data_2[4639:4632];
        layer3[1][7:0] = buffer_data_1[4607:4600];
        layer3[1][15:8] = buffer_data_1[4615:4608];
        layer3[1][23:16] = buffer_data_1[4623:4616];
        layer3[1][31:24] = buffer_data_1[4631:4624];
        layer3[1][39:32] = buffer_data_1[4639:4632];
        layer4[1][7:0] = buffer_data_0[4607:4600];
        layer4[1][15:8] = buffer_data_0[4615:4608];
        layer4[1][23:16] = buffer_data_0[4623:4616];
        layer4[1][31:24] = buffer_data_0[4631:4624];
        layer4[1][39:32] = buffer_data_0[4639:4632];
        layer0[2][7:0] = buffer_data_4[4615:4608];
        layer0[2][15:8] = buffer_data_4[4623:4616];
        layer0[2][23:16] = buffer_data_4[4631:4624];
        layer0[2][31:24] = buffer_data_4[4639:4632];
        layer0[2][39:32] = buffer_data_4[4647:4640];
        layer1[2][7:0] = buffer_data_3[4615:4608];
        layer1[2][15:8] = buffer_data_3[4623:4616];
        layer1[2][23:16] = buffer_data_3[4631:4624];
        layer1[2][31:24] = buffer_data_3[4639:4632];
        layer1[2][39:32] = buffer_data_3[4647:4640];
        layer2[2][7:0] = buffer_data_2[4615:4608];
        layer2[2][15:8] = buffer_data_2[4623:4616];
        layer2[2][23:16] = buffer_data_2[4631:4624];
        layer2[2][31:24] = buffer_data_2[4639:4632];
        layer2[2][39:32] = buffer_data_2[4647:4640];
        layer3[2][7:0] = buffer_data_1[4615:4608];
        layer3[2][15:8] = buffer_data_1[4623:4616];
        layer3[2][23:16] = buffer_data_1[4631:4624];
        layer3[2][31:24] = buffer_data_1[4639:4632];
        layer3[2][39:32] = buffer_data_1[4647:4640];
        layer4[2][7:0] = buffer_data_0[4615:4608];
        layer4[2][15:8] = buffer_data_0[4623:4616];
        layer4[2][23:16] = buffer_data_0[4631:4624];
        layer4[2][31:24] = buffer_data_0[4639:4632];
        layer4[2][39:32] = buffer_data_0[4647:4640];
        layer0[3][7:0] = buffer_data_4[4623:4616];
        layer0[3][15:8] = buffer_data_4[4631:4624];
        layer0[3][23:16] = buffer_data_4[4639:4632];
        layer0[3][31:24] = buffer_data_4[4647:4640];
        layer0[3][39:32] = buffer_data_4[4655:4648];
        layer1[3][7:0] = buffer_data_3[4623:4616];
        layer1[3][15:8] = buffer_data_3[4631:4624];
        layer1[3][23:16] = buffer_data_3[4639:4632];
        layer1[3][31:24] = buffer_data_3[4647:4640];
        layer1[3][39:32] = buffer_data_3[4655:4648];
        layer2[3][7:0] = buffer_data_2[4623:4616];
        layer2[3][15:8] = buffer_data_2[4631:4624];
        layer2[3][23:16] = buffer_data_2[4639:4632];
        layer2[3][31:24] = buffer_data_2[4647:4640];
        layer2[3][39:32] = buffer_data_2[4655:4648];
        layer3[3][7:0] = buffer_data_1[4623:4616];
        layer3[3][15:8] = buffer_data_1[4631:4624];
        layer3[3][23:16] = buffer_data_1[4639:4632];
        layer3[3][31:24] = buffer_data_1[4647:4640];
        layer3[3][39:32] = buffer_data_1[4655:4648];
        layer4[3][7:0] = buffer_data_0[4623:4616];
        layer4[3][15:8] = buffer_data_0[4631:4624];
        layer4[3][23:16] = buffer_data_0[4639:4632];
        layer4[3][31:24] = buffer_data_0[4647:4640];
        layer4[3][39:32] = buffer_data_0[4655:4648];
        layer0[4][7:0] = buffer_data_4[4631:4624];
        layer0[4][15:8] = buffer_data_4[4639:4632];
        layer0[4][23:16] = buffer_data_4[4647:4640];
        layer0[4][31:24] = buffer_data_4[4655:4648];
        layer0[4][39:32] = buffer_data_4[4663:4656];
        layer1[4][7:0] = buffer_data_3[4631:4624];
        layer1[4][15:8] = buffer_data_3[4639:4632];
        layer1[4][23:16] = buffer_data_3[4647:4640];
        layer1[4][31:24] = buffer_data_3[4655:4648];
        layer1[4][39:32] = buffer_data_3[4663:4656];
        layer2[4][7:0] = buffer_data_2[4631:4624];
        layer2[4][15:8] = buffer_data_2[4639:4632];
        layer2[4][23:16] = buffer_data_2[4647:4640];
        layer2[4][31:24] = buffer_data_2[4655:4648];
        layer2[4][39:32] = buffer_data_2[4663:4656];
        layer3[4][7:0] = buffer_data_1[4631:4624];
        layer3[4][15:8] = buffer_data_1[4639:4632];
        layer3[4][23:16] = buffer_data_1[4647:4640];
        layer3[4][31:24] = buffer_data_1[4655:4648];
        layer3[4][39:32] = buffer_data_1[4663:4656];
        layer4[4][7:0] = buffer_data_0[4631:4624];
        layer4[4][15:8] = buffer_data_0[4639:4632];
        layer4[4][23:16] = buffer_data_0[4647:4640];
        layer4[4][31:24] = buffer_data_0[4655:4648];
        layer4[4][39:32] = buffer_data_0[4663:4656];
        layer0[5][7:0] = buffer_data_4[4639:4632];
        layer0[5][15:8] = buffer_data_4[4647:4640];
        layer0[5][23:16] = buffer_data_4[4655:4648];
        layer0[5][31:24] = buffer_data_4[4663:4656];
        layer0[5][39:32] = buffer_data_4[4671:4664];
        layer1[5][7:0] = buffer_data_3[4639:4632];
        layer1[5][15:8] = buffer_data_3[4647:4640];
        layer1[5][23:16] = buffer_data_3[4655:4648];
        layer1[5][31:24] = buffer_data_3[4663:4656];
        layer1[5][39:32] = buffer_data_3[4671:4664];
        layer2[5][7:0] = buffer_data_2[4639:4632];
        layer2[5][15:8] = buffer_data_2[4647:4640];
        layer2[5][23:16] = buffer_data_2[4655:4648];
        layer2[5][31:24] = buffer_data_2[4663:4656];
        layer2[5][39:32] = buffer_data_2[4671:4664];
        layer3[5][7:0] = buffer_data_1[4639:4632];
        layer3[5][15:8] = buffer_data_1[4647:4640];
        layer3[5][23:16] = buffer_data_1[4655:4648];
        layer3[5][31:24] = buffer_data_1[4663:4656];
        layer3[5][39:32] = buffer_data_1[4671:4664];
        layer4[5][7:0] = buffer_data_0[4639:4632];
        layer4[5][15:8] = buffer_data_0[4647:4640];
        layer4[5][23:16] = buffer_data_0[4655:4648];
        layer4[5][31:24] = buffer_data_0[4663:4656];
        layer4[5][39:32] = buffer_data_0[4671:4664];
        layer0[6][7:0] = buffer_data_4[4647:4640];
        layer0[6][15:8] = buffer_data_4[4655:4648];
        layer0[6][23:16] = buffer_data_4[4663:4656];
        layer0[6][31:24] = buffer_data_4[4671:4664];
        layer0[6][39:32] = buffer_data_4[4679:4672];
        layer1[6][7:0] = buffer_data_3[4647:4640];
        layer1[6][15:8] = buffer_data_3[4655:4648];
        layer1[6][23:16] = buffer_data_3[4663:4656];
        layer1[6][31:24] = buffer_data_3[4671:4664];
        layer1[6][39:32] = buffer_data_3[4679:4672];
        layer2[6][7:0] = buffer_data_2[4647:4640];
        layer2[6][15:8] = buffer_data_2[4655:4648];
        layer2[6][23:16] = buffer_data_2[4663:4656];
        layer2[6][31:24] = buffer_data_2[4671:4664];
        layer2[6][39:32] = buffer_data_2[4679:4672];
        layer3[6][7:0] = buffer_data_1[4647:4640];
        layer3[6][15:8] = buffer_data_1[4655:4648];
        layer3[6][23:16] = buffer_data_1[4663:4656];
        layer3[6][31:24] = buffer_data_1[4671:4664];
        layer3[6][39:32] = buffer_data_1[4679:4672];
        layer4[6][7:0] = buffer_data_0[4647:4640];
        layer4[6][15:8] = buffer_data_0[4655:4648];
        layer4[6][23:16] = buffer_data_0[4663:4656];
        layer4[6][31:24] = buffer_data_0[4671:4664];
        layer4[6][39:32] = buffer_data_0[4679:4672];
        layer0[7][7:0] = buffer_data_4[4655:4648];
        layer0[7][15:8] = buffer_data_4[4663:4656];
        layer0[7][23:16] = buffer_data_4[4671:4664];
        layer0[7][31:24] = buffer_data_4[4679:4672];
        layer0[7][39:32] = buffer_data_4[4687:4680];
        layer1[7][7:0] = buffer_data_3[4655:4648];
        layer1[7][15:8] = buffer_data_3[4663:4656];
        layer1[7][23:16] = buffer_data_3[4671:4664];
        layer1[7][31:24] = buffer_data_3[4679:4672];
        layer1[7][39:32] = buffer_data_3[4687:4680];
        layer2[7][7:0] = buffer_data_2[4655:4648];
        layer2[7][15:8] = buffer_data_2[4663:4656];
        layer2[7][23:16] = buffer_data_2[4671:4664];
        layer2[7][31:24] = buffer_data_2[4679:4672];
        layer2[7][39:32] = buffer_data_2[4687:4680];
        layer3[7][7:0] = buffer_data_1[4655:4648];
        layer3[7][15:8] = buffer_data_1[4663:4656];
        layer3[7][23:16] = buffer_data_1[4671:4664];
        layer3[7][31:24] = buffer_data_1[4679:4672];
        layer3[7][39:32] = buffer_data_1[4687:4680];
        layer4[7][7:0] = buffer_data_0[4655:4648];
        layer4[7][15:8] = buffer_data_0[4663:4656];
        layer4[7][23:16] = buffer_data_0[4671:4664];
        layer4[7][31:24] = buffer_data_0[4679:4672];
        layer4[7][39:32] = buffer_data_0[4687:4680];
        layer0[8][7:0] = buffer_data_4[4663:4656];
        layer0[8][15:8] = buffer_data_4[4671:4664];
        layer0[8][23:16] = buffer_data_4[4679:4672];
        layer0[8][31:24] = buffer_data_4[4687:4680];
        layer0[8][39:32] = buffer_data_4[4695:4688];
        layer1[8][7:0] = buffer_data_3[4663:4656];
        layer1[8][15:8] = buffer_data_3[4671:4664];
        layer1[8][23:16] = buffer_data_3[4679:4672];
        layer1[8][31:24] = buffer_data_3[4687:4680];
        layer1[8][39:32] = buffer_data_3[4695:4688];
        layer2[8][7:0] = buffer_data_2[4663:4656];
        layer2[8][15:8] = buffer_data_2[4671:4664];
        layer2[8][23:16] = buffer_data_2[4679:4672];
        layer2[8][31:24] = buffer_data_2[4687:4680];
        layer2[8][39:32] = buffer_data_2[4695:4688];
        layer3[8][7:0] = buffer_data_1[4663:4656];
        layer3[8][15:8] = buffer_data_1[4671:4664];
        layer3[8][23:16] = buffer_data_1[4679:4672];
        layer3[8][31:24] = buffer_data_1[4687:4680];
        layer3[8][39:32] = buffer_data_1[4695:4688];
        layer4[8][7:0] = buffer_data_0[4663:4656];
        layer4[8][15:8] = buffer_data_0[4671:4664];
        layer4[8][23:16] = buffer_data_0[4679:4672];
        layer4[8][31:24] = buffer_data_0[4687:4680];
        layer4[8][39:32] = buffer_data_0[4695:4688];
        layer0[9][7:0] = buffer_data_4[4671:4664];
        layer0[9][15:8] = buffer_data_4[4679:4672];
        layer0[9][23:16] = buffer_data_4[4687:4680];
        layer0[9][31:24] = buffer_data_4[4695:4688];
        layer0[9][39:32] = buffer_data_4[4703:4696];
        layer1[9][7:0] = buffer_data_3[4671:4664];
        layer1[9][15:8] = buffer_data_3[4679:4672];
        layer1[9][23:16] = buffer_data_3[4687:4680];
        layer1[9][31:24] = buffer_data_3[4695:4688];
        layer1[9][39:32] = buffer_data_3[4703:4696];
        layer2[9][7:0] = buffer_data_2[4671:4664];
        layer2[9][15:8] = buffer_data_2[4679:4672];
        layer2[9][23:16] = buffer_data_2[4687:4680];
        layer2[9][31:24] = buffer_data_2[4695:4688];
        layer2[9][39:32] = buffer_data_2[4703:4696];
        layer3[9][7:0] = buffer_data_1[4671:4664];
        layer3[9][15:8] = buffer_data_1[4679:4672];
        layer3[9][23:16] = buffer_data_1[4687:4680];
        layer3[9][31:24] = buffer_data_1[4695:4688];
        layer3[9][39:32] = buffer_data_1[4703:4696];
        layer4[9][7:0] = buffer_data_0[4671:4664];
        layer4[9][15:8] = buffer_data_0[4679:4672];
        layer4[9][23:16] = buffer_data_0[4687:4680];
        layer4[9][31:24] = buffer_data_0[4695:4688];
        layer4[9][39:32] = buffer_data_0[4703:4696];
        layer0[10][7:0] = buffer_data_4[4679:4672];
        layer0[10][15:8] = buffer_data_4[4687:4680];
        layer0[10][23:16] = buffer_data_4[4695:4688];
        layer0[10][31:24] = buffer_data_4[4703:4696];
        layer0[10][39:32] = buffer_data_4[4711:4704];
        layer1[10][7:0] = buffer_data_3[4679:4672];
        layer1[10][15:8] = buffer_data_3[4687:4680];
        layer1[10][23:16] = buffer_data_3[4695:4688];
        layer1[10][31:24] = buffer_data_3[4703:4696];
        layer1[10][39:32] = buffer_data_3[4711:4704];
        layer2[10][7:0] = buffer_data_2[4679:4672];
        layer2[10][15:8] = buffer_data_2[4687:4680];
        layer2[10][23:16] = buffer_data_2[4695:4688];
        layer2[10][31:24] = buffer_data_2[4703:4696];
        layer2[10][39:32] = buffer_data_2[4711:4704];
        layer3[10][7:0] = buffer_data_1[4679:4672];
        layer3[10][15:8] = buffer_data_1[4687:4680];
        layer3[10][23:16] = buffer_data_1[4695:4688];
        layer3[10][31:24] = buffer_data_1[4703:4696];
        layer3[10][39:32] = buffer_data_1[4711:4704];
        layer4[10][7:0] = buffer_data_0[4679:4672];
        layer4[10][15:8] = buffer_data_0[4687:4680];
        layer4[10][23:16] = buffer_data_0[4695:4688];
        layer4[10][31:24] = buffer_data_0[4703:4696];
        layer4[10][39:32] = buffer_data_0[4711:4704];
        layer0[11][7:0] = buffer_data_4[4687:4680];
        layer0[11][15:8] = buffer_data_4[4695:4688];
        layer0[11][23:16] = buffer_data_4[4703:4696];
        layer0[11][31:24] = buffer_data_4[4711:4704];
        layer0[11][39:32] = buffer_data_4[4719:4712];
        layer1[11][7:0] = buffer_data_3[4687:4680];
        layer1[11][15:8] = buffer_data_3[4695:4688];
        layer1[11][23:16] = buffer_data_3[4703:4696];
        layer1[11][31:24] = buffer_data_3[4711:4704];
        layer1[11][39:32] = buffer_data_3[4719:4712];
        layer2[11][7:0] = buffer_data_2[4687:4680];
        layer2[11][15:8] = buffer_data_2[4695:4688];
        layer2[11][23:16] = buffer_data_2[4703:4696];
        layer2[11][31:24] = buffer_data_2[4711:4704];
        layer2[11][39:32] = buffer_data_2[4719:4712];
        layer3[11][7:0] = buffer_data_1[4687:4680];
        layer3[11][15:8] = buffer_data_1[4695:4688];
        layer3[11][23:16] = buffer_data_1[4703:4696];
        layer3[11][31:24] = buffer_data_1[4711:4704];
        layer3[11][39:32] = buffer_data_1[4719:4712];
        layer4[11][7:0] = buffer_data_0[4687:4680];
        layer4[11][15:8] = buffer_data_0[4695:4688];
        layer4[11][23:16] = buffer_data_0[4703:4696];
        layer4[11][31:24] = buffer_data_0[4711:4704];
        layer4[11][39:32] = buffer_data_0[4719:4712];
        layer0[12][7:0] = buffer_data_4[4695:4688];
        layer0[12][15:8] = buffer_data_4[4703:4696];
        layer0[12][23:16] = buffer_data_4[4711:4704];
        layer0[12][31:24] = buffer_data_4[4719:4712];
        layer0[12][39:32] = buffer_data_4[4727:4720];
        layer1[12][7:0] = buffer_data_3[4695:4688];
        layer1[12][15:8] = buffer_data_3[4703:4696];
        layer1[12][23:16] = buffer_data_3[4711:4704];
        layer1[12][31:24] = buffer_data_3[4719:4712];
        layer1[12][39:32] = buffer_data_3[4727:4720];
        layer2[12][7:0] = buffer_data_2[4695:4688];
        layer2[12][15:8] = buffer_data_2[4703:4696];
        layer2[12][23:16] = buffer_data_2[4711:4704];
        layer2[12][31:24] = buffer_data_2[4719:4712];
        layer2[12][39:32] = buffer_data_2[4727:4720];
        layer3[12][7:0] = buffer_data_1[4695:4688];
        layer3[12][15:8] = buffer_data_1[4703:4696];
        layer3[12][23:16] = buffer_data_1[4711:4704];
        layer3[12][31:24] = buffer_data_1[4719:4712];
        layer3[12][39:32] = buffer_data_1[4727:4720];
        layer4[12][7:0] = buffer_data_0[4695:4688];
        layer4[12][15:8] = buffer_data_0[4703:4696];
        layer4[12][23:16] = buffer_data_0[4711:4704];
        layer4[12][31:24] = buffer_data_0[4719:4712];
        layer4[12][39:32] = buffer_data_0[4727:4720];
        layer0[13][7:0] = buffer_data_4[4703:4696];
        layer0[13][15:8] = buffer_data_4[4711:4704];
        layer0[13][23:16] = buffer_data_4[4719:4712];
        layer0[13][31:24] = buffer_data_4[4727:4720];
        layer0[13][39:32] = buffer_data_4[4735:4728];
        layer1[13][7:0] = buffer_data_3[4703:4696];
        layer1[13][15:8] = buffer_data_3[4711:4704];
        layer1[13][23:16] = buffer_data_3[4719:4712];
        layer1[13][31:24] = buffer_data_3[4727:4720];
        layer1[13][39:32] = buffer_data_3[4735:4728];
        layer2[13][7:0] = buffer_data_2[4703:4696];
        layer2[13][15:8] = buffer_data_2[4711:4704];
        layer2[13][23:16] = buffer_data_2[4719:4712];
        layer2[13][31:24] = buffer_data_2[4727:4720];
        layer2[13][39:32] = buffer_data_2[4735:4728];
        layer3[13][7:0] = buffer_data_1[4703:4696];
        layer3[13][15:8] = buffer_data_1[4711:4704];
        layer3[13][23:16] = buffer_data_1[4719:4712];
        layer3[13][31:24] = buffer_data_1[4727:4720];
        layer3[13][39:32] = buffer_data_1[4735:4728];
        layer4[13][7:0] = buffer_data_0[4703:4696];
        layer4[13][15:8] = buffer_data_0[4711:4704];
        layer4[13][23:16] = buffer_data_0[4719:4712];
        layer4[13][31:24] = buffer_data_0[4727:4720];
        layer4[13][39:32] = buffer_data_0[4735:4728];
        layer0[14][7:0] = buffer_data_4[4711:4704];
        layer0[14][15:8] = buffer_data_4[4719:4712];
        layer0[14][23:16] = buffer_data_4[4727:4720];
        layer0[14][31:24] = buffer_data_4[4735:4728];
        layer0[14][39:32] = buffer_data_4[4743:4736];
        layer1[14][7:0] = buffer_data_3[4711:4704];
        layer1[14][15:8] = buffer_data_3[4719:4712];
        layer1[14][23:16] = buffer_data_3[4727:4720];
        layer1[14][31:24] = buffer_data_3[4735:4728];
        layer1[14][39:32] = buffer_data_3[4743:4736];
        layer2[14][7:0] = buffer_data_2[4711:4704];
        layer2[14][15:8] = buffer_data_2[4719:4712];
        layer2[14][23:16] = buffer_data_2[4727:4720];
        layer2[14][31:24] = buffer_data_2[4735:4728];
        layer2[14][39:32] = buffer_data_2[4743:4736];
        layer3[14][7:0] = buffer_data_1[4711:4704];
        layer3[14][15:8] = buffer_data_1[4719:4712];
        layer3[14][23:16] = buffer_data_1[4727:4720];
        layer3[14][31:24] = buffer_data_1[4735:4728];
        layer3[14][39:32] = buffer_data_1[4743:4736];
        layer4[14][7:0] = buffer_data_0[4711:4704];
        layer4[14][15:8] = buffer_data_0[4719:4712];
        layer4[14][23:16] = buffer_data_0[4727:4720];
        layer4[14][31:24] = buffer_data_0[4735:4728];
        layer4[14][39:32] = buffer_data_0[4743:4736];
        layer0[15][7:0] = buffer_data_4[4719:4712];
        layer0[15][15:8] = buffer_data_4[4727:4720];
        layer0[15][23:16] = buffer_data_4[4735:4728];
        layer0[15][31:24] = buffer_data_4[4743:4736];
        layer0[15][39:32] = buffer_data_4[4751:4744];
        layer1[15][7:0] = buffer_data_3[4719:4712];
        layer1[15][15:8] = buffer_data_3[4727:4720];
        layer1[15][23:16] = buffer_data_3[4735:4728];
        layer1[15][31:24] = buffer_data_3[4743:4736];
        layer1[15][39:32] = buffer_data_3[4751:4744];
        layer2[15][7:0] = buffer_data_2[4719:4712];
        layer2[15][15:8] = buffer_data_2[4727:4720];
        layer2[15][23:16] = buffer_data_2[4735:4728];
        layer2[15][31:24] = buffer_data_2[4743:4736];
        layer2[15][39:32] = buffer_data_2[4751:4744];
        layer3[15][7:0] = buffer_data_1[4719:4712];
        layer3[15][15:8] = buffer_data_1[4727:4720];
        layer3[15][23:16] = buffer_data_1[4735:4728];
        layer3[15][31:24] = buffer_data_1[4743:4736];
        layer3[15][39:32] = buffer_data_1[4751:4744];
        layer4[15][7:0] = buffer_data_0[4719:4712];
        layer4[15][15:8] = buffer_data_0[4727:4720];
        layer4[15][23:16] = buffer_data_0[4735:4728];
        layer4[15][31:24] = buffer_data_0[4743:4736];
        layer4[15][39:32] = buffer_data_0[4751:4744];
        layer0[16][7:0] = buffer_data_4[4727:4720];
        layer0[16][15:8] = buffer_data_4[4735:4728];
        layer0[16][23:16] = buffer_data_4[4743:4736];
        layer0[16][31:24] = buffer_data_4[4751:4744];
        layer0[16][39:32] = buffer_data_4[4759:4752];
        layer1[16][7:0] = buffer_data_3[4727:4720];
        layer1[16][15:8] = buffer_data_3[4735:4728];
        layer1[16][23:16] = buffer_data_3[4743:4736];
        layer1[16][31:24] = buffer_data_3[4751:4744];
        layer1[16][39:32] = buffer_data_3[4759:4752];
        layer2[16][7:0] = buffer_data_2[4727:4720];
        layer2[16][15:8] = buffer_data_2[4735:4728];
        layer2[16][23:16] = buffer_data_2[4743:4736];
        layer2[16][31:24] = buffer_data_2[4751:4744];
        layer2[16][39:32] = buffer_data_2[4759:4752];
        layer3[16][7:0] = buffer_data_1[4727:4720];
        layer3[16][15:8] = buffer_data_1[4735:4728];
        layer3[16][23:16] = buffer_data_1[4743:4736];
        layer3[16][31:24] = buffer_data_1[4751:4744];
        layer3[16][39:32] = buffer_data_1[4759:4752];
        layer4[16][7:0] = buffer_data_0[4727:4720];
        layer4[16][15:8] = buffer_data_0[4735:4728];
        layer4[16][23:16] = buffer_data_0[4743:4736];
        layer4[16][31:24] = buffer_data_0[4751:4744];
        layer4[16][39:32] = buffer_data_0[4759:4752];
        layer0[17][7:0] = buffer_data_4[4735:4728];
        layer0[17][15:8] = buffer_data_4[4743:4736];
        layer0[17][23:16] = buffer_data_4[4751:4744];
        layer0[17][31:24] = buffer_data_4[4759:4752];
        layer0[17][39:32] = buffer_data_4[4767:4760];
        layer1[17][7:0] = buffer_data_3[4735:4728];
        layer1[17][15:8] = buffer_data_3[4743:4736];
        layer1[17][23:16] = buffer_data_3[4751:4744];
        layer1[17][31:24] = buffer_data_3[4759:4752];
        layer1[17][39:32] = buffer_data_3[4767:4760];
        layer2[17][7:0] = buffer_data_2[4735:4728];
        layer2[17][15:8] = buffer_data_2[4743:4736];
        layer2[17][23:16] = buffer_data_2[4751:4744];
        layer2[17][31:24] = buffer_data_2[4759:4752];
        layer2[17][39:32] = buffer_data_2[4767:4760];
        layer3[17][7:0] = buffer_data_1[4735:4728];
        layer3[17][15:8] = buffer_data_1[4743:4736];
        layer3[17][23:16] = buffer_data_1[4751:4744];
        layer3[17][31:24] = buffer_data_1[4759:4752];
        layer3[17][39:32] = buffer_data_1[4767:4760];
        layer4[17][7:0] = buffer_data_0[4735:4728];
        layer4[17][15:8] = buffer_data_0[4743:4736];
        layer4[17][23:16] = buffer_data_0[4751:4744];
        layer4[17][31:24] = buffer_data_0[4759:4752];
        layer4[17][39:32] = buffer_data_0[4767:4760];
        layer0[18][7:0] = buffer_data_4[4743:4736];
        layer0[18][15:8] = buffer_data_4[4751:4744];
        layer0[18][23:16] = buffer_data_4[4759:4752];
        layer0[18][31:24] = buffer_data_4[4767:4760];
        layer0[18][39:32] = buffer_data_4[4775:4768];
        layer1[18][7:0] = buffer_data_3[4743:4736];
        layer1[18][15:8] = buffer_data_3[4751:4744];
        layer1[18][23:16] = buffer_data_3[4759:4752];
        layer1[18][31:24] = buffer_data_3[4767:4760];
        layer1[18][39:32] = buffer_data_3[4775:4768];
        layer2[18][7:0] = buffer_data_2[4743:4736];
        layer2[18][15:8] = buffer_data_2[4751:4744];
        layer2[18][23:16] = buffer_data_2[4759:4752];
        layer2[18][31:24] = buffer_data_2[4767:4760];
        layer2[18][39:32] = buffer_data_2[4775:4768];
        layer3[18][7:0] = buffer_data_1[4743:4736];
        layer3[18][15:8] = buffer_data_1[4751:4744];
        layer3[18][23:16] = buffer_data_1[4759:4752];
        layer3[18][31:24] = buffer_data_1[4767:4760];
        layer3[18][39:32] = buffer_data_1[4775:4768];
        layer4[18][7:0] = buffer_data_0[4743:4736];
        layer4[18][15:8] = buffer_data_0[4751:4744];
        layer4[18][23:16] = buffer_data_0[4759:4752];
        layer4[18][31:24] = buffer_data_0[4767:4760];
        layer4[18][39:32] = buffer_data_0[4775:4768];
        layer0[19][7:0] = buffer_data_4[4751:4744];
        layer0[19][15:8] = buffer_data_4[4759:4752];
        layer0[19][23:16] = buffer_data_4[4767:4760];
        layer0[19][31:24] = buffer_data_4[4775:4768];
        layer0[19][39:32] = buffer_data_4[4783:4776];
        layer1[19][7:0] = buffer_data_3[4751:4744];
        layer1[19][15:8] = buffer_data_3[4759:4752];
        layer1[19][23:16] = buffer_data_3[4767:4760];
        layer1[19][31:24] = buffer_data_3[4775:4768];
        layer1[19][39:32] = buffer_data_3[4783:4776];
        layer2[19][7:0] = buffer_data_2[4751:4744];
        layer2[19][15:8] = buffer_data_2[4759:4752];
        layer2[19][23:16] = buffer_data_2[4767:4760];
        layer2[19][31:24] = buffer_data_2[4775:4768];
        layer2[19][39:32] = buffer_data_2[4783:4776];
        layer3[19][7:0] = buffer_data_1[4751:4744];
        layer3[19][15:8] = buffer_data_1[4759:4752];
        layer3[19][23:16] = buffer_data_1[4767:4760];
        layer3[19][31:24] = buffer_data_1[4775:4768];
        layer3[19][39:32] = buffer_data_1[4783:4776];
        layer4[19][7:0] = buffer_data_0[4751:4744];
        layer4[19][15:8] = buffer_data_0[4759:4752];
        layer4[19][23:16] = buffer_data_0[4767:4760];
        layer4[19][31:24] = buffer_data_0[4775:4768];
        layer4[19][39:32] = buffer_data_0[4783:4776];
        layer0[20][7:0] = buffer_data_4[4759:4752];
        layer0[20][15:8] = buffer_data_4[4767:4760];
        layer0[20][23:16] = buffer_data_4[4775:4768];
        layer0[20][31:24] = buffer_data_4[4783:4776];
        layer0[20][39:32] = buffer_data_4[4791:4784];
        layer1[20][7:0] = buffer_data_3[4759:4752];
        layer1[20][15:8] = buffer_data_3[4767:4760];
        layer1[20][23:16] = buffer_data_3[4775:4768];
        layer1[20][31:24] = buffer_data_3[4783:4776];
        layer1[20][39:32] = buffer_data_3[4791:4784];
        layer2[20][7:0] = buffer_data_2[4759:4752];
        layer2[20][15:8] = buffer_data_2[4767:4760];
        layer2[20][23:16] = buffer_data_2[4775:4768];
        layer2[20][31:24] = buffer_data_2[4783:4776];
        layer2[20][39:32] = buffer_data_2[4791:4784];
        layer3[20][7:0] = buffer_data_1[4759:4752];
        layer3[20][15:8] = buffer_data_1[4767:4760];
        layer3[20][23:16] = buffer_data_1[4775:4768];
        layer3[20][31:24] = buffer_data_1[4783:4776];
        layer3[20][39:32] = buffer_data_1[4791:4784];
        layer4[20][7:0] = buffer_data_0[4759:4752];
        layer4[20][15:8] = buffer_data_0[4767:4760];
        layer4[20][23:16] = buffer_data_0[4775:4768];
        layer4[20][31:24] = buffer_data_0[4783:4776];
        layer4[20][39:32] = buffer_data_0[4791:4784];
        layer0[21][7:0] = buffer_data_4[4767:4760];
        layer0[21][15:8] = buffer_data_4[4775:4768];
        layer0[21][23:16] = buffer_data_4[4783:4776];
        layer0[21][31:24] = buffer_data_4[4791:4784];
        layer0[21][39:32] = buffer_data_4[4799:4792];
        layer1[21][7:0] = buffer_data_3[4767:4760];
        layer1[21][15:8] = buffer_data_3[4775:4768];
        layer1[21][23:16] = buffer_data_3[4783:4776];
        layer1[21][31:24] = buffer_data_3[4791:4784];
        layer1[21][39:32] = buffer_data_3[4799:4792];
        layer2[21][7:0] = buffer_data_2[4767:4760];
        layer2[21][15:8] = buffer_data_2[4775:4768];
        layer2[21][23:16] = buffer_data_2[4783:4776];
        layer2[21][31:24] = buffer_data_2[4791:4784];
        layer2[21][39:32] = buffer_data_2[4799:4792];
        layer3[21][7:0] = buffer_data_1[4767:4760];
        layer3[21][15:8] = buffer_data_1[4775:4768];
        layer3[21][23:16] = buffer_data_1[4783:4776];
        layer3[21][31:24] = buffer_data_1[4791:4784];
        layer3[21][39:32] = buffer_data_1[4799:4792];
        layer4[21][7:0] = buffer_data_0[4767:4760];
        layer4[21][15:8] = buffer_data_0[4775:4768];
        layer4[21][23:16] = buffer_data_0[4783:4776];
        layer4[21][31:24] = buffer_data_0[4791:4784];
        layer4[21][39:32] = buffer_data_0[4799:4792];
        layer0[22][7:0] = buffer_data_4[4775:4768];
        layer0[22][15:8] = buffer_data_4[4783:4776];
        layer0[22][23:16] = buffer_data_4[4791:4784];
        layer0[22][31:24] = buffer_data_4[4799:4792];
        layer0[22][39:32] = buffer_data_4[4807:4800];
        layer1[22][7:0] = buffer_data_3[4775:4768];
        layer1[22][15:8] = buffer_data_3[4783:4776];
        layer1[22][23:16] = buffer_data_3[4791:4784];
        layer1[22][31:24] = buffer_data_3[4799:4792];
        layer1[22][39:32] = buffer_data_3[4807:4800];
        layer2[22][7:0] = buffer_data_2[4775:4768];
        layer2[22][15:8] = buffer_data_2[4783:4776];
        layer2[22][23:16] = buffer_data_2[4791:4784];
        layer2[22][31:24] = buffer_data_2[4799:4792];
        layer2[22][39:32] = buffer_data_2[4807:4800];
        layer3[22][7:0] = buffer_data_1[4775:4768];
        layer3[22][15:8] = buffer_data_1[4783:4776];
        layer3[22][23:16] = buffer_data_1[4791:4784];
        layer3[22][31:24] = buffer_data_1[4799:4792];
        layer3[22][39:32] = buffer_data_1[4807:4800];
        layer4[22][7:0] = buffer_data_0[4775:4768];
        layer4[22][15:8] = buffer_data_0[4783:4776];
        layer4[22][23:16] = buffer_data_0[4791:4784];
        layer4[22][31:24] = buffer_data_0[4799:4792];
        layer4[22][39:32] = buffer_data_0[4807:4800];
        layer0[23][7:0] = buffer_data_4[4783:4776];
        layer0[23][15:8] = buffer_data_4[4791:4784];
        layer0[23][23:16] = buffer_data_4[4799:4792];
        layer0[23][31:24] = buffer_data_4[4807:4800];
        layer0[23][39:32] = buffer_data_4[4815:4808];
        layer1[23][7:0] = buffer_data_3[4783:4776];
        layer1[23][15:8] = buffer_data_3[4791:4784];
        layer1[23][23:16] = buffer_data_3[4799:4792];
        layer1[23][31:24] = buffer_data_3[4807:4800];
        layer1[23][39:32] = buffer_data_3[4815:4808];
        layer2[23][7:0] = buffer_data_2[4783:4776];
        layer2[23][15:8] = buffer_data_2[4791:4784];
        layer2[23][23:16] = buffer_data_2[4799:4792];
        layer2[23][31:24] = buffer_data_2[4807:4800];
        layer2[23][39:32] = buffer_data_2[4815:4808];
        layer3[23][7:0] = buffer_data_1[4783:4776];
        layer3[23][15:8] = buffer_data_1[4791:4784];
        layer3[23][23:16] = buffer_data_1[4799:4792];
        layer3[23][31:24] = buffer_data_1[4807:4800];
        layer3[23][39:32] = buffer_data_1[4815:4808];
        layer4[23][7:0] = buffer_data_0[4783:4776];
        layer4[23][15:8] = buffer_data_0[4791:4784];
        layer4[23][23:16] = buffer_data_0[4799:4792];
        layer4[23][31:24] = buffer_data_0[4807:4800];
        layer4[23][39:32] = buffer_data_0[4815:4808];
        layer0[24][7:0] = buffer_data_4[4791:4784];
        layer0[24][15:8] = buffer_data_4[4799:4792];
        layer0[24][23:16] = buffer_data_4[4807:4800];
        layer0[24][31:24] = buffer_data_4[4815:4808];
        layer0[24][39:32] = buffer_data_4[4823:4816];
        layer1[24][7:0] = buffer_data_3[4791:4784];
        layer1[24][15:8] = buffer_data_3[4799:4792];
        layer1[24][23:16] = buffer_data_3[4807:4800];
        layer1[24][31:24] = buffer_data_3[4815:4808];
        layer1[24][39:32] = buffer_data_3[4823:4816];
        layer2[24][7:0] = buffer_data_2[4791:4784];
        layer2[24][15:8] = buffer_data_2[4799:4792];
        layer2[24][23:16] = buffer_data_2[4807:4800];
        layer2[24][31:24] = buffer_data_2[4815:4808];
        layer2[24][39:32] = buffer_data_2[4823:4816];
        layer3[24][7:0] = buffer_data_1[4791:4784];
        layer3[24][15:8] = buffer_data_1[4799:4792];
        layer3[24][23:16] = buffer_data_1[4807:4800];
        layer3[24][31:24] = buffer_data_1[4815:4808];
        layer3[24][39:32] = buffer_data_1[4823:4816];
        layer4[24][7:0] = buffer_data_0[4791:4784];
        layer4[24][15:8] = buffer_data_0[4799:4792];
        layer4[24][23:16] = buffer_data_0[4807:4800];
        layer4[24][31:24] = buffer_data_0[4815:4808];
        layer4[24][39:32] = buffer_data_0[4823:4816];
        layer0[25][7:0] = buffer_data_4[4799:4792];
        layer0[25][15:8] = buffer_data_4[4807:4800];
        layer0[25][23:16] = buffer_data_4[4815:4808];
        layer0[25][31:24] = buffer_data_4[4823:4816];
        layer0[25][39:32] = buffer_data_4[4831:4824];
        layer1[25][7:0] = buffer_data_3[4799:4792];
        layer1[25][15:8] = buffer_data_3[4807:4800];
        layer1[25][23:16] = buffer_data_3[4815:4808];
        layer1[25][31:24] = buffer_data_3[4823:4816];
        layer1[25][39:32] = buffer_data_3[4831:4824];
        layer2[25][7:0] = buffer_data_2[4799:4792];
        layer2[25][15:8] = buffer_data_2[4807:4800];
        layer2[25][23:16] = buffer_data_2[4815:4808];
        layer2[25][31:24] = buffer_data_2[4823:4816];
        layer2[25][39:32] = buffer_data_2[4831:4824];
        layer3[25][7:0] = buffer_data_1[4799:4792];
        layer3[25][15:8] = buffer_data_1[4807:4800];
        layer3[25][23:16] = buffer_data_1[4815:4808];
        layer3[25][31:24] = buffer_data_1[4823:4816];
        layer3[25][39:32] = buffer_data_1[4831:4824];
        layer4[25][7:0] = buffer_data_0[4799:4792];
        layer4[25][15:8] = buffer_data_0[4807:4800];
        layer4[25][23:16] = buffer_data_0[4815:4808];
        layer4[25][31:24] = buffer_data_0[4823:4816];
        layer4[25][39:32] = buffer_data_0[4831:4824];
        layer0[26][7:0] = buffer_data_4[4807:4800];
        layer0[26][15:8] = buffer_data_4[4815:4808];
        layer0[26][23:16] = buffer_data_4[4823:4816];
        layer0[26][31:24] = buffer_data_4[4831:4824];
        layer0[26][39:32] = buffer_data_4[4839:4832];
        layer1[26][7:0] = buffer_data_3[4807:4800];
        layer1[26][15:8] = buffer_data_3[4815:4808];
        layer1[26][23:16] = buffer_data_3[4823:4816];
        layer1[26][31:24] = buffer_data_3[4831:4824];
        layer1[26][39:32] = buffer_data_3[4839:4832];
        layer2[26][7:0] = buffer_data_2[4807:4800];
        layer2[26][15:8] = buffer_data_2[4815:4808];
        layer2[26][23:16] = buffer_data_2[4823:4816];
        layer2[26][31:24] = buffer_data_2[4831:4824];
        layer2[26][39:32] = buffer_data_2[4839:4832];
        layer3[26][7:0] = buffer_data_1[4807:4800];
        layer3[26][15:8] = buffer_data_1[4815:4808];
        layer3[26][23:16] = buffer_data_1[4823:4816];
        layer3[26][31:24] = buffer_data_1[4831:4824];
        layer3[26][39:32] = buffer_data_1[4839:4832];
        layer4[26][7:0] = buffer_data_0[4807:4800];
        layer4[26][15:8] = buffer_data_0[4815:4808];
        layer4[26][23:16] = buffer_data_0[4823:4816];
        layer4[26][31:24] = buffer_data_0[4831:4824];
        layer4[26][39:32] = buffer_data_0[4839:4832];
        layer0[27][7:0] = buffer_data_4[4815:4808];
        layer0[27][15:8] = buffer_data_4[4823:4816];
        layer0[27][23:16] = buffer_data_4[4831:4824];
        layer0[27][31:24] = buffer_data_4[4839:4832];
        layer0[27][39:32] = buffer_data_4[4847:4840];
        layer1[27][7:0] = buffer_data_3[4815:4808];
        layer1[27][15:8] = buffer_data_3[4823:4816];
        layer1[27][23:16] = buffer_data_3[4831:4824];
        layer1[27][31:24] = buffer_data_3[4839:4832];
        layer1[27][39:32] = buffer_data_3[4847:4840];
        layer2[27][7:0] = buffer_data_2[4815:4808];
        layer2[27][15:8] = buffer_data_2[4823:4816];
        layer2[27][23:16] = buffer_data_2[4831:4824];
        layer2[27][31:24] = buffer_data_2[4839:4832];
        layer2[27][39:32] = buffer_data_2[4847:4840];
        layer3[27][7:0] = buffer_data_1[4815:4808];
        layer3[27][15:8] = buffer_data_1[4823:4816];
        layer3[27][23:16] = buffer_data_1[4831:4824];
        layer3[27][31:24] = buffer_data_1[4839:4832];
        layer3[27][39:32] = buffer_data_1[4847:4840];
        layer4[27][7:0] = buffer_data_0[4815:4808];
        layer4[27][15:8] = buffer_data_0[4823:4816];
        layer4[27][23:16] = buffer_data_0[4831:4824];
        layer4[27][31:24] = buffer_data_0[4839:4832];
        layer4[27][39:32] = buffer_data_0[4847:4840];
        layer0[28][7:0] = buffer_data_4[4823:4816];
        layer0[28][15:8] = buffer_data_4[4831:4824];
        layer0[28][23:16] = buffer_data_4[4839:4832];
        layer0[28][31:24] = buffer_data_4[4847:4840];
        layer0[28][39:32] = buffer_data_4[4855:4848];
        layer1[28][7:0] = buffer_data_3[4823:4816];
        layer1[28][15:8] = buffer_data_3[4831:4824];
        layer1[28][23:16] = buffer_data_3[4839:4832];
        layer1[28][31:24] = buffer_data_3[4847:4840];
        layer1[28][39:32] = buffer_data_3[4855:4848];
        layer2[28][7:0] = buffer_data_2[4823:4816];
        layer2[28][15:8] = buffer_data_2[4831:4824];
        layer2[28][23:16] = buffer_data_2[4839:4832];
        layer2[28][31:24] = buffer_data_2[4847:4840];
        layer2[28][39:32] = buffer_data_2[4855:4848];
        layer3[28][7:0] = buffer_data_1[4823:4816];
        layer3[28][15:8] = buffer_data_1[4831:4824];
        layer3[28][23:16] = buffer_data_1[4839:4832];
        layer3[28][31:24] = buffer_data_1[4847:4840];
        layer3[28][39:32] = buffer_data_1[4855:4848];
        layer4[28][7:0] = buffer_data_0[4823:4816];
        layer4[28][15:8] = buffer_data_0[4831:4824];
        layer4[28][23:16] = buffer_data_0[4839:4832];
        layer4[28][31:24] = buffer_data_0[4847:4840];
        layer4[28][39:32] = buffer_data_0[4855:4848];
        layer0[29][7:0] = buffer_data_4[4831:4824];
        layer0[29][15:8] = buffer_data_4[4839:4832];
        layer0[29][23:16] = buffer_data_4[4847:4840];
        layer0[29][31:24] = buffer_data_4[4855:4848];
        layer0[29][39:32] = buffer_data_4[4863:4856];
        layer1[29][7:0] = buffer_data_3[4831:4824];
        layer1[29][15:8] = buffer_data_3[4839:4832];
        layer1[29][23:16] = buffer_data_3[4847:4840];
        layer1[29][31:24] = buffer_data_3[4855:4848];
        layer1[29][39:32] = buffer_data_3[4863:4856];
        layer2[29][7:0] = buffer_data_2[4831:4824];
        layer2[29][15:8] = buffer_data_2[4839:4832];
        layer2[29][23:16] = buffer_data_2[4847:4840];
        layer2[29][31:24] = buffer_data_2[4855:4848];
        layer2[29][39:32] = buffer_data_2[4863:4856];
        layer3[29][7:0] = buffer_data_1[4831:4824];
        layer3[29][15:8] = buffer_data_1[4839:4832];
        layer3[29][23:16] = buffer_data_1[4847:4840];
        layer3[29][31:24] = buffer_data_1[4855:4848];
        layer3[29][39:32] = buffer_data_1[4863:4856];
        layer4[29][7:0] = buffer_data_0[4831:4824];
        layer4[29][15:8] = buffer_data_0[4839:4832];
        layer4[29][23:16] = buffer_data_0[4847:4840];
        layer4[29][31:24] = buffer_data_0[4855:4848];
        layer4[29][39:32] = buffer_data_0[4863:4856];
        layer0[30][7:0] = buffer_data_4[4839:4832];
        layer0[30][15:8] = buffer_data_4[4847:4840];
        layer0[30][23:16] = buffer_data_4[4855:4848];
        layer0[30][31:24] = buffer_data_4[4863:4856];
        layer0[30][39:32] = buffer_data_4[4871:4864];
        layer1[30][7:0] = buffer_data_3[4839:4832];
        layer1[30][15:8] = buffer_data_3[4847:4840];
        layer1[30][23:16] = buffer_data_3[4855:4848];
        layer1[30][31:24] = buffer_data_3[4863:4856];
        layer1[30][39:32] = buffer_data_3[4871:4864];
        layer2[30][7:0] = buffer_data_2[4839:4832];
        layer2[30][15:8] = buffer_data_2[4847:4840];
        layer2[30][23:16] = buffer_data_2[4855:4848];
        layer2[30][31:24] = buffer_data_2[4863:4856];
        layer2[30][39:32] = buffer_data_2[4871:4864];
        layer3[30][7:0] = buffer_data_1[4839:4832];
        layer3[30][15:8] = buffer_data_1[4847:4840];
        layer3[30][23:16] = buffer_data_1[4855:4848];
        layer3[30][31:24] = buffer_data_1[4863:4856];
        layer3[30][39:32] = buffer_data_1[4871:4864];
        layer4[30][7:0] = buffer_data_0[4839:4832];
        layer4[30][15:8] = buffer_data_0[4847:4840];
        layer4[30][23:16] = buffer_data_0[4855:4848];
        layer4[30][31:24] = buffer_data_0[4863:4856];
        layer4[30][39:32] = buffer_data_0[4871:4864];
        layer0[31][7:0] = buffer_data_4[4847:4840];
        layer0[31][15:8] = buffer_data_4[4855:4848];
        layer0[31][23:16] = buffer_data_4[4863:4856];
        layer0[31][31:24] = buffer_data_4[4871:4864];
        layer0[31][39:32] = buffer_data_4[4879:4872];
        layer1[31][7:0] = buffer_data_3[4847:4840];
        layer1[31][15:8] = buffer_data_3[4855:4848];
        layer1[31][23:16] = buffer_data_3[4863:4856];
        layer1[31][31:24] = buffer_data_3[4871:4864];
        layer1[31][39:32] = buffer_data_3[4879:4872];
        layer2[31][7:0] = buffer_data_2[4847:4840];
        layer2[31][15:8] = buffer_data_2[4855:4848];
        layer2[31][23:16] = buffer_data_2[4863:4856];
        layer2[31][31:24] = buffer_data_2[4871:4864];
        layer2[31][39:32] = buffer_data_2[4879:4872];
        layer3[31][7:0] = buffer_data_1[4847:4840];
        layer3[31][15:8] = buffer_data_1[4855:4848];
        layer3[31][23:16] = buffer_data_1[4863:4856];
        layer3[31][31:24] = buffer_data_1[4871:4864];
        layer3[31][39:32] = buffer_data_1[4879:4872];
        layer4[31][7:0] = buffer_data_0[4847:4840];
        layer4[31][15:8] = buffer_data_0[4855:4848];
        layer4[31][23:16] = buffer_data_0[4863:4856];
        layer4[31][31:24] = buffer_data_0[4871:4864];
        layer4[31][39:32] = buffer_data_0[4879:4872];
        layer0[32][7:0] = buffer_data_4[4855:4848];
        layer0[32][15:8] = buffer_data_4[4863:4856];
        layer0[32][23:16] = buffer_data_4[4871:4864];
        layer0[32][31:24] = buffer_data_4[4879:4872];
        layer0[32][39:32] = buffer_data_4[4887:4880];
        layer1[32][7:0] = buffer_data_3[4855:4848];
        layer1[32][15:8] = buffer_data_3[4863:4856];
        layer1[32][23:16] = buffer_data_3[4871:4864];
        layer1[32][31:24] = buffer_data_3[4879:4872];
        layer1[32][39:32] = buffer_data_3[4887:4880];
        layer2[32][7:0] = buffer_data_2[4855:4848];
        layer2[32][15:8] = buffer_data_2[4863:4856];
        layer2[32][23:16] = buffer_data_2[4871:4864];
        layer2[32][31:24] = buffer_data_2[4879:4872];
        layer2[32][39:32] = buffer_data_2[4887:4880];
        layer3[32][7:0] = buffer_data_1[4855:4848];
        layer3[32][15:8] = buffer_data_1[4863:4856];
        layer3[32][23:16] = buffer_data_1[4871:4864];
        layer3[32][31:24] = buffer_data_1[4879:4872];
        layer3[32][39:32] = buffer_data_1[4887:4880];
        layer4[32][7:0] = buffer_data_0[4855:4848];
        layer4[32][15:8] = buffer_data_0[4863:4856];
        layer4[32][23:16] = buffer_data_0[4871:4864];
        layer4[32][31:24] = buffer_data_0[4879:4872];
        layer4[32][39:32] = buffer_data_0[4887:4880];
        layer0[33][7:0] = buffer_data_4[4863:4856];
        layer0[33][15:8] = buffer_data_4[4871:4864];
        layer0[33][23:16] = buffer_data_4[4879:4872];
        layer0[33][31:24] = buffer_data_4[4887:4880];
        layer0[33][39:32] = buffer_data_4[4895:4888];
        layer1[33][7:0] = buffer_data_3[4863:4856];
        layer1[33][15:8] = buffer_data_3[4871:4864];
        layer1[33][23:16] = buffer_data_3[4879:4872];
        layer1[33][31:24] = buffer_data_3[4887:4880];
        layer1[33][39:32] = buffer_data_3[4895:4888];
        layer2[33][7:0] = buffer_data_2[4863:4856];
        layer2[33][15:8] = buffer_data_2[4871:4864];
        layer2[33][23:16] = buffer_data_2[4879:4872];
        layer2[33][31:24] = buffer_data_2[4887:4880];
        layer2[33][39:32] = buffer_data_2[4895:4888];
        layer3[33][7:0] = buffer_data_1[4863:4856];
        layer3[33][15:8] = buffer_data_1[4871:4864];
        layer3[33][23:16] = buffer_data_1[4879:4872];
        layer3[33][31:24] = buffer_data_1[4887:4880];
        layer3[33][39:32] = buffer_data_1[4895:4888];
        layer4[33][7:0] = buffer_data_0[4863:4856];
        layer4[33][15:8] = buffer_data_0[4871:4864];
        layer4[33][23:16] = buffer_data_0[4879:4872];
        layer4[33][31:24] = buffer_data_0[4887:4880];
        layer4[33][39:32] = buffer_data_0[4895:4888];
        layer0[34][7:0] = buffer_data_4[4871:4864];
        layer0[34][15:8] = buffer_data_4[4879:4872];
        layer0[34][23:16] = buffer_data_4[4887:4880];
        layer0[34][31:24] = buffer_data_4[4895:4888];
        layer0[34][39:32] = buffer_data_4[4903:4896];
        layer1[34][7:0] = buffer_data_3[4871:4864];
        layer1[34][15:8] = buffer_data_3[4879:4872];
        layer1[34][23:16] = buffer_data_3[4887:4880];
        layer1[34][31:24] = buffer_data_3[4895:4888];
        layer1[34][39:32] = buffer_data_3[4903:4896];
        layer2[34][7:0] = buffer_data_2[4871:4864];
        layer2[34][15:8] = buffer_data_2[4879:4872];
        layer2[34][23:16] = buffer_data_2[4887:4880];
        layer2[34][31:24] = buffer_data_2[4895:4888];
        layer2[34][39:32] = buffer_data_2[4903:4896];
        layer3[34][7:0] = buffer_data_1[4871:4864];
        layer3[34][15:8] = buffer_data_1[4879:4872];
        layer3[34][23:16] = buffer_data_1[4887:4880];
        layer3[34][31:24] = buffer_data_1[4895:4888];
        layer3[34][39:32] = buffer_data_1[4903:4896];
        layer4[34][7:0] = buffer_data_0[4871:4864];
        layer4[34][15:8] = buffer_data_0[4879:4872];
        layer4[34][23:16] = buffer_data_0[4887:4880];
        layer4[34][31:24] = buffer_data_0[4895:4888];
        layer4[34][39:32] = buffer_data_0[4903:4896];
        layer0[35][7:0] = buffer_data_4[4879:4872];
        layer0[35][15:8] = buffer_data_4[4887:4880];
        layer0[35][23:16] = buffer_data_4[4895:4888];
        layer0[35][31:24] = buffer_data_4[4903:4896];
        layer0[35][39:32] = buffer_data_4[4911:4904];
        layer1[35][7:0] = buffer_data_3[4879:4872];
        layer1[35][15:8] = buffer_data_3[4887:4880];
        layer1[35][23:16] = buffer_data_3[4895:4888];
        layer1[35][31:24] = buffer_data_3[4903:4896];
        layer1[35][39:32] = buffer_data_3[4911:4904];
        layer2[35][7:0] = buffer_data_2[4879:4872];
        layer2[35][15:8] = buffer_data_2[4887:4880];
        layer2[35][23:16] = buffer_data_2[4895:4888];
        layer2[35][31:24] = buffer_data_2[4903:4896];
        layer2[35][39:32] = buffer_data_2[4911:4904];
        layer3[35][7:0] = buffer_data_1[4879:4872];
        layer3[35][15:8] = buffer_data_1[4887:4880];
        layer3[35][23:16] = buffer_data_1[4895:4888];
        layer3[35][31:24] = buffer_data_1[4903:4896];
        layer3[35][39:32] = buffer_data_1[4911:4904];
        layer4[35][7:0] = buffer_data_0[4879:4872];
        layer4[35][15:8] = buffer_data_0[4887:4880];
        layer4[35][23:16] = buffer_data_0[4895:4888];
        layer4[35][31:24] = buffer_data_0[4903:4896];
        layer4[35][39:32] = buffer_data_0[4911:4904];
        layer0[36][7:0] = buffer_data_4[4887:4880];
        layer0[36][15:8] = buffer_data_4[4895:4888];
        layer0[36][23:16] = buffer_data_4[4903:4896];
        layer0[36][31:24] = buffer_data_4[4911:4904];
        layer0[36][39:32] = buffer_data_4[4919:4912];
        layer1[36][7:0] = buffer_data_3[4887:4880];
        layer1[36][15:8] = buffer_data_3[4895:4888];
        layer1[36][23:16] = buffer_data_3[4903:4896];
        layer1[36][31:24] = buffer_data_3[4911:4904];
        layer1[36][39:32] = buffer_data_3[4919:4912];
        layer2[36][7:0] = buffer_data_2[4887:4880];
        layer2[36][15:8] = buffer_data_2[4895:4888];
        layer2[36][23:16] = buffer_data_2[4903:4896];
        layer2[36][31:24] = buffer_data_2[4911:4904];
        layer2[36][39:32] = buffer_data_2[4919:4912];
        layer3[36][7:0] = buffer_data_1[4887:4880];
        layer3[36][15:8] = buffer_data_1[4895:4888];
        layer3[36][23:16] = buffer_data_1[4903:4896];
        layer3[36][31:24] = buffer_data_1[4911:4904];
        layer3[36][39:32] = buffer_data_1[4919:4912];
        layer4[36][7:0] = buffer_data_0[4887:4880];
        layer4[36][15:8] = buffer_data_0[4895:4888];
        layer4[36][23:16] = buffer_data_0[4903:4896];
        layer4[36][31:24] = buffer_data_0[4911:4904];
        layer4[36][39:32] = buffer_data_0[4919:4912];
        layer0[37][7:0] = buffer_data_4[4895:4888];
        layer0[37][15:8] = buffer_data_4[4903:4896];
        layer0[37][23:16] = buffer_data_4[4911:4904];
        layer0[37][31:24] = buffer_data_4[4919:4912];
        layer0[37][39:32] = buffer_data_4[4927:4920];
        layer1[37][7:0] = buffer_data_3[4895:4888];
        layer1[37][15:8] = buffer_data_3[4903:4896];
        layer1[37][23:16] = buffer_data_3[4911:4904];
        layer1[37][31:24] = buffer_data_3[4919:4912];
        layer1[37][39:32] = buffer_data_3[4927:4920];
        layer2[37][7:0] = buffer_data_2[4895:4888];
        layer2[37][15:8] = buffer_data_2[4903:4896];
        layer2[37][23:16] = buffer_data_2[4911:4904];
        layer2[37][31:24] = buffer_data_2[4919:4912];
        layer2[37][39:32] = buffer_data_2[4927:4920];
        layer3[37][7:0] = buffer_data_1[4895:4888];
        layer3[37][15:8] = buffer_data_1[4903:4896];
        layer3[37][23:16] = buffer_data_1[4911:4904];
        layer3[37][31:24] = buffer_data_1[4919:4912];
        layer3[37][39:32] = buffer_data_1[4927:4920];
        layer4[37][7:0] = buffer_data_0[4895:4888];
        layer4[37][15:8] = buffer_data_0[4903:4896];
        layer4[37][23:16] = buffer_data_0[4911:4904];
        layer4[37][31:24] = buffer_data_0[4919:4912];
        layer4[37][39:32] = buffer_data_0[4927:4920];
        layer0[38][7:0] = buffer_data_4[4903:4896];
        layer0[38][15:8] = buffer_data_4[4911:4904];
        layer0[38][23:16] = buffer_data_4[4919:4912];
        layer0[38][31:24] = buffer_data_4[4927:4920];
        layer0[38][39:32] = buffer_data_4[4935:4928];
        layer1[38][7:0] = buffer_data_3[4903:4896];
        layer1[38][15:8] = buffer_data_3[4911:4904];
        layer1[38][23:16] = buffer_data_3[4919:4912];
        layer1[38][31:24] = buffer_data_3[4927:4920];
        layer1[38][39:32] = buffer_data_3[4935:4928];
        layer2[38][7:0] = buffer_data_2[4903:4896];
        layer2[38][15:8] = buffer_data_2[4911:4904];
        layer2[38][23:16] = buffer_data_2[4919:4912];
        layer2[38][31:24] = buffer_data_2[4927:4920];
        layer2[38][39:32] = buffer_data_2[4935:4928];
        layer3[38][7:0] = buffer_data_1[4903:4896];
        layer3[38][15:8] = buffer_data_1[4911:4904];
        layer3[38][23:16] = buffer_data_1[4919:4912];
        layer3[38][31:24] = buffer_data_1[4927:4920];
        layer3[38][39:32] = buffer_data_1[4935:4928];
        layer4[38][7:0] = buffer_data_0[4903:4896];
        layer4[38][15:8] = buffer_data_0[4911:4904];
        layer4[38][23:16] = buffer_data_0[4919:4912];
        layer4[38][31:24] = buffer_data_0[4927:4920];
        layer4[38][39:32] = buffer_data_0[4935:4928];
        layer0[39][7:0] = buffer_data_4[4911:4904];
        layer0[39][15:8] = buffer_data_4[4919:4912];
        layer0[39][23:16] = buffer_data_4[4927:4920];
        layer0[39][31:24] = buffer_data_4[4935:4928];
        layer0[39][39:32] = buffer_data_4[4943:4936];
        layer1[39][7:0] = buffer_data_3[4911:4904];
        layer1[39][15:8] = buffer_data_3[4919:4912];
        layer1[39][23:16] = buffer_data_3[4927:4920];
        layer1[39][31:24] = buffer_data_3[4935:4928];
        layer1[39][39:32] = buffer_data_3[4943:4936];
        layer2[39][7:0] = buffer_data_2[4911:4904];
        layer2[39][15:8] = buffer_data_2[4919:4912];
        layer2[39][23:16] = buffer_data_2[4927:4920];
        layer2[39][31:24] = buffer_data_2[4935:4928];
        layer2[39][39:32] = buffer_data_2[4943:4936];
        layer3[39][7:0] = buffer_data_1[4911:4904];
        layer3[39][15:8] = buffer_data_1[4919:4912];
        layer3[39][23:16] = buffer_data_1[4927:4920];
        layer3[39][31:24] = buffer_data_1[4935:4928];
        layer3[39][39:32] = buffer_data_1[4943:4936];
        layer4[39][7:0] = buffer_data_0[4911:4904];
        layer4[39][15:8] = buffer_data_0[4919:4912];
        layer4[39][23:16] = buffer_data_0[4927:4920];
        layer4[39][31:24] = buffer_data_0[4935:4928];
        layer4[39][39:32] = buffer_data_0[4943:4936];
        layer0[40][7:0] = buffer_data_4[4919:4912];
        layer0[40][15:8] = buffer_data_4[4927:4920];
        layer0[40][23:16] = buffer_data_4[4935:4928];
        layer0[40][31:24] = buffer_data_4[4943:4936];
        layer0[40][39:32] = buffer_data_4[4951:4944];
        layer1[40][7:0] = buffer_data_3[4919:4912];
        layer1[40][15:8] = buffer_data_3[4927:4920];
        layer1[40][23:16] = buffer_data_3[4935:4928];
        layer1[40][31:24] = buffer_data_3[4943:4936];
        layer1[40][39:32] = buffer_data_3[4951:4944];
        layer2[40][7:0] = buffer_data_2[4919:4912];
        layer2[40][15:8] = buffer_data_2[4927:4920];
        layer2[40][23:16] = buffer_data_2[4935:4928];
        layer2[40][31:24] = buffer_data_2[4943:4936];
        layer2[40][39:32] = buffer_data_2[4951:4944];
        layer3[40][7:0] = buffer_data_1[4919:4912];
        layer3[40][15:8] = buffer_data_1[4927:4920];
        layer3[40][23:16] = buffer_data_1[4935:4928];
        layer3[40][31:24] = buffer_data_1[4943:4936];
        layer3[40][39:32] = buffer_data_1[4951:4944];
        layer4[40][7:0] = buffer_data_0[4919:4912];
        layer4[40][15:8] = buffer_data_0[4927:4920];
        layer4[40][23:16] = buffer_data_0[4935:4928];
        layer4[40][31:24] = buffer_data_0[4943:4936];
        layer4[40][39:32] = buffer_data_0[4951:4944];
        layer0[41][7:0] = buffer_data_4[4927:4920];
        layer0[41][15:8] = buffer_data_4[4935:4928];
        layer0[41][23:16] = buffer_data_4[4943:4936];
        layer0[41][31:24] = buffer_data_4[4951:4944];
        layer0[41][39:32] = buffer_data_4[4959:4952];
        layer1[41][7:0] = buffer_data_3[4927:4920];
        layer1[41][15:8] = buffer_data_3[4935:4928];
        layer1[41][23:16] = buffer_data_3[4943:4936];
        layer1[41][31:24] = buffer_data_3[4951:4944];
        layer1[41][39:32] = buffer_data_3[4959:4952];
        layer2[41][7:0] = buffer_data_2[4927:4920];
        layer2[41][15:8] = buffer_data_2[4935:4928];
        layer2[41][23:16] = buffer_data_2[4943:4936];
        layer2[41][31:24] = buffer_data_2[4951:4944];
        layer2[41][39:32] = buffer_data_2[4959:4952];
        layer3[41][7:0] = buffer_data_1[4927:4920];
        layer3[41][15:8] = buffer_data_1[4935:4928];
        layer3[41][23:16] = buffer_data_1[4943:4936];
        layer3[41][31:24] = buffer_data_1[4951:4944];
        layer3[41][39:32] = buffer_data_1[4959:4952];
        layer4[41][7:0] = buffer_data_0[4927:4920];
        layer4[41][15:8] = buffer_data_0[4935:4928];
        layer4[41][23:16] = buffer_data_0[4943:4936];
        layer4[41][31:24] = buffer_data_0[4951:4944];
        layer4[41][39:32] = buffer_data_0[4959:4952];
        layer0[42][7:0] = buffer_data_4[4935:4928];
        layer0[42][15:8] = buffer_data_4[4943:4936];
        layer0[42][23:16] = buffer_data_4[4951:4944];
        layer0[42][31:24] = buffer_data_4[4959:4952];
        layer0[42][39:32] = buffer_data_4[4967:4960];
        layer1[42][7:0] = buffer_data_3[4935:4928];
        layer1[42][15:8] = buffer_data_3[4943:4936];
        layer1[42][23:16] = buffer_data_3[4951:4944];
        layer1[42][31:24] = buffer_data_3[4959:4952];
        layer1[42][39:32] = buffer_data_3[4967:4960];
        layer2[42][7:0] = buffer_data_2[4935:4928];
        layer2[42][15:8] = buffer_data_2[4943:4936];
        layer2[42][23:16] = buffer_data_2[4951:4944];
        layer2[42][31:24] = buffer_data_2[4959:4952];
        layer2[42][39:32] = buffer_data_2[4967:4960];
        layer3[42][7:0] = buffer_data_1[4935:4928];
        layer3[42][15:8] = buffer_data_1[4943:4936];
        layer3[42][23:16] = buffer_data_1[4951:4944];
        layer3[42][31:24] = buffer_data_1[4959:4952];
        layer3[42][39:32] = buffer_data_1[4967:4960];
        layer4[42][7:0] = buffer_data_0[4935:4928];
        layer4[42][15:8] = buffer_data_0[4943:4936];
        layer4[42][23:16] = buffer_data_0[4951:4944];
        layer4[42][31:24] = buffer_data_0[4959:4952];
        layer4[42][39:32] = buffer_data_0[4967:4960];
        layer0[43][7:0] = buffer_data_4[4943:4936];
        layer0[43][15:8] = buffer_data_4[4951:4944];
        layer0[43][23:16] = buffer_data_4[4959:4952];
        layer0[43][31:24] = buffer_data_4[4967:4960];
        layer0[43][39:32] = buffer_data_4[4975:4968];
        layer1[43][7:0] = buffer_data_3[4943:4936];
        layer1[43][15:8] = buffer_data_3[4951:4944];
        layer1[43][23:16] = buffer_data_3[4959:4952];
        layer1[43][31:24] = buffer_data_3[4967:4960];
        layer1[43][39:32] = buffer_data_3[4975:4968];
        layer2[43][7:0] = buffer_data_2[4943:4936];
        layer2[43][15:8] = buffer_data_2[4951:4944];
        layer2[43][23:16] = buffer_data_2[4959:4952];
        layer2[43][31:24] = buffer_data_2[4967:4960];
        layer2[43][39:32] = buffer_data_2[4975:4968];
        layer3[43][7:0] = buffer_data_1[4943:4936];
        layer3[43][15:8] = buffer_data_1[4951:4944];
        layer3[43][23:16] = buffer_data_1[4959:4952];
        layer3[43][31:24] = buffer_data_1[4967:4960];
        layer3[43][39:32] = buffer_data_1[4975:4968];
        layer4[43][7:0] = buffer_data_0[4943:4936];
        layer4[43][15:8] = buffer_data_0[4951:4944];
        layer4[43][23:16] = buffer_data_0[4959:4952];
        layer4[43][31:24] = buffer_data_0[4967:4960];
        layer4[43][39:32] = buffer_data_0[4975:4968];
        layer0[44][7:0] = buffer_data_4[4951:4944];
        layer0[44][15:8] = buffer_data_4[4959:4952];
        layer0[44][23:16] = buffer_data_4[4967:4960];
        layer0[44][31:24] = buffer_data_4[4975:4968];
        layer0[44][39:32] = buffer_data_4[4983:4976];
        layer1[44][7:0] = buffer_data_3[4951:4944];
        layer1[44][15:8] = buffer_data_3[4959:4952];
        layer1[44][23:16] = buffer_data_3[4967:4960];
        layer1[44][31:24] = buffer_data_3[4975:4968];
        layer1[44][39:32] = buffer_data_3[4983:4976];
        layer2[44][7:0] = buffer_data_2[4951:4944];
        layer2[44][15:8] = buffer_data_2[4959:4952];
        layer2[44][23:16] = buffer_data_2[4967:4960];
        layer2[44][31:24] = buffer_data_2[4975:4968];
        layer2[44][39:32] = buffer_data_2[4983:4976];
        layer3[44][7:0] = buffer_data_1[4951:4944];
        layer3[44][15:8] = buffer_data_1[4959:4952];
        layer3[44][23:16] = buffer_data_1[4967:4960];
        layer3[44][31:24] = buffer_data_1[4975:4968];
        layer3[44][39:32] = buffer_data_1[4983:4976];
        layer4[44][7:0] = buffer_data_0[4951:4944];
        layer4[44][15:8] = buffer_data_0[4959:4952];
        layer4[44][23:16] = buffer_data_0[4967:4960];
        layer4[44][31:24] = buffer_data_0[4975:4968];
        layer4[44][39:32] = buffer_data_0[4983:4976];
        layer0[45][7:0] = buffer_data_4[4959:4952];
        layer0[45][15:8] = buffer_data_4[4967:4960];
        layer0[45][23:16] = buffer_data_4[4975:4968];
        layer0[45][31:24] = buffer_data_4[4983:4976];
        layer0[45][39:32] = buffer_data_4[4991:4984];
        layer1[45][7:0] = buffer_data_3[4959:4952];
        layer1[45][15:8] = buffer_data_3[4967:4960];
        layer1[45][23:16] = buffer_data_3[4975:4968];
        layer1[45][31:24] = buffer_data_3[4983:4976];
        layer1[45][39:32] = buffer_data_3[4991:4984];
        layer2[45][7:0] = buffer_data_2[4959:4952];
        layer2[45][15:8] = buffer_data_2[4967:4960];
        layer2[45][23:16] = buffer_data_2[4975:4968];
        layer2[45][31:24] = buffer_data_2[4983:4976];
        layer2[45][39:32] = buffer_data_2[4991:4984];
        layer3[45][7:0] = buffer_data_1[4959:4952];
        layer3[45][15:8] = buffer_data_1[4967:4960];
        layer3[45][23:16] = buffer_data_1[4975:4968];
        layer3[45][31:24] = buffer_data_1[4983:4976];
        layer3[45][39:32] = buffer_data_1[4991:4984];
        layer4[45][7:0] = buffer_data_0[4959:4952];
        layer4[45][15:8] = buffer_data_0[4967:4960];
        layer4[45][23:16] = buffer_data_0[4975:4968];
        layer4[45][31:24] = buffer_data_0[4983:4976];
        layer4[45][39:32] = buffer_data_0[4991:4984];
        layer0[46][7:0] = buffer_data_4[4967:4960];
        layer0[46][15:8] = buffer_data_4[4975:4968];
        layer0[46][23:16] = buffer_data_4[4983:4976];
        layer0[46][31:24] = buffer_data_4[4991:4984];
        layer0[46][39:32] = buffer_data_4[4999:4992];
        layer1[46][7:0] = buffer_data_3[4967:4960];
        layer1[46][15:8] = buffer_data_3[4975:4968];
        layer1[46][23:16] = buffer_data_3[4983:4976];
        layer1[46][31:24] = buffer_data_3[4991:4984];
        layer1[46][39:32] = buffer_data_3[4999:4992];
        layer2[46][7:0] = buffer_data_2[4967:4960];
        layer2[46][15:8] = buffer_data_2[4975:4968];
        layer2[46][23:16] = buffer_data_2[4983:4976];
        layer2[46][31:24] = buffer_data_2[4991:4984];
        layer2[46][39:32] = buffer_data_2[4999:4992];
        layer3[46][7:0] = buffer_data_1[4967:4960];
        layer3[46][15:8] = buffer_data_1[4975:4968];
        layer3[46][23:16] = buffer_data_1[4983:4976];
        layer3[46][31:24] = buffer_data_1[4991:4984];
        layer3[46][39:32] = buffer_data_1[4999:4992];
        layer4[46][7:0] = buffer_data_0[4967:4960];
        layer4[46][15:8] = buffer_data_0[4975:4968];
        layer4[46][23:16] = buffer_data_0[4983:4976];
        layer4[46][31:24] = buffer_data_0[4991:4984];
        layer4[46][39:32] = buffer_data_0[4999:4992];
        layer0[47][7:0] = buffer_data_4[4975:4968];
        layer0[47][15:8] = buffer_data_4[4983:4976];
        layer0[47][23:16] = buffer_data_4[4991:4984];
        layer0[47][31:24] = buffer_data_4[4999:4992];
        layer0[47][39:32] = buffer_data_4[5007:5000];
        layer1[47][7:0] = buffer_data_3[4975:4968];
        layer1[47][15:8] = buffer_data_3[4983:4976];
        layer1[47][23:16] = buffer_data_3[4991:4984];
        layer1[47][31:24] = buffer_data_3[4999:4992];
        layer1[47][39:32] = buffer_data_3[5007:5000];
        layer2[47][7:0] = buffer_data_2[4975:4968];
        layer2[47][15:8] = buffer_data_2[4983:4976];
        layer2[47][23:16] = buffer_data_2[4991:4984];
        layer2[47][31:24] = buffer_data_2[4999:4992];
        layer2[47][39:32] = buffer_data_2[5007:5000];
        layer3[47][7:0] = buffer_data_1[4975:4968];
        layer3[47][15:8] = buffer_data_1[4983:4976];
        layer3[47][23:16] = buffer_data_1[4991:4984];
        layer3[47][31:24] = buffer_data_1[4999:4992];
        layer3[47][39:32] = buffer_data_1[5007:5000];
        layer4[47][7:0] = buffer_data_0[4975:4968];
        layer4[47][15:8] = buffer_data_0[4983:4976];
        layer4[47][23:16] = buffer_data_0[4991:4984];
        layer4[47][31:24] = buffer_data_0[4999:4992];
        layer4[47][39:32] = buffer_data_0[5007:5000];
        layer0[48][7:0] = buffer_data_4[4983:4976];
        layer0[48][15:8] = buffer_data_4[4991:4984];
        layer0[48][23:16] = buffer_data_4[4999:4992];
        layer0[48][31:24] = buffer_data_4[5007:5000];
        layer0[48][39:32] = buffer_data_4[5015:5008];
        layer1[48][7:0] = buffer_data_3[4983:4976];
        layer1[48][15:8] = buffer_data_3[4991:4984];
        layer1[48][23:16] = buffer_data_3[4999:4992];
        layer1[48][31:24] = buffer_data_3[5007:5000];
        layer1[48][39:32] = buffer_data_3[5015:5008];
        layer2[48][7:0] = buffer_data_2[4983:4976];
        layer2[48][15:8] = buffer_data_2[4991:4984];
        layer2[48][23:16] = buffer_data_2[4999:4992];
        layer2[48][31:24] = buffer_data_2[5007:5000];
        layer2[48][39:32] = buffer_data_2[5015:5008];
        layer3[48][7:0] = buffer_data_1[4983:4976];
        layer3[48][15:8] = buffer_data_1[4991:4984];
        layer3[48][23:16] = buffer_data_1[4999:4992];
        layer3[48][31:24] = buffer_data_1[5007:5000];
        layer3[48][39:32] = buffer_data_1[5015:5008];
        layer4[48][7:0] = buffer_data_0[4983:4976];
        layer4[48][15:8] = buffer_data_0[4991:4984];
        layer4[48][23:16] = buffer_data_0[4999:4992];
        layer4[48][31:24] = buffer_data_0[5007:5000];
        layer4[48][39:32] = buffer_data_0[5015:5008];
        layer0[49][7:0] = buffer_data_4[4991:4984];
        layer0[49][15:8] = buffer_data_4[4999:4992];
        layer0[49][23:16] = buffer_data_4[5007:5000];
        layer0[49][31:24] = buffer_data_4[5015:5008];
        layer0[49][39:32] = buffer_data_4[5023:5016];
        layer1[49][7:0] = buffer_data_3[4991:4984];
        layer1[49][15:8] = buffer_data_3[4999:4992];
        layer1[49][23:16] = buffer_data_3[5007:5000];
        layer1[49][31:24] = buffer_data_3[5015:5008];
        layer1[49][39:32] = buffer_data_3[5023:5016];
        layer2[49][7:0] = buffer_data_2[4991:4984];
        layer2[49][15:8] = buffer_data_2[4999:4992];
        layer2[49][23:16] = buffer_data_2[5007:5000];
        layer2[49][31:24] = buffer_data_2[5015:5008];
        layer2[49][39:32] = buffer_data_2[5023:5016];
        layer3[49][7:0] = buffer_data_1[4991:4984];
        layer3[49][15:8] = buffer_data_1[4999:4992];
        layer3[49][23:16] = buffer_data_1[5007:5000];
        layer3[49][31:24] = buffer_data_1[5015:5008];
        layer3[49][39:32] = buffer_data_1[5023:5016];
        layer4[49][7:0] = buffer_data_0[4991:4984];
        layer4[49][15:8] = buffer_data_0[4999:4992];
        layer4[49][23:16] = buffer_data_0[5007:5000];
        layer4[49][31:24] = buffer_data_0[5015:5008];
        layer4[49][39:32] = buffer_data_0[5023:5016];
        layer0[50][7:0] = buffer_data_4[4999:4992];
        layer0[50][15:8] = buffer_data_4[5007:5000];
        layer0[50][23:16] = buffer_data_4[5015:5008];
        layer0[50][31:24] = buffer_data_4[5023:5016];
        layer0[50][39:32] = buffer_data_4[5031:5024];
        layer1[50][7:0] = buffer_data_3[4999:4992];
        layer1[50][15:8] = buffer_data_3[5007:5000];
        layer1[50][23:16] = buffer_data_3[5015:5008];
        layer1[50][31:24] = buffer_data_3[5023:5016];
        layer1[50][39:32] = buffer_data_3[5031:5024];
        layer2[50][7:0] = buffer_data_2[4999:4992];
        layer2[50][15:8] = buffer_data_2[5007:5000];
        layer2[50][23:16] = buffer_data_2[5015:5008];
        layer2[50][31:24] = buffer_data_2[5023:5016];
        layer2[50][39:32] = buffer_data_2[5031:5024];
        layer3[50][7:0] = buffer_data_1[4999:4992];
        layer3[50][15:8] = buffer_data_1[5007:5000];
        layer3[50][23:16] = buffer_data_1[5015:5008];
        layer3[50][31:24] = buffer_data_1[5023:5016];
        layer3[50][39:32] = buffer_data_1[5031:5024];
        layer4[50][7:0] = buffer_data_0[4999:4992];
        layer4[50][15:8] = buffer_data_0[5007:5000];
        layer4[50][23:16] = buffer_data_0[5015:5008];
        layer4[50][31:24] = buffer_data_0[5023:5016];
        layer4[50][39:32] = buffer_data_0[5031:5024];
        layer0[51][7:0] = buffer_data_4[5007:5000];
        layer0[51][15:8] = buffer_data_4[5015:5008];
        layer0[51][23:16] = buffer_data_4[5023:5016];
        layer0[51][31:24] = buffer_data_4[5031:5024];
        layer0[51][39:32] = buffer_data_4[5039:5032];
        layer1[51][7:0] = buffer_data_3[5007:5000];
        layer1[51][15:8] = buffer_data_3[5015:5008];
        layer1[51][23:16] = buffer_data_3[5023:5016];
        layer1[51][31:24] = buffer_data_3[5031:5024];
        layer1[51][39:32] = buffer_data_3[5039:5032];
        layer2[51][7:0] = buffer_data_2[5007:5000];
        layer2[51][15:8] = buffer_data_2[5015:5008];
        layer2[51][23:16] = buffer_data_2[5023:5016];
        layer2[51][31:24] = buffer_data_2[5031:5024];
        layer2[51][39:32] = buffer_data_2[5039:5032];
        layer3[51][7:0] = buffer_data_1[5007:5000];
        layer3[51][15:8] = buffer_data_1[5015:5008];
        layer3[51][23:16] = buffer_data_1[5023:5016];
        layer3[51][31:24] = buffer_data_1[5031:5024];
        layer3[51][39:32] = buffer_data_1[5039:5032];
        layer4[51][7:0] = buffer_data_0[5007:5000];
        layer4[51][15:8] = buffer_data_0[5015:5008];
        layer4[51][23:16] = buffer_data_0[5023:5016];
        layer4[51][31:24] = buffer_data_0[5031:5024];
        layer4[51][39:32] = buffer_data_0[5039:5032];
        layer0[52][7:0] = buffer_data_4[5015:5008];
        layer0[52][15:8] = buffer_data_4[5023:5016];
        layer0[52][23:16] = buffer_data_4[5031:5024];
        layer0[52][31:24] = buffer_data_4[5039:5032];
        layer0[52][39:32] = buffer_data_4[5047:5040];
        layer1[52][7:0] = buffer_data_3[5015:5008];
        layer1[52][15:8] = buffer_data_3[5023:5016];
        layer1[52][23:16] = buffer_data_3[5031:5024];
        layer1[52][31:24] = buffer_data_3[5039:5032];
        layer1[52][39:32] = buffer_data_3[5047:5040];
        layer2[52][7:0] = buffer_data_2[5015:5008];
        layer2[52][15:8] = buffer_data_2[5023:5016];
        layer2[52][23:16] = buffer_data_2[5031:5024];
        layer2[52][31:24] = buffer_data_2[5039:5032];
        layer2[52][39:32] = buffer_data_2[5047:5040];
        layer3[52][7:0] = buffer_data_1[5015:5008];
        layer3[52][15:8] = buffer_data_1[5023:5016];
        layer3[52][23:16] = buffer_data_1[5031:5024];
        layer3[52][31:24] = buffer_data_1[5039:5032];
        layer3[52][39:32] = buffer_data_1[5047:5040];
        layer4[52][7:0] = buffer_data_0[5015:5008];
        layer4[52][15:8] = buffer_data_0[5023:5016];
        layer4[52][23:16] = buffer_data_0[5031:5024];
        layer4[52][31:24] = buffer_data_0[5039:5032];
        layer4[52][39:32] = buffer_data_0[5047:5040];
        layer0[53][7:0] = buffer_data_4[5023:5016];
        layer0[53][15:8] = buffer_data_4[5031:5024];
        layer0[53][23:16] = buffer_data_4[5039:5032];
        layer0[53][31:24] = buffer_data_4[5047:5040];
        layer0[53][39:32] = buffer_data_4[5055:5048];
        layer1[53][7:0] = buffer_data_3[5023:5016];
        layer1[53][15:8] = buffer_data_3[5031:5024];
        layer1[53][23:16] = buffer_data_3[5039:5032];
        layer1[53][31:24] = buffer_data_3[5047:5040];
        layer1[53][39:32] = buffer_data_3[5055:5048];
        layer2[53][7:0] = buffer_data_2[5023:5016];
        layer2[53][15:8] = buffer_data_2[5031:5024];
        layer2[53][23:16] = buffer_data_2[5039:5032];
        layer2[53][31:24] = buffer_data_2[5047:5040];
        layer2[53][39:32] = buffer_data_2[5055:5048];
        layer3[53][7:0] = buffer_data_1[5023:5016];
        layer3[53][15:8] = buffer_data_1[5031:5024];
        layer3[53][23:16] = buffer_data_1[5039:5032];
        layer3[53][31:24] = buffer_data_1[5047:5040];
        layer3[53][39:32] = buffer_data_1[5055:5048];
        layer4[53][7:0] = buffer_data_0[5023:5016];
        layer4[53][15:8] = buffer_data_0[5031:5024];
        layer4[53][23:16] = buffer_data_0[5039:5032];
        layer4[53][31:24] = buffer_data_0[5047:5040];
        layer4[53][39:32] = buffer_data_0[5055:5048];
        layer0[54][7:0] = buffer_data_4[5031:5024];
        layer0[54][15:8] = buffer_data_4[5039:5032];
        layer0[54][23:16] = buffer_data_4[5047:5040];
        layer0[54][31:24] = buffer_data_4[5055:5048];
        layer0[54][39:32] = buffer_data_4[5063:5056];
        layer1[54][7:0] = buffer_data_3[5031:5024];
        layer1[54][15:8] = buffer_data_3[5039:5032];
        layer1[54][23:16] = buffer_data_3[5047:5040];
        layer1[54][31:24] = buffer_data_3[5055:5048];
        layer1[54][39:32] = buffer_data_3[5063:5056];
        layer2[54][7:0] = buffer_data_2[5031:5024];
        layer2[54][15:8] = buffer_data_2[5039:5032];
        layer2[54][23:16] = buffer_data_2[5047:5040];
        layer2[54][31:24] = buffer_data_2[5055:5048];
        layer2[54][39:32] = buffer_data_2[5063:5056];
        layer3[54][7:0] = buffer_data_1[5031:5024];
        layer3[54][15:8] = buffer_data_1[5039:5032];
        layer3[54][23:16] = buffer_data_1[5047:5040];
        layer3[54][31:24] = buffer_data_1[5055:5048];
        layer3[54][39:32] = buffer_data_1[5063:5056];
        layer4[54][7:0] = buffer_data_0[5031:5024];
        layer4[54][15:8] = buffer_data_0[5039:5032];
        layer4[54][23:16] = buffer_data_0[5047:5040];
        layer4[54][31:24] = buffer_data_0[5055:5048];
        layer4[54][39:32] = buffer_data_0[5063:5056];
        layer0[55][7:0] = buffer_data_4[5039:5032];
        layer0[55][15:8] = buffer_data_4[5047:5040];
        layer0[55][23:16] = buffer_data_4[5055:5048];
        layer0[55][31:24] = buffer_data_4[5063:5056];
        layer0[55][39:32] = buffer_data_4[5071:5064];
        layer1[55][7:0] = buffer_data_3[5039:5032];
        layer1[55][15:8] = buffer_data_3[5047:5040];
        layer1[55][23:16] = buffer_data_3[5055:5048];
        layer1[55][31:24] = buffer_data_3[5063:5056];
        layer1[55][39:32] = buffer_data_3[5071:5064];
        layer2[55][7:0] = buffer_data_2[5039:5032];
        layer2[55][15:8] = buffer_data_2[5047:5040];
        layer2[55][23:16] = buffer_data_2[5055:5048];
        layer2[55][31:24] = buffer_data_2[5063:5056];
        layer2[55][39:32] = buffer_data_2[5071:5064];
        layer3[55][7:0] = buffer_data_1[5039:5032];
        layer3[55][15:8] = buffer_data_1[5047:5040];
        layer3[55][23:16] = buffer_data_1[5055:5048];
        layer3[55][31:24] = buffer_data_1[5063:5056];
        layer3[55][39:32] = buffer_data_1[5071:5064];
        layer4[55][7:0] = buffer_data_0[5039:5032];
        layer4[55][15:8] = buffer_data_0[5047:5040];
        layer4[55][23:16] = buffer_data_0[5055:5048];
        layer4[55][31:24] = buffer_data_0[5063:5056];
        layer4[55][39:32] = buffer_data_0[5071:5064];
        layer0[56][7:0] = buffer_data_4[5047:5040];
        layer0[56][15:8] = buffer_data_4[5055:5048];
        layer0[56][23:16] = buffer_data_4[5063:5056];
        layer0[56][31:24] = buffer_data_4[5071:5064];
        layer0[56][39:32] = buffer_data_4[5079:5072];
        layer1[56][7:0] = buffer_data_3[5047:5040];
        layer1[56][15:8] = buffer_data_3[5055:5048];
        layer1[56][23:16] = buffer_data_3[5063:5056];
        layer1[56][31:24] = buffer_data_3[5071:5064];
        layer1[56][39:32] = buffer_data_3[5079:5072];
        layer2[56][7:0] = buffer_data_2[5047:5040];
        layer2[56][15:8] = buffer_data_2[5055:5048];
        layer2[56][23:16] = buffer_data_2[5063:5056];
        layer2[56][31:24] = buffer_data_2[5071:5064];
        layer2[56][39:32] = buffer_data_2[5079:5072];
        layer3[56][7:0] = buffer_data_1[5047:5040];
        layer3[56][15:8] = buffer_data_1[5055:5048];
        layer3[56][23:16] = buffer_data_1[5063:5056];
        layer3[56][31:24] = buffer_data_1[5071:5064];
        layer3[56][39:32] = buffer_data_1[5079:5072];
        layer4[56][7:0] = buffer_data_0[5047:5040];
        layer4[56][15:8] = buffer_data_0[5055:5048];
        layer4[56][23:16] = buffer_data_0[5063:5056];
        layer4[56][31:24] = buffer_data_0[5071:5064];
        layer4[56][39:32] = buffer_data_0[5079:5072];
        layer0[57][7:0] = buffer_data_4[5055:5048];
        layer0[57][15:8] = buffer_data_4[5063:5056];
        layer0[57][23:16] = buffer_data_4[5071:5064];
        layer0[57][31:24] = buffer_data_4[5079:5072];
        layer0[57][39:32] = buffer_data_4[5087:5080];
        layer1[57][7:0] = buffer_data_3[5055:5048];
        layer1[57][15:8] = buffer_data_3[5063:5056];
        layer1[57][23:16] = buffer_data_3[5071:5064];
        layer1[57][31:24] = buffer_data_3[5079:5072];
        layer1[57][39:32] = buffer_data_3[5087:5080];
        layer2[57][7:0] = buffer_data_2[5055:5048];
        layer2[57][15:8] = buffer_data_2[5063:5056];
        layer2[57][23:16] = buffer_data_2[5071:5064];
        layer2[57][31:24] = buffer_data_2[5079:5072];
        layer2[57][39:32] = buffer_data_2[5087:5080];
        layer3[57][7:0] = buffer_data_1[5055:5048];
        layer3[57][15:8] = buffer_data_1[5063:5056];
        layer3[57][23:16] = buffer_data_1[5071:5064];
        layer3[57][31:24] = buffer_data_1[5079:5072];
        layer3[57][39:32] = buffer_data_1[5087:5080];
        layer4[57][7:0] = buffer_data_0[5055:5048];
        layer4[57][15:8] = buffer_data_0[5063:5056];
        layer4[57][23:16] = buffer_data_0[5071:5064];
        layer4[57][31:24] = buffer_data_0[5079:5072];
        layer4[57][39:32] = buffer_data_0[5087:5080];
        layer0[58][7:0] = buffer_data_4[5063:5056];
        layer0[58][15:8] = buffer_data_4[5071:5064];
        layer0[58][23:16] = buffer_data_4[5079:5072];
        layer0[58][31:24] = buffer_data_4[5087:5080];
        layer0[58][39:32] = buffer_data_4[5095:5088];
        layer1[58][7:0] = buffer_data_3[5063:5056];
        layer1[58][15:8] = buffer_data_3[5071:5064];
        layer1[58][23:16] = buffer_data_3[5079:5072];
        layer1[58][31:24] = buffer_data_3[5087:5080];
        layer1[58][39:32] = buffer_data_3[5095:5088];
        layer2[58][7:0] = buffer_data_2[5063:5056];
        layer2[58][15:8] = buffer_data_2[5071:5064];
        layer2[58][23:16] = buffer_data_2[5079:5072];
        layer2[58][31:24] = buffer_data_2[5087:5080];
        layer2[58][39:32] = buffer_data_2[5095:5088];
        layer3[58][7:0] = buffer_data_1[5063:5056];
        layer3[58][15:8] = buffer_data_1[5071:5064];
        layer3[58][23:16] = buffer_data_1[5079:5072];
        layer3[58][31:24] = buffer_data_1[5087:5080];
        layer3[58][39:32] = buffer_data_1[5095:5088];
        layer4[58][7:0] = buffer_data_0[5063:5056];
        layer4[58][15:8] = buffer_data_0[5071:5064];
        layer4[58][23:16] = buffer_data_0[5079:5072];
        layer4[58][31:24] = buffer_data_0[5087:5080];
        layer4[58][39:32] = buffer_data_0[5095:5088];
        layer0[59][7:0] = buffer_data_4[5071:5064];
        layer0[59][15:8] = buffer_data_4[5079:5072];
        layer0[59][23:16] = buffer_data_4[5087:5080];
        layer0[59][31:24] = buffer_data_4[5095:5088];
        layer0[59][39:32] = buffer_data_4[5103:5096];
        layer1[59][7:0] = buffer_data_3[5071:5064];
        layer1[59][15:8] = buffer_data_3[5079:5072];
        layer1[59][23:16] = buffer_data_3[5087:5080];
        layer1[59][31:24] = buffer_data_3[5095:5088];
        layer1[59][39:32] = buffer_data_3[5103:5096];
        layer2[59][7:0] = buffer_data_2[5071:5064];
        layer2[59][15:8] = buffer_data_2[5079:5072];
        layer2[59][23:16] = buffer_data_2[5087:5080];
        layer2[59][31:24] = buffer_data_2[5095:5088];
        layer2[59][39:32] = buffer_data_2[5103:5096];
        layer3[59][7:0] = buffer_data_1[5071:5064];
        layer3[59][15:8] = buffer_data_1[5079:5072];
        layer3[59][23:16] = buffer_data_1[5087:5080];
        layer3[59][31:24] = buffer_data_1[5095:5088];
        layer3[59][39:32] = buffer_data_1[5103:5096];
        layer4[59][7:0] = buffer_data_0[5071:5064];
        layer4[59][15:8] = buffer_data_0[5079:5072];
        layer4[59][23:16] = buffer_data_0[5087:5080];
        layer4[59][31:24] = buffer_data_0[5095:5088];
        layer4[59][39:32] = buffer_data_0[5103:5096];
        layer0[60][7:0] = buffer_data_4[5079:5072];
        layer0[60][15:8] = buffer_data_4[5087:5080];
        layer0[60][23:16] = buffer_data_4[5095:5088];
        layer0[60][31:24] = buffer_data_4[5103:5096];
        layer0[60][39:32] = buffer_data_4[5111:5104];
        layer1[60][7:0] = buffer_data_3[5079:5072];
        layer1[60][15:8] = buffer_data_3[5087:5080];
        layer1[60][23:16] = buffer_data_3[5095:5088];
        layer1[60][31:24] = buffer_data_3[5103:5096];
        layer1[60][39:32] = buffer_data_3[5111:5104];
        layer2[60][7:0] = buffer_data_2[5079:5072];
        layer2[60][15:8] = buffer_data_2[5087:5080];
        layer2[60][23:16] = buffer_data_2[5095:5088];
        layer2[60][31:24] = buffer_data_2[5103:5096];
        layer2[60][39:32] = buffer_data_2[5111:5104];
        layer3[60][7:0] = buffer_data_1[5079:5072];
        layer3[60][15:8] = buffer_data_1[5087:5080];
        layer3[60][23:16] = buffer_data_1[5095:5088];
        layer3[60][31:24] = buffer_data_1[5103:5096];
        layer3[60][39:32] = buffer_data_1[5111:5104];
        layer4[60][7:0] = buffer_data_0[5079:5072];
        layer4[60][15:8] = buffer_data_0[5087:5080];
        layer4[60][23:16] = buffer_data_0[5095:5088];
        layer4[60][31:24] = buffer_data_0[5103:5096];
        layer4[60][39:32] = buffer_data_0[5111:5104];
        layer0[61][7:0] = buffer_data_4[5087:5080];
        layer0[61][15:8] = buffer_data_4[5095:5088];
        layer0[61][23:16] = buffer_data_4[5103:5096];
        layer0[61][31:24] = buffer_data_4[5111:5104];
        layer0[61][39:32] = buffer_data_4[5119:5112];
        layer1[61][7:0] = buffer_data_3[5087:5080];
        layer1[61][15:8] = buffer_data_3[5095:5088];
        layer1[61][23:16] = buffer_data_3[5103:5096];
        layer1[61][31:24] = buffer_data_3[5111:5104];
        layer1[61][39:32] = buffer_data_3[5119:5112];
        layer2[61][7:0] = buffer_data_2[5087:5080];
        layer2[61][15:8] = buffer_data_2[5095:5088];
        layer2[61][23:16] = buffer_data_2[5103:5096];
        layer2[61][31:24] = buffer_data_2[5111:5104];
        layer2[61][39:32] = buffer_data_2[5119:5112];
        layer3[61][7:0] = buffer_data_1[5087:5080];
        layer3[61][15:8] = buffer_data_1[5095:5088];
        layer3[61][23:16] = buffer_data_1[5103:5096];
        layer3[61][31:24] = buffer_data_1[5111:5104];
        layer3[61][39:32] = buffer_data_1[5119:5112];
        layer4[61][7:0] = buffer_data_0[5087:5080];
        layer4[61][15:8] = buffer_data_0[5095:5088];
        layer4[61][23:16] = buffer_data_0[5103:5096];
        layer4[61][31:24] = buffer_data_0[5111:5104];
        layer4[61][39:32] = buffer_data_0[5119:5112];
        layer0[62][7:0] = buffer_data_4[5095:5088];
        layer0[62][15:8] = buffer_data_4[5103:5096];
        layer0[62][23:16] = buffer_data_4[5111:5104];
        layer0[62][31:24] = 0;
        layer0[62][39:32] = 0;
        layer1[62][7:0] = buffer_data_3[5095:5088];
        layer1[62][15:8] = buffer_data_3[5103:5096];
        layer1[62][23:16] = buffer_data_3[5111:5104];
        layer1[62][31:24] = 0;
        layer1[62][39:32] = 0;
        layer2[62][7:0] = buffer_data_2[5095:5088];
        layer2[62][15:8] = buffer_data_2[5103:5096];
        layer2[62][23:16] = buffer_data_2[5111:5104];
        layer2[62][31:24] = 0;
        layer2[62][39:32] = 0;
        layer3[62][7:0] = buffer_data_1[5095:5088];
        layer3[62][15:8] = buffer_data_1[5103:5096];
        layer3[62][23:16] = buffer_data_1[5111:5104];
        layer3[62][31:24] = 0;
        layer3[62][39:32] = 0;
        layer4[62][7:0] = buffer_data_0[5095:5088];
        layer4[62][15:8] = buffer_data_0[5103:5096];
        layer4[62][23:16] = buffer_data_0[5111:5104];
        layer4[62][31:24] = 0;
        layer4[62][39:32] = 0;
        layer0[63][7:0] = buffer_data_4[5103:5096];
        layer0[63][15:8] = buffer_data_4[5111:5104];
        layer0[63][23:16] = 0;
        layer0[63][31:24] = 0;
        layer0[63][39:32] = 0;
        layer1[63][7:0] = buffer_data_3[5103:5096];
        layer1[63][15:8] = buffer_data_3[5111:5104];
        layer1[63][23:16] = 0;
        layer1[63][31:24] = 0;
        layer1[63][39:32] = 0;
        layer2[63][7:0] = buffer_data_2[5103:5096];
        layer2[63][15:8] = buffer_data_2[5111:5104];
        layer2[63][23:16] = 0;
        layer2[63][31:24] = 0;
        layer2[63][39:32] = 0;
        layer3[63][7:0] = buffer_data_1[5103:5096];
        layer3[63][15:8] = buffer_data_1[5111:5104];
        layer3[63][23:16] = 0;
        layer3[63][31:24] = 0;
        layer3[63][39:32] = 0;
        layer4[63][7:0] = buffer_data_0[5103:5096];
        layer4[63][15:8] = buffer_data_0[5111:5104];
        layer4[63][23:16] = 0;
        layer4[63][31:24] = 0;
        layer4[63][39:32] = 0;
    end
  endcase
end

wire  [39:0]  kernel_img_mul_0[0:24];
assign kernel_img_mul_0[0] = layer0[0][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_0[1] = layer0[0][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_0[2] = layer0[0][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_0[3] = layer0[0][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_0[4] = layer0[0][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_0[5] = layer1[0][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_0[6] = layer1[0][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_0[7] = layer1[0][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_0[8] = layer1[0][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_0[9] = layer1[0][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_0[10] = layer2[0][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_0[11] = layer2[0][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_0[12] = layer2[0][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_0[13] = layer2[0][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_0[14] = layer2[0][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_0[15] = layer3[0][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_0[16] = layer3[0][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_0[17] = layer3[0][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_0[18] = layer3[0][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_0[19] = layer3[0][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_0[20] = layer4[0][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_0[21] = layer4[0][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_0[22] = layer4[0][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_0[23] = layer4[0][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_0[24] = layer4[0][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_0 = kernel_img_mul_0[0] + kernel_img_mul_0[1] + kernel_img_mul_0[2] + 
                kernel_img_mul_0[3] + kernel_img_mul_0[4] + kernel_img_mul_0[5] + 
                kernel_img_mul_0[6] + kernel_img_mul_0[7] + kernel_img_mul_0[8] + 
                kernel_img_mul_0[9] + kernel_img_mul_0[10] + kernel_img_mul_0[11] + 
                kernel_img_mul_0[12] + kernel_img_mul_0[13] + kernel_img_mul_0[14] + 
                kernel_img_mul_0[15] + kernel_img_mul_0[16] + kernel_img_mul_0[17] + 
                kernel_img_mul_0[18] + kernel_img_mul_0[19] + kernel_img_mul_0[20] + 
                kernel_img_mul_0[21] + kernel_img_mul_0[22] + kernel_img_mul_0[23] + 
                kernel_img_mul_0[24];
wire  [39:0]  kernel_img_mul_1[0:24];
assign kernel_img_mul_1[0] = layer0[1][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_1[1] = layer0[1][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_1[2] = layer0[1][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_1[3] = layer0[1][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_1[4] = layer0[1][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_1[5] = layer1[1][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_1[6] = layer1[1][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_1[7] = layer1[1][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_1[8] = layer1[1][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_1[9] = layer1[1][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_1[10] = layer2[1][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_1[11] = layer2[1][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_1[12] = layer2[1][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_1[13] = layer2[1][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_1[14] = layer2[1][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_1[15] = layer3[1][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_1[16] = layer3[1][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_1[17] = layer3[1][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_1[18] = layer3[1][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_1[19] = layer3[1][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_1[20] = layer4[1][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_1[21] = layer4[1][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_1[22] = layer4[1][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_1[23] = layer4[1][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_1[24] = layer4[1][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_1 = kernel_img_mul_1[0] + kernel_img_mul_1[1] + kernel_img_mul_1[2] + 
                kernel_img_mul_1[3] + kernel_img_mul_1[4] + kernel_img_mul_1[5] + 
                kernel_img_mul_1[6] + kernel_img_mul_1[7] + kernel_img_mul_1[8] + 
                kernel_img_mul_1[9] + kernel_img_mul_1[10] + kernel_img_mul_1[11] + 
                kernel_img_mul_1[12] + kernel_img_mul_1[13] + kernel_img_mul_1[14] + 
                kernel_img_mul_1[15] + kernel_img_mul_1[16] + kernel_img_mul_1[17] + 
                kernel_img_mul_1[18] + kernel_img_mul_1[19] + kernel_img_mul_1[20] + 
                kernel_img_mul_1[21] + kernel_img_mul_1[22] + kernel_img_mul_1[23] + 
                kernel_img_mul_1[24];
wire  [39:0]  kernel_img_mul_2[0:24];
assign kernel_img_mul_2[0] = layer0[2][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_2[1] = layer0[2][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_2[2] = layer0[2][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_2[3] = layer0[2][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_2[4] = layer0[2][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_2[5] = layer1[2][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_2[6] = layer1[2][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_2[7] = layer1[2][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_2[8] = layer1[2][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_2[9] = layer1[2][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_2[10] = layer2[2][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_2[11] = layer2[2][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_2[12] = layer2[2][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_2[13] = layer2[2][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_2[14] = layer2[2][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_2[15] = layer3[2][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_2[16] = layer3[2][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_2[17] = layer3[2][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_2[18] = layer3[2][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_2[19] = layer3[2][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_2[20] = layer4[2][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_2[21] = layer4[2][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_2[22] = layer4[2][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_2[23] = layer4[2][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_2[24] = layer4[2][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_2 = kernel_img_mul_2[0] + kernel_img_mul_2[1] + kernel_img_mul_2[2] + 
                kernel_img_mul_2[3] + kernel_img_mul_2[4] + kernel_img_mul_2[5] + 
                kernel_img_mul_2[6] + kernel_img_mul_2[7] + kernel_img_mul_2[8] + 
                kernel_img_mul_2[9] + kernel_img_mul_2[10] + kernel_img_mul_2[11] + 
                kernel_img_mul_2[12] + kernel_img_mul_2[13] + kernel_img_mul_2[14] + 
                kernel_img_mul_2[15] + kernel_img_mul_2[16] + kernel_img_mul_2[17] + 
                kernel_img_mul_2[18] + kernel_img_mul_2[19] + kernel_img_mul_2[20] + 
                kernel_img_mul_2[21] + kernel_img_mul_2[22] + kernel_img_mul_2[23] + 
                kernel_img_mul_2[24];
wire  [39:0]  kernel_img_mul_3[0:24];
assign kernel_img_mul_3[0] = layer0[3][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_3[1] = layer0[3][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_3[2] = layer0[3][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_3[3] = layer0[3][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_3[4] = layer0[3][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_3[5] = layer1[3][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_3[6] = layer1[3][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_3[7] = layer1[3][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_3[8] = layer1[3][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_3[9] = layer1[3][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_3[10] = layer2[3][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_3[11] = layer2[3][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_3[12] = layer2[3][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_3[13] = layer2[3][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_3[14] = layer2[3][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_3[15] = layer3[3][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_3[16] = layer3[3][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_3[17] = layer3[3][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_3[18] = layer3[3][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_3[19] = layer3[3][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_3[20] = layer4[3][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_3[21] = layer4[3][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_3[22] = layer4[3][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_3[23] = layer4[3][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_3[24] = layer4[3][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_3 = kernel_img_mul_3[0] + kernel_img_mul_3[1] + kernel_img_mul_3[2] + 
                kernel_img_mul_3[3] + kernel_img_mul_3[4] + kernel_img_mul_3[5] + 
                kernel_img_mul_3[6] + kernel_img_mul_3[7] + kernel_img_mul_3[8] + 
                kernel_img_mul_3[9] + kernel_img_mul_3[10] + kernel_img_mul_3[11] + 
                kernel_img_mul_3[12] + kernel_img_mul_3[13] + kernel_img_mul_3[14] + 
                kernel_img_mul_3[15] + kernel_img_mul_3[16] + kernel_img_mul_3[17] + 
                kernel_img_mul_3[18] + kernel_img_mul_3[19] + kernel_img_mul_3[20] + 
                kernel_img_mul_3[21] + kernel_img_mul_3[22] + kernel_img_mul_3[23] + 
                kernel_img_mul_3[24];
wire  [39:0]  kernel_img_mul_4[0:24];
assign kernel_img_mul_4[0] = layer0[4][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_4[1] = layer0[4][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_4[2] = layer0[4][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_4[3] = layer0[4][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_4[4] = layer0[4][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_4[5] = layer1[4][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_4[6] = layer1[4][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_4[7] = layer1[4][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_4[8] = layer1[4][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_4[9] = layer1[4][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_4[10] = layer2[4][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_4[11] = layer2[4][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_4[12] = layer2[4][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_4[13] = layer2[4][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_4[14] = layer2[4][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_4[15] = layer3[4][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_4[16] = layer3[4][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_4[17] = layer3[4][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_4[18] = layer3[4][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_4[19] = layer3[4][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_4[20] = layer4[4][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_4[21] = layer4[4][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_4[22] = layer4[4][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_4[23] = layer4[4][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_4[24] = layer4[4][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_4 = kernel_img_mul_4[0] + kernel_img_mul_4[1] + kernel_img_mul_4[2] + 
                kernel_img_mul_4[3] + kernel_img_mul_4[4] + kernel_img_mul_4[5] + 
                kernel_img_mul_4[6] + kernel_img_mul_4[7] + kernel_img_mul_4[8] + 
                kernel_img_mul_4[9] + kernel_img_mul_4[10] + kernel_img_mul_4[11] + 
                kernel_img_mul_4[12] + kernel_img_mul_4[13] + kernel_img_mul_4[14] + 
                kernel_img_mul_4[15] + kernel_img_mul_4[16] + kernel_img_mul_4[17] + 
                kernel_img_mul_4[18] + kernel_img_mul_4[19] + kernel_img_mul_4[20] + 
                kernel_img_mul_4[21] + kernel_img_mul_4[22] + kernel_img_mul_4[23] + 
                kernel_img_mul_4[24];
wire  [39:0]  kernel_img_mul_5[0:24];
assign kernel_img_mul_5[0] = layer0[5][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_5[1] = layer0[5][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_5[2] = layer0[5][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_5[3] = layer0[5][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_5[4] = layer0[5][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_5[5] = layer1[5][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_5[6] = layer1[5][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_5[7] = layer1[5][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_5[8] = layer1[5][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_5[9] = layer1[5][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_5[10] = layer2[5][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_5[11] = layer2[5][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_5[12] = layer2[5][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_5[13] = layer2[5][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_5[14] = layer2[5][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_5[15] = layer3[5][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_5[16] = layer3[5][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_5[17] = layer3[5][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_5[18] = layer3[5][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_5[19] = layer3[5][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_5[20] = layer4[5][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_5[21] = layer4[5][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_5[22] = layer4[5][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_5[23] = layer4[5][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_5[24] = layer4[5][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_5 = kernel_img_mul_5[0] + kernel_img_mul_5[1] + kernel_img_mul_5[2] + 
                kernel_img_mul_5[3] + kernel_img_mul_5[4] + kernel_img_mul_5[5] + 
                kernel_img_mul_5[6] + kernel_img_mul_5[7] + kernel_img_mul_5[8] + 
                kernel_img_mul_5[9] + kernel_img_mul_5[10] + kernel_img_mul_5[11] + 
                kernel_img_mul_5[12] + kernel_img_mul_5[13] + kernel_img_mul_5[14] + 
                kernel_img_mul_5[15] + kernel_img_mul_5[16] + kernel_img_mul_5[17] + 
                kernel_img_mul_5[18] + kernel_img_mul_5[19] + kernel_img_mul_5[20] + 
                kernel_img_mul_5[21] + kernel_img_mul_5[22] + kernel_img_mul_5[23] + 
                kernel_img_mul_5[24];
wire  [39:0]  kernel_img_mul_6[0:24];
assign kernel_img_mul_6[0] = layer0[6][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_6[1] = layer0[6][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_6[2] = layer0[6][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_6[3] = layer0[6][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_6[4] = layer0[6][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_6[5] = layer1[6][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_6[6] = layer1[6][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_6[7] = layer1[6][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_6[8] = layer1[6][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_6[9] = layer1[6][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_6[10] = layer2[6][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_6[11] = layer2[6][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_6[12] = layer2[6][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_6[13] = layer2[6][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_6[14] = layer2[6][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_6[15] = layer3[6][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_6[16] = layer3[6][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_6[17] = layer3[6][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_6[18] = layer3[6][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_6[19] = layer3[6][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_6[20] = layer4[6][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_6[21] = layer4[6][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_6[22] = layer4[6][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_6[23] = layer4[6][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_6[24] = layer4[6][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_6 = kernel_img_mul_6[0] + kernel_img_mul_6[1] + kernel_img_mul_6[2] + 
                kernel_img_mul_6[3] + kernel_img_mul_6[4] + kernel_img_mul_6[5] + 
                kernel_img_mul_6[6] + kernel_img_mul_6[7] + kernel_img_mul_6[8] + 
                kernel_img_mul_6[9] + kernel_img_mul_6[10] + kernel_img_mul_6[11] + 
                kernel_img_mul_6[12] + kernel_img_mul_6[13] + kernel_img_mul_6[14] + 
                kernel_img_mul_6[15] + kernel_img_mul_6[16] + kernel_img_mul_6[17] + 
                kernel_img_mul_6[18] + kernel_img_mul_6[19] + kernel_img_mul_6[20] + 
                kernel_img_mul_6[21] + kernel_img_mul_6[22] + kernel_img_mul_6[23] + 
                kernel_img_mul_6[24];
wire  [39:0]  kernel_img_mul_7[0:24];
assign kernel_img_mul_7[0] = layer0[7][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_7[1] = layer0[7][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_7[2] = layer0[7][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_7[3] = layer0[7][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_7[4] = layer0[7][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_7[5] = layer1[7][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_7[6] = layer1[7][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_7[7] = layer1[7][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_7[8] = layer1[7][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_7[9] = layer1[7][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_7[10] = layer2[7][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_7[11] = layer2[7][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_7[12] = layer2[7][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_7[13] = layer2[7][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_7[14] = layer2[7][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_7[15] = layer3[7][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_7[16] = layer3[7][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_7[17] = layer3[7][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_7[18] = layer3[7][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_7[19] = layer3[7][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_7[20] = layer4[7][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_7[21] = layer4[7][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_7[22] = layer4[7][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_7[23] = layer4[7][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_7[24] = layer4[7][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_7 = kernel_img_mul_7[0] + kernel_img_mul_7[1] + kernel_img_mul_7[2] + 
                kernel_img_mul_7[3] + kernel_img_mul_7[4] + kernel_img_mul_7[5] + 
                kernel_img_mul_7[6] + kernel_img_mul_7[7] + kernel_img_mul_7[8] + 
                kernel_img_mul_7[9] + kernel_img_mul_7[10] + kernel_img_mul_7[11] + 
                kernel_img_mul_7[12] + kernel_img_mul_7[13] + kernel_img_mul_7[14] + 
                kernel_img_mul_7[15] + kernel_img_mul_7[16] + kernel_img_mul_7[17] + 
                kernel_img_mul_7[18] + kernel_img_mul_7[19] + kernel_img_mul_7[20] + 
                kernel_img_mul_7[21] + kernel_img_mul_7[22] + kernel_img_mul_7[23] + 
                kernel_img_mul_7[24];
wire  [39:0]  kernel_img_mul_8[0:24];
assign kernel_img_mul_8[0] = layer0[8][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_8[1] = layer0[8][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_8[2] = layer0[8][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_8[3] = layer0[8][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_8[4] = layer0[8][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_8[5] = layer1[8][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_8[6] = layer1[8][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_8[7] = layer1[8][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_8[8] = layer1[8][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_8[9] = layer1[8][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_8[10] = layer2[8][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_8[11] = layer2[8][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_8[12] = layer2[8][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_8[13] = layer2[8][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_8[14] = layer2[8][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_8[15] = layer3[8][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_8[16] = layer3[8][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_8[17] = layer3[8][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_8[18] = layer3[8][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_8[19] = layer3[8][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_8[20] = layer4[8][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_8[21] = layer4[8][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_8[22] = layer4[8][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_8[23] = layer4[8][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_8[24] = layer4[8][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_8 = kernel_img_mul_8[0] + kernel_img_mul_8[1] + kernel_img_mul_8[2] + 
                kernel_img_mul_8[3] + kernel_img_mul_8[4] + kernel_img_mul_8[5] + 
                kernel_img_mul_8[6] + kernel_img_mul_8[7] + kernel_img_mul_8[8] + 
                kernel_img_mul_8[9] + kernel_img_mul_8[10] + kernel_img_mul_8[11] + 
                kernel_img_mul_8[12] + kernel_img_mul_8[13] + kernel_img_mul_8[14] + 
                kernel_img_mul_8[15] + kernel_img_mul_8[16] + kernel_img_mul_8[17] + 
                kernel_img_mul_8[18] + kernel_img_mul_8[19] + kernel_img_mul_8[20] + 
                kernel_img_mul_8[21] + kernel_img_mul_8[22] + kernel_img_mul_8[23] + 
                kernel_img_mul_8[24];
wire  [39:0]  kernel_img_mul_9[0:24];
assign kernel_img_mul_9[0] = layer0[9][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_9[1] = layer0[9][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_9[2] = layer0[9][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_9[3] = layer0[9][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_9[4] = layer0[9][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_9[5] = layer1[9][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_9[6] = layer1[9][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_9[7] = layer1[9][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_9[8] = layer1[9][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_9[9] = layer1[9][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_9[10] = layer2[9][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_9[11] = layer2[9][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_9[12] = layer2[9][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_9[13] = layer2[9][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_9[14] = layer2[9][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_9[15] = layer3[9][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_9[16] = layer3[9][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_9[17] = layer3[9][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_9[18] = layer3[9][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_9[19] = layer3[9][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_9[20] = layer4[9][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_9[21] = layer4[9][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_9[22] = layer4[9][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_9[23] = layer4[9][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_9[24] = layer4[9][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_9 = kernel_img_mul_9[0] + kernel_img_mul_9[1] + kernel_img_mul_9[2] + 
                kernel_img_mul_9[3] + kernel_img_mul_9[4] + kernel_img_mul_9[5] + 
                kernel_img_mul_9[6] + kernel_img_mul_9[7] + kernel_img_mul_9[8] + 
                kernel_img_mul_9[9] + kernel_img_mul_9[10] + kernel_img_mul_9[11] + 
                kernel_img_mul_9[12] + kernel_img_mul_9[13] + kernel_img_mul_9[14] + 
                kernel_img_mul_9[15] + kernel_img_mul_9[16] + kernel_img_mul_9[17] + 
                kernel_img_mul_9[18] + kernel_img_mul_9[19] + kernel_img_mul_9[20] + 
                kernel_img_mul_9[21] + kernel_img_mul_9[22] + kernel_img_mul_9[23] + 
                kernel_img_mul_9[24];
wire  [39:0]  kernel_img_mul_10[0:24];
assign kernel_img_mul_10[0] = layer0[10][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_10[1] = layer0[10][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_10[2] = layer0[10][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_10[3] = layer0[10][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_10[4] = layer0[10][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_10[5] = layer1[10][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_10[6] = layer1[10][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_10[7] = layer1[10][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_10[8] = layer1[10][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_10[9] = layer1[10][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_10[10] = layer2[10][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_10[11] = layer2[10][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_10[12] = layer2[10][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_10[13] = layer2[10][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_10[14] = layer2[10][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_10[15] = layer3[10][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_10[16] = layer3[10][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_10[17] = layer3[10][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_10[18] = layer3[10][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_10[19] = layer3[10][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_10[20] = layer4[10][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_10[21] = layer4[10][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_10[22] = layer4[10][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_10[23] = layer4[10][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_10[24] = layer4[10][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_10 = kernel_img_mul_10[0] + kernel_img_mul_10[1] + kernel_img_mul_10[2] + 
                kernel_img_mul_10[3] + kernel_img_mul_10[4] + kernel_img_mul_10[5] + 
                kernel_img_mul_10[6] + kernel_img_mul_10[7] + kernel_img_mul_10[8] + 
                kernel_img_mul_10[9] + kernel_img_mul_10[10] + kernel_img_mul_10[11] + 
                kernel_img_mul_10[12] + kernel_img_mul_10[13] + kernel_img_mul_10[14] + 
                kernel_img_mul_10[15] + kernel_img_mul_10[16] + kernel_img_mul_10[17] + 
                kernel_img_mul_10[18] + kernel_img_mul_10[19] + kernel_img_mul_10[20] + 
                kernel_img_mul_10[21] + kernel_img_mul_10[22] + kernel_img_mul_10[23] + 
                kernel_img_mul_10[24];
wire  [39:0]  kernel_img_mul_11[0:24];
assign kernel_img_mul_11[0] = layer0[11][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_11[1] = layer0[11][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_11[2] = layer0[11][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_11[3] = layer0[11][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_11[4] = layer0[11][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_11[5] = layer1[11][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_11[6] = layer1[11][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_11[7] = layer1[11][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_11[8] = layer1[11][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_11[9] = layer1[11][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_11[10] = layer2[11][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_11[11] = layer2[11][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_11[12] = layer2[11][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_11[13] = layer2[11][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_11[14] = layer2[11][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_11[15] = layer3[11][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_11[16] = layer3[11][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_11[17] = layer3[11][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_11[18] = layer3[11][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_11[19] = layer3[11][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_11[20] = layer4[11][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_11[21] = layer4[11][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_11[22] = layer4[11][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_11[23] = layer4[11][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_11[24] = layer4[11][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_11 = kernel_img_mul_11[0] + kernel_img_mul_11[1] + kernel_img_mul_11[2] + 
                kernel_img_mul_11[3] + kernel_img_mul_11[4] + kernel_img_mul_11[5] + 
                kernel_img_mul_11[6] + kernel_img_mul_11[7] + kernel_img_mul_11[8] + 
                kernel_img_mul_11[9] + kernel_img_mul_11[10] + kernel_img_mul_11[11] + 
                kernel_img_mul_11[12] + kernel_img_mul_11[13] + kernel_img_mul_11[14] + 
                kernel_img_mul_11[15] + kernel_img_mul_11[16] + kernel_img_mul_11[17] + 
                kernel_img_mul_11[18] + kernel_img_mul_11[19] + kernel_img_mul_11[20] + 
                kernel_img_mul_11[21] + kernel_img_mul_11[22] + kernel_img_mul_11[23] + 
                kernel_img_mul_11[24];
wire  [39:0]  kernel_img_mul_12[0:24];
assign kernel_img_mul_12[0] = layer0[12][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_12[1] = layer0[12][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_12[2] = layer0[12][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_12[3] = layer0[12][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_12[4] = layer0[12][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_12[5] = layer1[12][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_12[6] = layer1[12][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_12[7] = layer1[12][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_12[8] = layer1[12][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_12[9] = layer1[12][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_12[10] = layer2[12][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_12[11] = layer2[12][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_12[12] = layer2[12][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_12[13] = layer2[12][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_12[14] = layer2[12][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_12[15] = layer3[12][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_12[16] = layer3[12][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_12[17] = layer3[12][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_12[18] = layer3[12][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_12[19] = layer3[12][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_12[20] = layer4[12][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_12[21] = layer4[12][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_12[22] = layer4[12][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_12[23] = layer4[12][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_12[24] = layer4[12][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_12 = kernel_img_mul_12[0] + kernel_img_mul_12[1] + kernel_img_mul_12[2] + 
                kernel_img_mul_12[3] + kernel_img_mul_12[4] + kernel_img_mul_12[5] + 
                kernel_img_mul_12[6] + kernel_img_mul_12[7] + kernel_img_mul_12[8] + 
                kernel_img_mul_12[9] + kernel_img_mul_12[10] + kernel_img_mul_12[11] + 
                kernel_img_mul_12[12] + kernel_img_mul_12[13] + kernel_img_mul_12[14] + 
                kernel_img_mul_12[15] + kernel_img_mul_12[16] + kernel_img_mul_12[17] + 
                kernel_img_mul_12[18] + kernel_img_mul_12[19] + kernel_img_mul_12[20] + 
                kernel_img_mul_12[21] + kernel_img_mul_12[22] + kernel_img_mul_12[23] + 
                kernel_img_mul_12[24];
wire  [39:0]  kernel_img_mul_13[0:24];
assign kernel_img_mul_13[0] = layer0[13][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_13[1] = layer0[13][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_13[2] = layer0[13][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_13[3] = layer0[13][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_13[4] = layer0[13][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_13[5] = layer1[13][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_13[6] = layer1[13][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_13[7] = layer1[13][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_13[8] = layer1[13][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_13[9] = layer1[13][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_13[10] = layer2[13][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_13[11] = layer2[13][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_13[12] = layer2[13][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_13[13] = layer2[13][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_13[14] = layer2[13][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_13[15] = layer3[13][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_13[16] = layer3[13][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_13[17] = layer3[13][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_13[18] = layer3[13][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_13[19] = layer3[13][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_13[20] = layer4[13][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_13[21] = layer4[13][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_13[22] = layer4[13][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_13[23] = layer4[13][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_13[24] = layer4[13][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_13 = kernel_img_mul_13[0] + kernel_img_mul_13[1] + kernel_img_mul_13[2] + 
                kernel_img_mul_13[3] + kernel_img_mul_13[4] + kernel_img_mul_13[5] + 
                kernel_img_mul_13[6] + kernel_img_mul_13[7] + kernel_img_mul_13[8] + 
                kernel_img_mul_13[9] + kernel_img_mul_13[10] + kernel_img_mul_13[11] + 
                kernel_img_mul_13[12] + kernel_img_mul_13[13] + kernel_img_mul_13[14] + 
                kernel_img_mul_13[15] + kernel_img_mul_13[16] + kernel_img_mul_13[17] + 
                kernel_img_mul_13[18] + kernel_img_mul_13[19] + kernel_img_mul_13[20] + 
                kernel_img_mul_13[21] + kernel_img_mul_13[22] + kernel_img_mul_13[23] + 
                kernel_img_mul_13[24];
wire  [39:0]  kernel_img_mul_14[0:24];
assign kernel_img_mul_14[0] = layer0[14][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_14[1] = layer0[14][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_14[2] = layer0[14][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_14[3] = layer0[14][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_14[4] = layer0[14][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_14[5] = layer1[14][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_14[6] = layer1[14][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_14[7] = layer1[14][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_14[8] = layer1[14][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_14[9] = layer1[14][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_14[10] = layer2[14][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_14[11] = layer2[14][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_14[12] = layer2[14][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_14[13] = layer2[14][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_14[14] = layer2[14][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_14[15] = layer3[14][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_14[16] = layer3[14][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_14[17] = layer3[14][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_14[18] = layer3[14][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_14[19] = layer3[14][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_14[20] = layer4[14][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_14[21] = layer4[14][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_14[22] = layer4[14][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_14[23] = layer4[14][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_14[24] = layer4[14][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_14 = kernel_img_mul_14[0] + kernel_img_mul_14[1] + kernel_img_mul_14[2] + 
                kernel_img_mul_14[3] + kernel_img_mul_14[4] + kernel_img_mul_14[5] + 
                kernel_img_mul_14[6] + kernel_img_mul_14[7] + kernel_img_mul_14[8] + 
                kernel_img_mul_14[9] + kernel_img_mul_14[10] + kernel_img_mul_14[11] + 
                kernel_img_mul_14[12] + kernel_img_mul_14[13] + kernel_img_mul_14[14] + 
                kernel_img_mul_14[15] + kernel_img_mul_14[16] + kernel_img_mul_14[17] + 
                kernel_img_mul_14[18] + kernel_img_mul_14[19] + kernel_img_mul_14[20] + 
                kernel_img_mul_14[21] + kernel_img_mul_14[22] + kernel_img_mul_14[23] + 
                kernel_img_mul_14[24];
wire  [39:0]  kernel_img_mul_15[0:24];
assign kernel_img_mul_15[0] = layer0[15][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_15[1] = layer0[15][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_15[2] = layer0[15][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_15[3] = layer0[15][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_15[4] = layer0[15][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_15[5] = layer1[15][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_15[6] = layer1[15][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_15[7] = layer1[15][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_15[8] = layer1[15][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_15[9] = layer1[15][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_15[10] = layer2[15][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_15[11] = layer2[15][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_15[12] = layer2[15][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_15[13] = layer2[15][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_15[14] = layer2[15][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_15[15] = layer3[15][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_15[16] = layer3[15][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_15[17] = layer3[15][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_15[18] = layer3[15][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_15[19] = layer3[15][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_15[20] = layer4[15][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_15[21] = layer4[15][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_15[22] = layer4[15][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_15[23] = layer4[15][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_15[24] = layer4[15][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_15 = kernel_img_mul_15[0] + kernel_img_mul_15[1] + kernel_img_mul_15[2] + 
                kernel_img_mul_15[3] + kernel_img_mul_15[4] + kernel_img_mul_15[5] + 
                kernel_img_mul_15[6] + kernel_img_mul_15[7] + kernel_img_mul_15[8] + 
                kernel_img_mul_15[9] + kernel_img_mul_15[10] + kernel_img_mul_15[11] + 
                kernel_img_mul_15[12] + kernel_img_mul_15[13] + kernel_img_mul_15[14] + 
                kernel_img_mul_15[15] + kernel_img_mul_15[16] + kernel_img_mul_15[17] + 
                kernel_img_mul_15[18] + kernel_img_mul_15[19] + kernel_img_mul_15[20] + 
                kernel_img_mul_15[21] + kernel_img_mul_15[22] + kernel_img_mul_15[23] + 
                kernel_img_mul_15[24];
wire  [39:0]  kernel_img_mul_16[0:24];
assign kernel_img_mul_16[0] = layer0[16][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_16[1] = layer0[16][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_16[2] = layer0[16][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_16[3] = layer0[16][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_16[4] = layer0[16][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_16[5] = layer1[16][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_16[6] = layer1[16][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_16[7] = layer1[16][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_16[8] = layer1[16][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_16[9] = layer1[16][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_16[10] = layer2[16][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_16[11] = layer2[16][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_16[12] = layer2[16][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_16[13] = layer2[16][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_16[14] = layer2[16][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_16[15] = layer3[16][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_16[16] = layer3[16][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_16[17] = layer3[16][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_16[18] = layer3[16][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_16[19] = layer3[16][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_16[20] = layer4[16][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_16[21] = layer4[16][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_16[22] = layer4[16][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_16[23] = layer4[16][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_16[24] = layer4[16][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_16 = kernel_img_mul_16[0] + kernel_img_mul_16[1] + kernel_img_mul_16[2] + 
                kernel_img_mul_16[3] + kernel_img_mul_16[4] + kernel_img_mul_16[5] + 
                kernel_img_mul_16[6] + kernel_img_mul_16[7] + kernel_img_mul_16[8] + 
                kernel_img_mul_16[9] + kernel_img_mul_16[10] + kernel_img_mul_16[11] + 
                kernel_img_mul_16[12] + kernel_img_mul_16[13] + kernel_img_mul_16[14] + 
                kernel_img_mul_16[15] + kernel_img_mul_16[16] + kernel_img_mul_16[17] + 
                kernel_img_mul_16[18] + kernel_img_mul_16[19] + kernel_img_mul_16[20] + 
                kernel_img_mul_16[21] + kernel_img_mul_16[22] + kernel_img_mul_16[23] + 
                kernel_img_mul_16[24];
wire  [39:0]  kernel_img_mul_17[0:24];
assign kernel_img_mul_17[0] = layer0[17][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_17[1] = layer0[17][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_17[2] = layer0[17][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_17[3] = layer0[17][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_17[4] = layer0[17][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_17[5] = layer1[17][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_17[6] = layer1[17][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_17[7] = layer1[17][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_17[8] = layer1[17][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_17[9] = layer1[17][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_17[10] = layer2[17][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_17[11] = layer2[17][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_17[12] = layer2[17][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_17[13] = layer2[17][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_17[14] = layer2[17][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_17[15] = layer3[17][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_17[16] = layer3[17][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_17[17] = layer3[17][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_17[18] = layer3[17][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_17[19] = layer3[17][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_17[20] = layer4[17][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_17[21] = layer4[17][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_17[22] = layer4[17][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_17[23] = layer4[17][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_17[24] = layer4[17][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_17 = kernel_img_mul_17[0] + kernel_img_mul_17[1] + kernel_img_mul_17[2] + 
                kernel_img_mul_17[3] + kernel_img_mul_17[4] + kernel_img_mul_17[5] + 
                kernel_img_mul_17[6] + kernel_img_mul_17[7] + kernel_img_mul_17[8] + 
                kernel_img_mul_17[9] + kernel_img_mul_17[10] + kernel_img_mul_17[11] + 
                kernel_img_mul_17[12] + kernel_img_mul_17[13] + kernel_img_mul_17[14] + 
                kernel_img_mul_17[15] + kernel_img_mul_17[16] + kernel_img_mul_17[17] + 
                kernel_img_mul_17[18] + kernel_img_mul_17[19] + kernel_img_mul_17[20] + 
                kernel_img_mul_17[21] + kernel_img_mul_17[22] + kernel_img_mul_17[23] + 
                kernel_img_mul_17[24];
wire  [39:0]  kernel_img_mul_18[0:24];
assign kernel_img_mul_18[0] = layer0[18][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_18[1] = layer0[18][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_18[2] = layer0[18][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_18[3] = layer0[18][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_18[4] = layer0[18][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_18[5] = layer1[18][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_18[6] = layer1[18][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_18[7] = layer1[18][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_18[8] = layer1[18][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_18[9] = layer1[18][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_18[10] = layer2[18][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_18[11] = layer2[18][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_18[12] = layer2[18][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_18[13] = layer2[18][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_18[14] = layer2[18][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_18[15] = layer3[18][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_18[16] = layer3[18][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_18[17] = layer3[18][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_18[18] = layer3[18][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_18[19] = layer3[18][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_18[20] = layer4[18][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_18[21] = layer4[18][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_18[22] = layer4[18][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_18[23] = layer4[18][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_18[24] = layer4[18][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_18 = kernel_img_mul_18[0] + kernel_img_mul_18[1] + kernel_img_mul_18[2] + 
                kernel_img_mul_18[3] + kernel_img_mul_18[4] + kernel_img_mul_18[5] + 
                kernel_img_mul_18[6] + kernel_img_mul_18[7] + kernel_img_mul_18[8] + 
                kernel_img_mul_18[9] + kernel_img_mul_18[10] + kernel_img_mul_18[11] + 
                kernel_img_mul_18[12] + kernel_img_mul_18[13] + kernel_img_mul_18[14] + 
                kernel_img_mul_18[15] + kernel_img_mul_18[16] + kernel_img_mul_18[17] + 
                kernel_img_mul_18[18] + kernel_img_mul_18[19] + kernel_img_mul_18[20] + 
                kernel_img_mul_18[21] + kernel_img_mul_18[22] + kernel_img_mul_18[23] + 
                kernel_img_mul_18[24];
wire  [39:0]  kernel_img_mul_19[0:24];
assign kernel_img_mul_19[0] = layer0[19][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_19[1] = layer0[19][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_19[2] = layer0[19][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_19[3] = layer0[19][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_19[4] = layer0[19][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_19[5] = layer1[19][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_19[6] = layer1[19][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_19[7] = layer1[19][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_19[8] = layer1[19][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_19[9] = layer1[19][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_19[10] = layer2[19][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_19[11] = layer2[19][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_19[12] = layer2[19][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_19[13] = layer2[19][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_19[14] = layer2[19][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_19[15] = layer3[19][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_19[16] = layer3[19][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_19[17] = layer3[19][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_19[18] = layer3[19][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_19[19] = layer3[19][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_19[20] = layer4[19][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_19[21] = layer4[19][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_19[22] = layer4[19][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_19[23] = layer4[19][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_19[24] = layer4[19][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_19 = kernel_img_mul_19[0] + kernel_img_mul_19[1] + kernel_img_mul_19[2] + 
                kernel_img_mul_19[3] + kernel_img_mul_19[4] + kernel_img_mul_19[5] + 
                kernel_img_mul_19[6] + kernel_img_mul_19[7] + kernel_img_mul_19[8] + 
                kernel_img_mul_19[9] + kernel_img_mul_19[10] + kernel_img_mul_19[11] + 
                kernel_img_mul_19[12] + kernel_img_mul_19[13] + kernel_img_mul_19[14] + 
                kernel_img_mul_19[15] + kernel_img_mul_19[16] + kernel_img_mul_19[17] + 
                kernel_img_mul_19[18] + kernel_img_mul_19[19] + kernel_img_mul_19[20] + 
                kernel_img_mul_19[21] + kernel_img_mul_19[22] + kernel_img_mul_19[23] + 
                kernel_img_mul_19[24];
wire  [39:0]  kernel_img_mul_20[0:24];
assign kernel_img_mul_20[0] = layer0[20][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_20[1] = layer0[20][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_20[2] = layer0[20][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_20[3] = layer0[20][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_20[4] = layer0[20][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_20[5] = layer1[20][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_20[6] = layer1[20][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_20[7] = layer1[20][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_20[8] = layer1[20][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_20[9] = layer1[20][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_20[10] = layer2[20][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_20[11] = layer2[20][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_20[12] = layer2[20][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_20[13] = layer2[20][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_20[14] = layer2[20][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_20[15] = layer3[20][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_20[16] = layer3[20][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_20[17] = layer3[20][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_20[18] = layer3[20][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_20[19] = layer3[20][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_20[20] = layer4[20][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_20[21] = layer4[20][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_20[22] = layer4[20][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_20[23] = layer4[20][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_20[24] = layer4[20][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_20 = kernel_img_mul_20[0] + kernel_img_mul_20[1] + kernel_img_mul_20[2] + 
                kernel_img_mul_20[3] + kernel_img_mul_20[4] + kernel_img_mul_20[5] + 
                kernel_img_mul_20[6] + kernel_img_mul_20[7] + kernel_img_mul_20[8] + 
                kernel_img_mul_20[9] + kernel_img_mul_20[10] + kernel_img_mul_20[11] + 
                kernel_img_mul_20[12] + kernel_img_mul_20[13] + kernel_img_mul_20[14] + 
                kernel_img_mul_20[15] + kernel_img_mul_20[16] + kernel_img_mul_20[17] + 
                kernel_img_mul_20[18] + kernel_img_mul_20[19] + kernel_img_mul_20[20] + 
                kernel_img_mul_20[21] + kernel_img_mul_20[22] + kernel_img_mul_20[23] + 
                kernel_img_mul_20[24];
wire  [39:0]  kernel_img_mul_21[0:24];
assign kernel_img_mul_21[0] = layer0[21][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_21[1] = layer0[21][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_21[2] = layer0[21][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_21[3] = layer0[21][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_21[4] = layer0[21][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_21[5] = layer1[21][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_21[6] = layer1[21][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_21[7] = layer1[21][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_21[8] = layer1[21][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_21[9] = layer1[21][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_21[10] = layer2[21][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_21[11] = layer2[21][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_21[12] = layer2[21][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_21[13] = layer2[21][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_21[14] = layer2[21][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_21[15] = layer3[21][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_21[16] = layer3[21][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_21[17] = layer3[21][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_21[18] = layer3[21][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_21[19] = layer3[21][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_21[20] = layer4[21][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_21[21] = layer4[21][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_21[22] = layer4[21][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_21[23] = layer4[21][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_21[24] = layer4[21][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_21 = kernel_img_mul_21[0] + kernel_img_mul_21[1] + kernel_img_mul_21[2] + 
                kernel_img_mul_21[3] + kernel_img_mul_21[4] + kernel_img_mul_21[5] + 
                kernel_img_mul_21[6] + kernel_img_mul_21[7] + kernel_img_mul_21[8] + 
                kernel_img_mul_21[9] + kernel_img_mul_21[10] + kernel_img_mul_21[11] + 
                kernel_img_mul_21[12] + kernel_img_mul_21[13] + kernel_img_mul_21[14] + 
                kernel_img_mul_21[15] + kernel_img_mul_21[16] + kernel_img_mul_21[17] + 
                kernel_img_mul_21[18] + kernel_img_mul_21[19] + kernel_img_mul_21[20] + 
                kernel_img_mul_21[21] + kernel_img_mul_21[22] + kernel_img_mul_21[23] + 
                kernel_img_mul_21[24];
wire  [39:0]  kernel_img_mul_22[0:24];
assign kernel_img_mul_22[0] = layer0[22][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_22[1] = layer0[22][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_22[2] = layer0[22][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_22[3] = layer0[22][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_22[4] = layer0[22][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_22[5] = layer1[22][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_22[6] = layer1[22][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_22[7] = layer1[22][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_22[8] = layer1[22][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_22[9] = layer1[22][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_22[10] = layer2[22][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_22[11] = layer2[22][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_22[12] = layer2[22][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_22[13] = layer2[22][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_22[14] = layer2[22][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_22[15] = layer3[22][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_22[16] = layer3[22][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_22[17] = layer3[22][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_22[18] = layer3[22][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_22[19] = layer3[22][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_22[20] = layer4[22][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_22[21] = layer4[22][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_22[22] = layer4[22][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_22[23] = layer4[22][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_22[24] = layer4[22][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_22 = kernel_img_mul_22[0] + kernel_img_mul_22[1] + kernel_img_mul_22[2] + 
                kernel_img_mul_22[3] + kernel_img_mul_22[4] + kernel_img_mul_22[5] + 
                kernel_img_mul_22[6] + kernel_img_mul_22[7] + kernel_img_mul_22[8] + 
                kernel_img_mul_22[9] + kernel_img_mul_22[10] + kernel_img_mul_22[11] + 
                kernel_img_mul_22[12] + kernel_img_mul_22[13] + kernel_img_mul_22[14] + 
                kernel_img_mul_22[15] + kernel_img_mul_22[16] + kernel_img_mul_22[17] + 
                kernel_img_mul_22[18] + kernel_img_mul_22[19] + kernel_img_mul_22[20] + 
                kernel_img_mul_22[21] + kernel_img_mul_22[22] + kernel_img_mul_22[23] + 
                kernel_img_mul_22[24];
wire  [39:0]  kernel_img_mul_23[0:24];
assign kernel_img_mul_23[0] = layer0[23][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_23[1] = layer0[23][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_23[2] = layer0[23][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_23[3] = layer0[23][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_23[4] = layer0[23][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_23[5] = layer1[23][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_23[6] = layer1[23][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_23[7] = layer1[23][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_23[8] = layer1[23][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_23[9] = layer1[23][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_23[10] = layer2[23][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_23[11] = layer2[23][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_23[12] = layer2[23][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_23[13] = layer2[23][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_23[14] = layer2[23][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_23[15] = layer3[23][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_23[16] = layer3[23][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_23[17] = layer3[23][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_23[18] = layer3[23][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_23[19] = layer3[23][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_23[20] = layer4[23][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_23[21] = layer4[23][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_23[22] = layer4[23][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_23[23] = layer4[23][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_23[24] = layer4[23][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_23 = kernel_img_mul_23[0] + kernel_img_mul_23[1] + kernel_img_mul_23[2] + 
                kernel_img_mul_23[3] + kernel_img_mul_23[4] + kernel_img_mul_23[5] + 
                kernel_img_mul_23[6] + kernel_img_mul_23[7] + kernel_img_mul_23[8] + 
                kernel_img_mul_23[9] + kernel_img_mul_23[10] + kernel_img_mul_23[11] + 
                kernel_img_mul_23[12] + kernel_img_mul_23[13] + kernel_img_mul_23[14] + 
                kernel_img_mul_23[15] + kernel_img_mul_23[16] + kernel_img_mul_23[17] + 
                kernel_img_mul_23[18] + kernel_img_mul_23[19] + kernel_img_mul_23[20] + 
                kernel_img_mul_23[21] + kernel_img_mul_23[22] + kernel_img_mul_23[23] + 
                kernel_img_mul_23[24];
wire  [39:0]  kernel_img_mul_24[0:24];
assign kernel_img_mul_24[0] = layer0[24][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_24[1] = layer0[24][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_24[2] = layer0[24][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_24[3] = layer0[24][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_24[4] = layer0[24][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_24[5] = layer1[24][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_24[6] = layer1[24][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_24[7] = layer1[24][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_24[8] = layer1[24][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_24[9] = layer1[24][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_24[10] = layer2[24][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_24[11] = layer2[24][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_24[12] = layer2[24][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_24[13] = layer2[24][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_24[14] = layer2[24][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_24[15] = layer3[24][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_24[16] = layer3[24][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_24[17] = layer3[24][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_24[18] = layer3[24][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_24[19] = layer3[24][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_24[20] = layer4[24][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_24[21] = layer4[24][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_24[22] = layer4[24][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_24[23] = layer4[24][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_24[24] = layer4[24][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_24 = kernel_img_mul_24[0] + kernel_img_mul_24[1] + kernel_img_mul_24[2] + 
                kernel_img_mul_24[3] + kernel_img_mul_24[4] + kernel_img_mul_24[5] + 
                kernel_img_mul_24[6] + kernel_img_mul_24[7] + kernel_img_mul_24[8] + 
                kernel_img_mul_24[9] + kernel_img_mul_24[10] + kernel_img_mul_24[11] + 
                kernel_img_mul_24[12] + kernel_img_mul_24[13] + kernel_img_mul_24[14] + 
                kernel_img_mul_24[15] + kernel_img_mul_24[16] + kernel_img_mul_24[17] + 
                kernel_img_mul_24[18] + kernel_img_mul_24[19] + kernel_img_mul_24[20] + 
                kernel_img_mul_24[21] + kernel_img_mul_24[22] + kernel_img_mul_24[23] + 
                kernel_img_mul_24[24];
wire  [39:0]  kernel_img_mul_25[0:24];
assign kernel_img_mul_25[0] = layer0[25][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_25[1] = layer0[25][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_25[2] = layer0[25][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_25[3] = layer0[25][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_25[4] = layer0[25][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_25[5] = layer1[25][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_25[6] = layer1[25][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_25[7] = layer1[25][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_25[8] = layer1[25][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_25[9] = layer1[25][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_25[10] = layer2[25][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_25[11] = layer2[25][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_25[12] = layer2[25][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_25[13] = layer2[25][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_25[14] = layer2[25][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_25[15] = layer3[25][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_25[16] = layer3[25][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_25[17] = layer3[25][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_25[18] = layer3[25][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_25[19] = layer3[25][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_25[20] = layer4[25][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_25[21] = layer4[25][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_25[22] = layer4[25][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_25[23] = layer4[25][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_25[24] = layer4[25][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_25 = kernel_img_mul_25[0] + kernel_img_mul_25[1] + kernel_img_mul_25[2] + 
                kernel_img_mul_25[3] + kernel_img_mul_25[4] + kernel_img_mul_25[5] + 
                kernel_img_mul_25[6] + kernel_img_mul_25[7] + kernel_img_mul_25[8] + 
                kernel_img_mul_25[9] + kernel_img_mul_25[10] + kernel_img_mul_25[11] + 
                kernel_img_mul_25[12] + kernel_img_mul_25[13] + kernel_img_mul_25[14] + 
                kernel_img_mul_25[15] + kernel_img_mul_25[16] + kernel_img_mul_25[17] + 
                kernel_img_mul_25[18] + kernel_img_mul_25[19] + kernel_img_mul_25[20] + 
                kernel_img_mul_25[21] + kernel_img_mul_25[22] + kernel_img_mul_25[23] + 
                kernel_img_mul_25[24];
wire  [39:0]  kernel_img_mul_26[0:24];
assign kernel_img_mul_26[0] = layer0[26][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_26[1] = layer0[26][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_26[2] = layer0[26][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_26[3] = layer0[26][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_26[4] = layer0[26][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_26[5] = layer1[26][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_26[6] = layer1[26][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_26[7] = layer1[26][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_26[8] = layer1[26][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_26[9] = layer1[26][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_26[10] = layer2[26][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_26[11] = layer2[26][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_26[12] = layer2[26][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_26[13] = layer2[26][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_26[14] = layer2[26][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_26[15] = layer3[26][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_26[16] = layer3[26][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_26[17] = layer3[26][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_26[18] = layer3[26][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_26[19] = layer3[26][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_26[20] = layer4[26][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_26[21] = layer4[26][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_26[22] = layer4[26][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_26[23] = layer4[26][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_26[24] = layer4[26][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_26 = kernel_img_mul_26[0] + kernel_img_mul_26[1] + kernel_img_mul_26[2] + 
                kernel_img_mul_26[3] + kernel_img_mul_26[4] + kernel_img_mul_26[5] + 
                kernel_img_mul_26[6] + kernel_img_mul_26[7] + kernel_img_mul_26[8] + 
                kernel_img_mul_26[9] + kernel_img_mul_26[10] + kernel_img_mul_26[11] + 
                kernel_img_mul_26[12] + kernel_img_mul_26[13] + kernel_img_mul_26[14] + 
                kernel_img_mul_26[15] + kernel_img_mul_26[16] + kernel_img_mul_26[17] + 
                kernel_img_mul_26[18] + kernel_img_mul_26[19] + kernel_img_mul_26[20] + 
                kernel_img_mul_26[21] + kernel_img_mul_26[22] + kernel_img_mul_26[23] + 
                kernel_img_mul_26[24];
wire  [39:0]  kernel_img_mul_27[0:24];
assign kernel_img_mul_27[0] = layer0[27][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_27[1] = layer0[27][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_27[2] = layer0[27][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_27[3] = layer0[27][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_27[4] = layer0[27][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_27[5] = layer1[27][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_27[6] = layer1[27][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_27[7] = layer1[27][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_27[8] = layer1[27][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_27[9] = layer1[27][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_27[10] = layer2[27][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_27[11] = layer2[27][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_27[12] = layer2[27][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_27[13] = layer2[27][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_27[14] = layer2[27][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_27[15] = layer3[27][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_27[16] = layer3[27][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_27[17] = layer3[27][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_27[18] = layer3[27][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_27[19] = layer3[27][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_27[20] = layer4[27][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_27[21] = layer4[27][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_27[22] = layer4[27][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_27[23] = layer4[27][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_27[24] = layer4[27][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_27 = kernel_img_mul_27[0] + kernel_img_mul_27[1] + kernel_img_mul_27[2] + 
                kernel_img_mul_27[3] + kernel_img_mul_27[4] + kernel_img_mul_27[5] + 
                kernel_img_mul_27[6] + kernel_img_mul_27[7] + kernel_img_mul_27[8] + 
                kernel_img_mul_27[9] + kernel_img_mul_27[10] + kernel_img_mul_27[11] + 
                kernel_img_mul_27[12] + kernel_img_mul_27[13] + kernel_img_mul_27[14] + 
                kernel_img_mul_27[15] + kernel_img_mul_27[16] + kernel_img_mul_27[17] + 
                kernel_img_mul_27[18] + kernel_img_mul_27[19] + kernel_img_mul_27[20] + 
                kernel_img_mul_27[21] + kernel_img_mul_27[22] + kernel_img_mul_27[23] + 
                kernel_img_mul_27[24];
wire  [39:0]  kernel_img_mul_28[0:24];
assign kernel_img_mul_28[0] = layer0[28][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_28[1] = layer0[28][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_28[2] = layer0[28][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_28[3] = layer0[28][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_28[4] = layer0[28][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_28[5] = layer1[28][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_28[6] = layer1[28][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_28[7] = layer1[28][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_28[8] = layer1[28][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_28[9] = layer1[28][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_28[10] = layer2[28][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_28[11] = layer2[28][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_28[12] = layer2[28][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_28[13] = layer2[28][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_28[14] = layer2[28][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_28[15] = layer3[28][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_28[16] = layer3[28][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_28[17] = layer3[28][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_28[18] = layer3[28][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_28[19] = layer3[28][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_28[20] = layer4[28][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_28[21] = layer4[28][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_28[22] = layer4[28][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_28[23] = layer4[28][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_28[24] = layer4[28][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_28 = kernel_img_mul_28[0] + kernel_img_mul_28[1] + kernel_img_mul_28[2] + 
                kernel_img_mul_28[3] + kernel_img_mul_28[4] + kernel_img_mul_28[5] + 
                kernel_img_mul_28[6] + kernel_img_mul_28[7] + kernel_img_mul_28[8] + 
                kernel_img_mul_28[9] + kernel_img_mul_28[10] + kernel_img_mul_28[11] + 
                kernel_img_mul_28[12] + kernel_img_mul_28[13] + kernel_img_mul_28[14] + 
                kernel_img_mul_28[15] + kernel_img_mul_28[16] + kernel_img_mul_28[17] + 
                kernel_img_mul_28[18] + kernel_img_mul_28[19] + kernel_img_mul_28[20] + 
                kernel_img_mul_28[21] + kernel_img_mul_28[22] + kernel_img_mul_28[23] + 
                kernel_img_mul_28[24];
wire  [39:0]  kernel_img_mul_29[0:24];
assign kernel_img_mul_29[0] = layer0[29][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_29[1] = layer0[29][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_29[2] = layer0[29][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_29[3] = layer0[29][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_29[4] = layer0[29][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_29[5] = layer1[29][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_29[6] = layer1[29][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_29[7] = layer1[29][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_29[8] = layer1[29][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_29[9] = layer1[29][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_29[10] = layer2[29][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_29[11] = layer2[29][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_29[12] = layer2[29][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_29[13] = layer2[29][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_29[14] = layer2[29][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_29[15] = layer3[29][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_29[16] = layer3[29][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_29[17] = layer3[29][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_29[18] = layer3[29][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_29[19] = layer3[29][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_29[20] = layer4[29][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_29[21] = layer4[29][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_29[22] = layer4[29][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_29[23] = layer4[29][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_29[24] = layer4[29][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_29 = kernel_img_mul_29[0] + kernel_img_mul_29[1] + kernel_img_mul_29[2] + 
                kernel_img_mul_29[3] + kernel_img_mul_29[4] + kernel_img_mul_29[5] + 
                kernel_img_mul_29[6] + kernel_img_mul_29[7] + kernel_img_mul_29[8] + 
                kernel_img_mul_29[9] + kernel_img_mul_29[10] + kernel_img_mul_29[11] + 
                kernel_img_mul_29[12] + kernel_img_mul_29[13] + kernel_img_mul_29[14] + 
                kernel_img_mul_29[15] + kernel_img_mul_29[16] + kernel_img_mul_29[17] + 
                kernel_img_mul_29[18] + kernel_img_mul_29[19] + kernel_img_mul_29[20] + 
                kernel_img_mul_29[21] + kernel_img_mul_29[22] + kernel_img_mul_29[23] + 
                kernel_img_mul_29[24];
wire  [39:0]  kernel_img_mul_30[0:24];
assign kernel_img_mul_30[0] = layer0[30][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_30[1] = layer0[30][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_30[2] = layer0[30][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_30[3] = layer0[30][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_30[4] = layer0[30][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_30[5] = layer1[30][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_30[6] = layer1[30][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_30[7] = layer1[30][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_30[8] = layer1[30][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_30[9] = layer1[30][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_30[10] = layer2[30][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_30[11] = layer2[30][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_30[12] = layer2[30][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_30[13] = layer2[30][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_30[14] = layer2[30][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_30[15] = layer3[30][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_30[16] = layer3[30][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_30[17] = layer3[30][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_30[18] = layer3[30][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_30[19] = layer3[30][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_30[20] = layer4[30][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_30[21] = layer4[30][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_30[22] = layer4[30][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_30[23] = layer4[30][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_30[24] = layer4[30][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_30 = kernel_img_mul_30[0] + kernel_img_mul_30[1] + kernel_img_mul_30[2] + 
                kernel_img_mul_30[3] + kernel_img_mul_30[4] + kernel_img_mul_30[5] + 
                kernel_img_mul_30[6] + kernel_img_mul_30[7] + kernel_img_mul_30[8] + 
                kernel_img_mul_30[9] + kernel_img_mul_30[10] + kernel_img_mul_30[11] + 
                kernel_img_mul_30[12] + kernel_img_mul_30[13] + kernel_img_mul_30[14] + 
                kernel_img_mul_30[15] + kernel_img_mul_30[16] + kernel_img_mul_30[17] + 
                kernel_img_mul_30[18] + kernel_img_mul_30[19] + kernel_img_mul_30[20] + 
                kernel_img_mul_30[21] + kernel_img_mul_30[22] + kernel_img_mul_30[23] + 
                kernel_img_mul_30[24];
wire  [39:0]  kernel_img_mul_31[0:24];
assign kernel_img_mul_31[0] = layer0[31][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_31[1] = layer0[31][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_31[2] = layer0[31][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_31[3] = layer0[31][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_31[4] = layer0[31][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_31[5] = layer1[31][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_31[6] = layer1[31][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_31[7] = layer1[31][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_31[8] = layer1[31][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_31[9] = layer1[31][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_31[10] = layer2[31][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_31[11] = layer2[31][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_31[12] = layer2[31][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_31[13] = layer2[31][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_31[14] = layer2[31][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_31[15] = layer3[31][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_31[16] = layer3[31][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_31[17] = layer3[31][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_31[18] = layer3[31][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_31[19] = layer3[31][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_31[20] = layer4[31][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_31[21] = layer4[31][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_31[22] = layer4[31][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_31[23] = layer4[31][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_31[24] = layer4[31][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_31 = kernel_img_mul_31[0] + kernel_img_mul_31[1] + kernel_img_mul_31[2] + 
                kernel_img_mul_31[3] + kernel_img_mul_31[4] + kernel_img_mul_31[5] + 
                kernel_img_mul_31[6] + kernel_img_mul_31[7] + kernel_img_mul_31[8] + 
                kernel_img_mul_31[9] + kernel_img_mul_31[10] + kernel_img_mul_31[11] + 
                kernel_img_mul_31[12] + kernel_img_mul_31[13] + kernel_img_mul_31[14] + 
                kernel_img_mul_31[15] + kernel_img_mul_31[16] + kernel_img_mul_31[17] + 
                kernel_img_mul_31[18] + kernel_img_mul_31[19] + kernel_img_mul_31[20] + 
                kernel_img_mul_31[21] + kernel_img_mul_31[22] + kernel_img_mul_31[23] + 
                kernel_img_mul_31[24];
wire  [39:0]  kernel_img_mul_32[0:24];
assign kernel_img_mul_32[0] = layer0[32][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_32[1] = layer0[32][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_32[2] = layer0[32][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_32[3] = layer0[32][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_32[4] = layer0[32][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_32[5] = layer1[32][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_32[6] = layer1[32][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_32[7] = layer1[32][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_32[8] = layer1[32][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_32[9] = layer1[32][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_32[10] = layer2[32][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_32[11] = layer2[32][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_32[12] = layer2[32][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_32[13] = layer2[32][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_32[14] = layer2[32][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_32[15] = layer3[32][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_32[16] = layer3[32][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_32[17] = layer3[32][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_32[18] = layer3[32][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_32[19] = layer3[32][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_32[20] = layer4[32][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_32[21] = layer4[32][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_32[22] = layer4[32][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_32[23] = layer4[32][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_32[24] = layer4[32][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_32 = kernel_img_mul_32[0] + kernel_img_mul_32[1] + kernel_img_mul_32[2] + 
                kernel_img_mul_32[3] + kernel_img_mul_32[4] + kernel_img_mul_32[5] + 
                kernel_img_mul_32[6] + kernel_img_mul_32[7] + kernel_img_mul_32[8] + 
                kernel_img_mul_32[9] + kernel_img_mul_32[10] + kernel_img_mul_32[11] + 
                kernel_img_mul_32[12] + kernel_img_mul_32[13] + kernel_img_mul_32[14] + 
                kernel_img_mul_32[15] + kernel_img_mul_32[16] + kernel_img_mul_32[17] + 
                kernel_img_mul_32[18] + kernel_img_mul_32[19] + kernel_img_mul_32[20] + 
                kernel_img_mul_32[21] + kernel_img_mul_32[22] + kernel_img_mul_32[23] + 
                kernel_img_mul_32[24];
wire  [39:0]  kernel_img_mul_33[0:24];
assign kernel_img_mul_33[0] = layer0[33][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_33[1] = layer0[33][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_33[2] = layer0[33][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_33[3] = layer0[33][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_33[4] = layer0[33][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_33[5] = layer1[33][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_33[6] = layer1[33][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_33[7] = layer1[33][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_33[8] = layer1[33][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_33[9] = layer1[33][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_33[10] = layer2[33][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_33[11] = layer2[33][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_33[12] = layer2[33][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_33[13] = layer2[33][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_33[14] = layer2[33][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_33[15] = layer3[33][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_33[16] = layer3[33][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_33[17] = layer3[33][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_33[18] = layer3[33][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_33[19] = layer3[33][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_33[20] = layer4[33][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_33[21] = layer4[33][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_33[22] = layer4[33][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_33[23] = layer4[33][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_33[24] = layer4[33][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_33 = kernel_img_mul_33[0] + kernel_img_mul_33[1] + kernel_img_mul_33[2] + 
                kernel_img_mul_33[3] + kernel_img_mul_33[4] + kernel_img_mul_33[5] + 
                kernel_img_mul_33[6] + kernel_img_mul_33[7] + kernel_img_mul_33[8] + 
                kernel_img_mul_33[9] + kernel_img_mul_33[10] + kernel_img_mul_33[11] + 
                kernel_img_mul_33[12] + kernel_img_mul_33[13] + kernel_img_mul_33[14] + 
                kernel_img_mul_33[15] + kernel_img_mul_33[16] + kernel_img_mul_33[17] + 
                kernel_img_mul_33[18] + kernel_img_mul_33[19] + kernel_img_mul_33[20] + 
                kernel_img_mul_33[21] + kernel_img_mul_33[22] + kernel_img_mul_33[23] + 
                kernel_img_mul_33[24];
wire  [39:0]  kernel_img_mul_34[0:24];
assign kernel_img_mul_34[0] = layer0[34][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_34[1] = layer0[34][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_34[2] = layer0[34][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_34[3] = layer0[34][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_34[4] = layer0[34][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_34[5] = layer1[34][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_34[6] = layer1[34][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_34[7] = layer1[34][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_34[8] = layer1[34][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_34[9] = layer1[34][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_34[10] = layer2[34][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_34[11] = layer2[34][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_34[12] = layer2[34][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_34[13] = layer2[34][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_34[14] = layer2[34][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_34[15] = layer3[34][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_34[16] = layer3[34][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_34[17] = layer3[34][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_34[18] = layer3[34][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_34[19] = layer3[34][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_34[20] = layer4[34][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_34[21] = layer4[34][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_34[22] = layer4[34][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_34[23] = layer4[34][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_34[24] = layer4[34][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_34 = kernel_img_mul_34[0] + kernel_img_mul_34[1] + kernel_img_mul_34[2] + 
                kernel_img_mul_34[3] + kernel_img_mul_34[4] + kernel_img_mul_34[5] + 
                kernel_img_mul_34[6] + kernel_img_mul_34[7] + kernel_img_mul_34[8] + 
                kernel_img_mul_34[9] + kernel_img_mul_34[10] + kernel_img_mul_34[11] + 
                kernel_img_mul_34[12] + kernel_img_mul_34[13] + kernel_img_mul_34[14] + 
                kernel_img_mul_34[15] + kernel_img_mul_34[16] + kernel_img_mul_34[17] + 
                kernel_img_mul_34[18] + kernel_img_mul_34[19] + kernel_img_mul_34[20] + 
                kernel_img_mul_34[21] + kernel_img_mul_34[22] + kernel_img_mul_34[23] + 
                kernel_img_mul_34[24];
wire  [39:0]  kernel_img_mul_35[0:24];
assign kernel_img_mul_35[0] = layer0[35][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_35[1] = layer0[35][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_35[2] = layer0[35][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_35[3] = layer0[35][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_35[4] = layer0[35][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_35[5] = layer1[35][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_35[6] = layer1[35][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_35[7] = layer1[35][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_35[8] = layer1[35][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_35[9] = layer1[35][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_35[10] = layer2[35][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_35[11] = layer2[35][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_35[12] = layer2[35][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_35[13] = layer2[35][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_35[14] = layer2[35][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_35[15] = layer3[35][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_35[16] = layer3[35][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_35[17] = layer3[35][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_35[18] = layer3[35][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_35[19] = layer3[35][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_35[20] = layer4[35][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_35[21] = layer4[35][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_35[22] = layer4[35][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_35[23] = layer4[35][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_35[24] = layer4[35][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_35 = kernel_img_mul_35[0] + kernel_img_mul_35[1] + kernel_img_mul_35[2] + 
                kernel_img_mul_35[3] + kernel_img_mul_35[4] + kernel_img_mul_35[5] + 
                kernel_img_mul_35[6] + kernel_img_mul_35[7] + kernel_img_mul_35[8] + 
                kernel_img_mul_35[9] + kernel_img_mul_35[10] + kernel_img_mul_35[11] + 
                kernel_img_mul_35[12] + kernel_img_mul_35[13] + kernel_img_mul_35[14] + 
                kernel_img_mul_35[15] + kernel_img_mul_35[16] + kernel_img_mul_35[17] + 
                kernel_img_mul_35[18] + kernel_img_mul_35[19] + kernel_img_mul_35[20] + 
                kernel_img_mul_35[21] + kernel_img_mul_35[22] + kernel_img_mul_35[23] + 
                kernel_img_mul_35[24];
wire  [39:0]  kernel_img_mul_36[0:24];
assign kernel_img_mul_36[0] = layer0[36][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_36[1] = layer0[36][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_36[2] = layer0[36][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_36[3] = layer0[36][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_36[4] = layer0[36][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_36[5] = layer1[36][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_36[6] = layer1[36][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_36[7] = layer1[36][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_36[8] = layer1[36][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_36[9] = layer1[36][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_36[10] = layer2[36][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_36[11] = layer2[36][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_36[12] = layer2[36][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_36[13] = layer2[36][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_36[14] = layer2[36][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_36[15] = layer3[36][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_36[16] = layer3[36][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_36[17] = layer3[36][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_36[18] = layer3[36][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_36[19] = layer3[36][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_36[20] = layer4[36][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_36[21] = layer4[36][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_36[22] = layer4[36][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_36[23] = layer4[36][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_36[24] = layer4[36][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_36 = kernel_img_mul_36[0] + kernel_img_mul_36[1] + kernel_img_mul_36[2] + 
                kernel_img_mul_36[3] + kernel_img_mul_36[4] + kernel_img_mul_36[5] + 
                kernel_img_mul_36[6] + kernel_img_mul_36[7] + kernel_img_mul_36[8] + 
                kernel_img_mul_36[9] + kernel_img_mul_36[10] + kernel_img_mul_36[11] + 
                kernel_img_mul_36[12] + kernel_img_mul_36[13] + kernel_img_mul_36[14] + 
                kernel_img_mul_36[15] + kernel_img_mul_36[16] + kernel_img_mul_36[17] + 
                kernel_img_mul_36[18] + kernel_img_mul_36[19] + kernel_img_mul_36[20] + 
                kernel_img_mul_36[21] + kernel_img_mul_36[22] + kernel_img_mul_36[23] + 
                kernel_img_mul_36[24];
wire  [39:0]  kernel_img_mul_37[0:24];
assign kernel_img_mul_37[0] = layer0[37][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_37[1] = layer0[37][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_37[2] = layer0[37][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_37[3] = layer0[37][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_37[4] = layer0[37][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_37[5] = layer1[37][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_37[6] = layer1[37][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_37[7] = layer1[37][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_37[8] = layer1[37][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_37[9] = layer1[37][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_37[10] = layer2[37][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_37[11] = layer2[37][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_37[12] = layer2[37][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_37[13] = layer2[37][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_37[14] = layer2[37][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_37[15] = layer3[37][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_37[16] = layer3[37][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_37[17] = layer3[37][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_37[18] = layer3[37][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_37[19] = layer3[37][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_37[20] = layer4[37][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_37[21] = layer4[37][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_37[22] = layer4[37][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_37[23] = layer4[37][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_37[24] = layer4[37][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_37 = kernel_img_mul_37[0] + kernel_img_mul_37[1] + kernel_img_mul_37[2] + 
                kernel_img_mul_37[3] + kernel_img_mul_37[4] + kernel_img_mul_37[5] + 
                kernel_img_mul_37[6] + kernel_img_mul_37[7] + kernel_img_mul_37[8] + 
                kernel_img_mul_37[9] + kernel_img_mul_37[10] + kernel_img_mul_37[11] + 
                kernel_img_mul_37[12] + kernel_img_mul_37[13] + kernel_img_mul_37[14] + 
                kernel_img_mul_37[15] + kernel_img_mul_37[16] + kernel_img_mul_37[17] + 
                kernel_img_mul_37[18] + kernel_img_mul_37[19] + kernel_img_mul_37[20] + 
                kernel_img_mul_37[21] + kernel_img_mul_37[22] + kernel_img_mul_37[23] + 
                kernel_img_mul_37[24];
wire  [39:0]  kernel_img_mul_38[0:24];
assign kernel_img_mul_38[0] = layer0[38][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_38[1] = layer0[38][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_38[2] = layer0[38][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_38[3] = layer0[38][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_38[4] = layer0[38][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_38[5] = layer1[38][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_38[6] = layer1[38][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_38[7] = layer1[38][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_38[8] = layer1[38][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_38[9] = layer1[38][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_38[10] = layer2[38][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_38[11] = layer2[38][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_38[12] = layer2[38][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_38[13] = layer2[38][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_38[14] = layer2[38][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_38[15] = layer3[38][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_38[16] = layer3[38][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_38[17] = layer3[38][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_38[18] = layer3[38][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_38[19] = layer3[38][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_38[20] = layer4[38][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_38[21] = layer4[38][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_38[22] = layer4[38][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_38[23] = layer4[38][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_38[24] = layer4[38][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_38 = kernel_img_mul_38[0] + kernel_img_mul_38[1] + kernel_img_mul_38[2] + 
                kernel_img_mul_38[3] + kernel_img_mul_38[4] + kernel_img_mul_38[5] + 
                kernel_img_mul_38[6] + kernel_img_mul_38[7] + kernel_img_mul_38[8] + 
                kernel_img_mul_38[9] + kernel_img_mul_38[10] + kernel_img_mul_38[11] + 
                kernel_img_mul_38[12] + kernel_img_mul_38[13] + kernel_img_mul_38[14] + 
                kernel_img_mul_38[15] + kernel_img_mul_38[16] + kernel_img_mul_38[17] + 
                kernel_img_mul_38[18] + kernel_img_mul_38[19] + kernel_img_mul_38[20] + 
                kernel_img_mul_38[21] + kernel_img_mul_38[22] + kernel_img_mul_38[23] + 
                kernel_img_mul_38[24];
wire  [39:0]  kernel_img_mul_39[0:24];
assign kernel_img_mul_39[0] = layer0[39][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_39[1] = layer0[39][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_39[2] = layer0[39][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_39[3] = layer0[39][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_39[4] = layer0[39][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_39[5] = layer1[39][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_39[6] = layer1[39][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_39[7] = layer1[39][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_39[8] = layer1[39][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_39[9] = layer1[39][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_39[10] = layer2[39][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_39[11] = layer2[39][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_39[12] = layer2[39][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_39[13] = layer2[39][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_39[14] = layer2[39][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_39[15] = layer3[39][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_39[16] = layer3[39][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_39[17] = layer3[39][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_39[18] = layer3[39][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_39[19] = layer3[39][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_39[20] = layer4[39][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_39[21] = layer4[39][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_39[22] = layer4[39][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_39[23] = layer4[39][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_39[24] = layer4[39][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_39 = kernel_img_mul_39[0] + kernel_img_mul_39[1] + kernel_img_mul_39[2] + 
                kernel_img_mul_39[3] + kernel_img_mul_39[4] + kernel_img_mul_39[5] + 
                kernel_img_mul_39[6] + kernel_img_mul_39[7] + kernel_img_mul_39[8] + 
                kernel_img_mul_39[9] + kernel_img_mul_39[10] + kernel_img_mul_39[11] + 
                kernel_img_mul_39[12] + kernel_img_mul_39[13] + kernel_img_mul_39[14] + 
                kernel_img_mul_39[15] + kernel_img_mul_39[16] + kernel_img_mul_39[17] + 
                kernel_img_mul_39[18] + kernel_img_mul_39[19] + kernel_img_mul_39[20] + 
                kernel_img_mul_39[21] + kernel_img_mul_39[22] + kernel_img_mul_39[23] + 
                kernel_img_mul_39[24];
wire  [39:0]  kernel_img_mul_40[0:24];
assign kernel_img_mul_40[0] = layer0[40][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_40[1] = layer0[40][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_40[2] = layer0[40][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_40[3] = layer0[40][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_40[4] = layer0[40][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_40[5] = layer1[40][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_40[6] = layer1[40][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_40[7] = layer1[40][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_40[8] = layer1[40][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_40[9] = layer1[40][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_40[10] = layer2[40][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_40[11] = layer2[40][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_40[12] = layer2[40][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_40[13] = layer2[40][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_40[14] = layer2[40][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_40[15] = layer3[40][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_40[16] = layer3[40][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_40[17] = layer3[40][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_40[18] = layer3[40][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_40[19] = layer3[40][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_40[20] = layer4[40][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_40[21] = layer4[40][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_40[22] = layer4[40][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_40[23] = layer4[40][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_40[24] = layer4[40][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_40 = kernel_img_mul_40[0] + kernel_img_mul_40[1] + kernel_img_mul_40[2] + 
                kernel_img_mul_40[3] + kernel_img_mul_40[4] + kernel_img_mul_40[5] + 
                kernel_img_mul_40[6] + kernel_img_mul_40[7] + kernel_img_mul_40[8] + 
                kernel_img_mul_40[9] + kernel_img_mul_40[10] + kernel_img_mul_40[11] + 
                kernel_img_mul_40[12] + kernel_img_mul_40[13] + kernel_img_mul_40[14] + 
                kernel_img_mul_40[15] + kernel_img_mul_40[16] + kernel_img_mul_40[17] + 
                kernel_img_mul_40[18] + kernel_img_mul_40[19] + kernel_img_mul_40[20] + 
                kernel_img_mul_40[21] + kernel_img_mul_40[22] + kernel_img_mul_40[23] + 
                kernel_img_mul_40[24];
wire  [39:0]  kernel_img_mul_41[0:24];
assign kernel_img_mul_41[0] = layer0[41][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_41[1] = layer0[41][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_41[2] = layer0[41][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_41[3] = layer0[41][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_41[4] = layer0[41][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_41[5] = layer1[41][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_41[6] = layer1[41][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_41[7] = layer1[41][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_41[8] = layer1[41][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_41[9] = layer1[41][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_41[10] = layer2[41][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_41[11] = layer2[41][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_41[12] = layer2[41][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_41[13] = layer2[41][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_41[14] = layer2[41][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_41[15] = layer3[41][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_41[16] = layer3[41][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_41[17] = layer3[41][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_41[18] = layer3[41][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_41[19] = layer3[41][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_41[20] = layer4[41][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_41[21] = layer4[41][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_41[22] = layer4[41][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_41[23] = layer4[41][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_41[24] = layer4[41][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_41 = kernel_img_mul_41[0] + kernel_img_mul_41[1] + kernel_img_mul_41[2] + 
                kernel_img_mul_41[3] + kernel_img_mul_41[4] + kernel_img_mul_41[5] + 
                kernel_img_mul_41[6] + kernel_img_mul_41[7] + kernel_img_mul_41[8] + 
                kernel_img_mul_41[9] + kernel_img_mul_41[10] + kernel_img_mul_41[11] + 
                kernel_img_mul_41[12] + kernel_img_mul_41[13] + kernel_img_mul_41[14] + 
                kernel_img_mul_41[15] + kernel_img_mul_41[16] + kernel_img_mul_41[17] + 
                kernel_img_mul_41[18] + kernel_img_mul_41[19] + kernel_img_mul_41[20] + 
                kernel_img_mul_41[21] + kernel_img_mul_41[22] + kernel_img_mul_41[23] + 
                kernel_img_mul_41[24];
wire  [39:0]  kernel_img_mul_42[0:24];
assign kernel_img_mul_42[0] = layer0[42][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_42[1] = layer0[42][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_42[2] = layer0[42][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_42[3] = layer0[42][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_42[4] = layer0[42][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_42[5] = layer1[42][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_42[6] = layer1[42][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_42[7] = layer1[42][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_42[8] = layer1[42][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_42[9] = layer1[42][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_42[10] = layer2[42][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_42[11] = layer2[42][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_42[12] = layer2[42][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_42[13] = layer2[42][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_42[14] = layer2[42][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_42[15] = layer3[42][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_42[16] = layer3[42][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_42[17] = layer3[42][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_42[18] = layer3[42][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_42[19] = layer3[42][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_42[20] = layer4[42][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_42[21] = layer4[42][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_42[22] = layer4[42][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_42[23] = layer4[42][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_42[24] = layer4[42][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_42 = kernel_img_mul_42[0] + kernel_img_mul_42[1] + kernel_img_mul_42[2] + 
                kernel_img_mul_42[3] + kernel_img_mul_42[4] + kernel_img_mul_42[5] + 
                kernel_img_mul_42[6] + kernel_img_mul_42[7] + kernel_img_mul_42[8] + 
                kernel_img_mul_42[9] + kernel_img_mul_42[10] + kernel_img_mul_42[11] + 
                kernel_img_mul_42[12] + kernel_img_mul_42[13] + kernel_img_mul_42[14] + 
                kernel_img_mul_42[15] + kernel_img_mul_42[16] + kernel_img_mul_42[17] + 
                kernel_img_mul_42[18] + kernel_img_mul_42[19] + kernel_img_mul_42[20] + 
                kernel_img_mul_42[21] + kernel_img_mul_42[22] + kernel_img_mul_42[23] + 
                kernel_img_mul_42[24];
wire  [39:0]  kernel_img_mul_43[0:24];
assign kernel_img_mul_43[0] = layer0[43][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_43[1] = layer0[43][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_43[2] = layer0[43][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_43[3] = layer0[43][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_43[4] = layer0[43][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_43[5] = layer1[43][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_43[6] = layer1[43][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_43[7] = layer1[43][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_43[8] = layer1[43][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_43[9] = layer1[43][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_43[10] = layer2[43][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_43[11] = layer2[43][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_43[12] = layer2[43][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_43[13] = layer2[43][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_43[14] = layer2[43][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_43[15] = layer3[43][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_43[16] = layer3[43][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_43[17] = layer3[43][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_43[18] = layer3[43][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_43[19] = layer3[43][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_43[20] = layer4[43][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_43[21] = layer4[43][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_43[22] = layer4[43][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_43[23] = layer4[43][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_43[24] = layer4[43][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_43 = kernel_img_mul_43[0] + kernel_img_mul_43[1] + kernel_img_mul_43[2] + 
                kernel_img_mul_43[3] + kernel_img_mul_43[4] + kernel_img_mul_43[5] + 
                kernel_img_mul_43[6] + kernel_img_mul_43[7] + kernel_img_mul_43[8] + 
                kernel_img_mul_43[9] + kernel_img_mul_43[10] + kernel_img_mul_43[11] + 
                kernel_img_mul_43[12] + kernel_img_mul_43[13] + kernel_img_mul_43[14] + 
                kernel_img_mul_43[15] + kernel_img_mul_43[16] + kernel_img_mul_43[17] + 
                kernel_img_mul_43[18] + kernel_img_mul_43[19] + kernel_img_mul_43[20] + 
                kernel_img_mul_43[21] + kernel_img_mul_43[22] + kernel_img_mul_43[23] + 
                kernel_img_mul_43[24];
wire  [39:0]  kernel_img_mul_44[0:24];
assign kernel_img_mul_44[0] = layer0[44][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_44[1] = layer0[44][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_44[2] = layer0[44][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_44[3] = layer0[44][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_44[4] = layer0[44][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_44[5] = layer1[44][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_44[6] = layer1[44][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_44[7] = layer1[44][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_44[8] = layer1[44][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_44[9] = layer1[44][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_44[10] = layer2[44][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_44[11] = layer2[44][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_44[12] = layer2[44][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_44[13] = layer2[44][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_44[14] = layer2[44][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_44[15] = layer3[44][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_44[16] = layer3[44][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_44[17] = layer3[44][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_44[18] = layer3[44][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_44[19] = layer3[44][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_44[20] = layer4[44][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_44[21] = layer4[44][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_44[22] = layer4[44][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_44[23] = layer4[44][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_44[24] = layer4[44][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_44 = kernel_img_mul_44[0] + kernel_img_mul_44[1] + kernel_img_mul_44[2] + 
                kernel_img_mul_44[3] + kernel_img_mul_44[4] + kernel_img_mul_44[5] + 
                kernel_img_mul_44[6] + kernel_img_mul_44[7] + kernel_img_mul_44[8] + 
                kernel_img_mul_44[9] + kernel_img_mul_44[10] + kernel_img_mul_44[11] + 
                kernel_img_mul_44[12] + kernel_img_mul_44[13] + kernel_img_mul_44[14] + 
                kernel_img_mul_44[15] + kernel_img_mul_44[16] + kernel_img_mul_44[17] + 
                kernel_img_mul_44[18] + kernel_img_mul_44[19] + kernel_img_mul_44[20] + 
                kernel_img_mul_44[21] + kernel_img_mul_44[22] + kernel_img_mul_44[23] + 
                kernel_img_mul_44[24];
wire  [39:0]  kernel_img_mul_45[0:24];
assign kernel_img_mul_45[0] = layer0[45][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_45[1] = layer0[45][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_45[2] = layer0[45][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_45[3] = layer0[45][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_45[4] = layer0[45][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_45[5] = layer1[45][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_45[6] = layer1[45][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_45[7] = layer1[45][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_45[8] = layer1[45][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_45[9] = layer1[45][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_45[10] = layer2[45][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_45[11] = layer2[45][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_45[12] = layer2[45][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_45[13] = layer2[45][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_45[14] = layer2[45][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_45[15] = layer3[45][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_45[16] = layer3[45][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_45[17] = layer3[45][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_45[18] = layer3[45][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_45[19] = layer3[45][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_45[20] = layer4[45][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_45[21] = layer4[45][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_45[22] = layer4[45][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_45[23] = layer4[45][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_45[24] = layer4[45][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_45 = kernel_img_mul_45[0] + kernel_img_mul_45[1] + kernel_img_mul_45[2] + 
                kernel_img_mul_45[3] + kernel_img_mul_45[4] + kernel_img_mul_45[5] + 
                kernel_img_mul_45[6] + kernel_img_mul_45[7] + kernel_img_mul_45[8] + 
                kernel_img_mul_45[9] + kernel_img_mul_45[10] + kernel_img_mul_45[11] + 
                kernel_img_mul_45[12] + kernel_img_mul_45[13] + kernel_img_mul_45[14] + 
                kernel_img_mul_45[15] + kernel_img_mul_45[16] + kernel_img_mul_45[17] + 
                kernel_img_mul_45[18] + kernel_img_mul_45[19] + kernel_img_mul_45[20] + 
                kernel_img_mul_45[21] + kernel_img_mul_45[22] + kernel_img_mul_45[23] + 
                kernel_img_mul_45[24];
wire  [39:0]  kernel_img_mul_46[0:24];
assign kernel_img_mul_46[0] = layer0[46][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_46[1] = layer0[46][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_46[2] = layer0[46][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_46[3] = layer0[46][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_46[4] = layer0[46][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_46[5] = layer1[46][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_46[6] = layer1[46][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_46[7] = layer1[46][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_46[8] = layer1[46][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_46[9] = layer1[46][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_46[10] = layer2[46][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_46[11] = layer2[46][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_46[12] = layer2[46][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_46[13] = layer2[46][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_46[14] = layer2[46][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_46[15] = layer3[46][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_46[16] = layer3[46][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_46[17] = layer3[46][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_46[18] = layer3[46][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_46[19] = layer3[46][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_46[20] = layer4[46][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_46[21] = layer4[46][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_46[22] = layer4[46][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_46[23] = layer4[46][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_46[24] = layer4[46][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_46 = kernel_img_mul_46[0] + kernel_img_mul_46[1] + kernel_img_mul_46[2] + 
                kernel_img_mul_46[3] + kernel_img_mul_46[4] + kernel_img_mul_46[5] + 
                kernel_img_mul_46[6] + kernel_img_mul_46[7] + kernel_img_mul_46[8] + 
                kernel_img_mul_46[9] + kernel_img_mul_46[10] + kernel_img_mul_46[11] + 
                kernel_img_mul_46[12] + kernel_img_mul_46[13] + kernel_img_mul_46[14] + 
                kernel_img_mul_46[15] + kernel_img_mul_46[16] + kernel_img_mul_46[17] + 
                kernel_img_mul_46[18] + kernel_img_mul_46[19] + kernel_img_mul_46[20] + 
                kernel_img_mul_46[21] + kernel_img_mul_46[22] + kernel_img_mul_46[23] + 
                kernel_img_mul_46[24];
wire  [39:0]  kernel_img_mul_47[0:24];
assign kernel_img_mul_47[0] = layer0[47][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_47[1] = layer0[47][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_47[2] = layer0[47][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_47[3] = layer0[47][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_47[4] = layer0[47][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_47[5] = layer1[47][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_47[6] = layer1[47][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_47[7] = layer1[47][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_47[8] = layer1[47][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_47[9] = layer1[47][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_47[10] = layer2[47][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_47[11] = layer2[47][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_47[12] = layer2[47][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_47[13] = layer2[47][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_47[14] = layer2[47][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_47[15] = layer3[47][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_47[16] = layer3[47][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_47[17] = layer3[47][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_47[18] = layer3[47][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_47[19] = layer3[47][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_47[20] = layer4[47][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_47[21] = layer4[47][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_47[22] = layer4[47][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_47[23] = layer4[47][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_47[24] = layer4[47][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_47 = kernel_img_mul_47[0] + kernel_img_mul_47[1] + kernel_img_mul_47[2] + 
                kernel_img_mul_47[3] + kernel_img_mul_47[4] + kernel_img_mul_47[5] + 
                kernel_img_mul_47[6] + kernel_img_mul_47[7] + kernel_img_mul_47[8] + 
                kernel_img_mul_47[9] + kernel_img_mul_47[10] + kernel_img_mul_47[11] + 
                kernel_img_mul_47[12] + kernel_img_mul_47[13] + kernel_img_mul_47[14] + 
                kernel_img_mul_47[15] + kernel_img_mul_47[16] + kernel_img_mul_47[17] + 
                kernel_img_mul_47[18] + kernel_img_mul_47[19] + kernel_img_mul_47[20] + 
                kernel_img_mul_47[21] + kernel_img_mul_47[22] + kernel_img_mul_47[23] + 
                kernel_img_mul_47[24];
wire  [39:0]  kernel_img_mul_48[0:24];
assign kernel_img_mul_48[0] = layer0[48][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_48[1] = layer0[48][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_48[2] = layer0[48][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_48[3] = layer0[48][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_48[4] = layer0[48][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_48[5] = layer1[48][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_48[6] = layer1[48][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_48[7] = layer1[48][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_48[8] = layer1[48][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_48[9] = layer1[48][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_48[10] = layer2[48][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_48[11] = layer2[48][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_48[12] = layer2[48][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_48[13] = layer2[48][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_48[14] = layer2[48][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_48[15] = layer3[48][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_48[16] = layer3[48][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_48[17] = layer3[48][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_48[18] = layer3[48][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_48[19] = layer3[48][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_48[20] = layer4[48][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_48[21] = layer4[48][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_48[22] = layer4[48][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_48[23] = layer4[48][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_48[24] = layer4[48][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_48 = kernel_img_mul_48[0] + kernel_img_mul_48[1] + kernel_img_mul_48[2] + 
                kernel_img_mul_48[3] + kernel_img_mul_48[4] + kernel_img_mul_48[5] + 
                kernel_img_mul_48[6] + kernel_img_mul_48[7] + kernel_img_mul_48[8] + 
                kernel_img_mul_48[9] + kernel_img_mul_48[10] + kernel_img_mul_48[11] + 
                kernel_img_mul_48[12] + kernel_img_mul_48[13] + kernel_img_mul_48[14] + 
                kernel_img_mul_48[15] + kernel_img_mul_48[16] + kernel_img_mul_48[17] + 
                kernel_img_mul_48[18] + kernel_img_mul_48[19] + kernel_img_mul_48[20] + 
                kernel_img_mul_48[21] + kernel_img_mul_48[22] + kernel_img_mul_48[23] + 
                kernel_img_mul_48[24];
wire  [39:0]  kernel_img_mul_49[0:24];
assign kernel_img_mul_49[0] = layer0[49][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_49[1] = layer0[49][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_49[2] = layer0[49][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_49[3] = layer0[49][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_49[4] = layer0[49][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_49[5] = layer1[49][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_49[6] = layer1[49][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_49[7] = layer1[49][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_49[8] = layer1[49][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_49[9] = layer1[49][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_49[10] = layer2[49][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_49[11] = layer2[49][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_49[12] = layer2[49][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_49[13] = layer2[49][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_49[14] = layer2[49][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_49[15] = layer3[49][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_49[16] = layer3[49][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_49[17] = layer3[49][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_49[18] = layer3[49][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_49[19] = layer3[49][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_49[20] = layer4[49][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_49[21] = layer4[49][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_49[22] = layer4[49][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_49[23] = layer4[49][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_49[24] = layer4[49][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_49 = kernel_img_mul_49[0] + kernel_img_mul_49[1] + kernel_img_mul_49[2] + 
                kernel_img_mul_49[3] + kernel_img_mul_49[4] + kernel_img_mul_49[5] + 
                kernel_img_mul_49[6] + kernel_img_mul_49[7] + kernel_img_mul_49[8] + 
                kernel_img_mul_49[9] + kernel_img_mul_49[10] + kernel_img_mul_49[11] + 
                kernel_img_mul_49[12] + kernel_img_mul_49[13] + kernel_img_mul_49[14] + 
                kernel_img_mul_49[15] + kernel_img_mul_49[16] + kernel_img_mul_49[17] + 
                kernel_img_mul_49[18] + kernel_img_mul_49[19] + kernel_img_mul_49[20] + 
                kernel_img_mul_49[21] + kernel_img_mul_49[22] + kernel_img_mul_49[23] + 
                kernel_img_mul_49[24];
wire  [39:0]  kernel_img_mul_50[0:24];
assign kernel_img_mul_50[0] = layer0[50][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_50[1] = layer0[50][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_50[2] = layer0[50][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_50[3] = layer0[50][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_50[4] = layer0[50][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_50[5] = layer1[50][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_50[6] = layer1[50][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_50[7] = layer1[50][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_50[8] = layer1[50][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_50[9] = layer1[50][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_50[10] = layer2[50][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_50[11] = layer2[50][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_50[12] = layer2[50][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_50[13] = layer2[50][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_50[14] = layer2[50][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_50[15] = layer3[50][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_50[16] = layer3[50][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_50[17] = layer3[50][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_50[18] = layer3[50][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_50[19] = layer3[50][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_50[20] = layer4[50][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_50[21] = layer4[50][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_50[22] = layer4[50][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_50[23] = layer4[50][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_50[24] = layer4[50][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_50 = kernel_img_mul_50[0] + kernel_img_mul_50[1] + kernel_img_mul_50[2] + 
                kernel_img_mul_50[3] + kernel_img_mul_50[4] + kernel_img_mul_50[5] + 
                kernel_img_mul_50[6] + kernel_img_mul_50[7] + kernel_img_mul_50[8] + 
                kernel_img_mul_50[9] + kernel_img_mul_50[10] + kernel_img_mul_50[11] + 
                kernel_img_mul_50[12] + kernel_img_mul_50[13] + kernel_img_mul_50[14] + 
                kernel_img_mul_50[15] + kernel_img_mul_50[16] + kernel_img_mul_50[17] + 
                kernel_img_mul_50[18] + kernel_img_mul_50[19] + kernel_img_mul_50[20] + 
                kernel_img_mul_50[21] + kernel_img_mul_50[22] + kernel_img_mul_50[23] + 
                kernel_img_mul_50[24];
wire  [39:0]  kernel_img_mul_51[0:24];
assign kernel_img_mul_51[0] = layer0[51][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_51[1] = layer0[51][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_51[2] = layer0[51][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_51[3] = layer0[51][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_51[4] = layer0[51][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_51[5] = layer1[51][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_51[6] = layer1[51][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_51[7] = layer1[51][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_51[8] = layer1[51][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_51[9] = layer1[51][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_51[10] = layer2[51][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_51[11] = layer2[51][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_51[12] = layer2[51][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_51[13] = layer2[51][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_51[14] = layer2[51][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_51[15] = layer3[51][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_51[16] = layer3[51][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_51[17] = layer3[51][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_51[18] = layer3[51][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_51[19] = layer3[51][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_51[20] = layer4[51][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_51[21] = layer4[51][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_51[22] = layer4[51][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_51[23] = layer4[51][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_51[24] = layer4[51][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_51 = kernel_img_mul_51[0] + kernel_img_mul_51[1] + kernel_img_mul_51[2] + 
                kernel_img_mul_51[3] + kernel_img_mul_51[4] + kernel_img_mul_51[5] + 
                kernel_img_mul_51[6] + kernel_img_mul_51[7] + kernel_img_mul_51[8] + 
                kernel_img_mul_51[9] + kernel_img_mul_51[10] + kernel_img_mul_51[11] + 
                kernel_img_mul_51[12] + kernel_img_mul_51[13] + kernel_img_mul_51[14] + 
                kernel_img_mul_51[15] + kernel_img_mul_51[16] + kernel_img_mul_51[17] + 
                kernel_img_mul_51[18] + kernel_img_mul_51[19] + kernel_img_mul_51[20] + 
                kernel_img_mul_51[21] + kernel_img_mul_51[22] + kernel_img_mul_51[23] + 
                kernel_img_mul_51[24];
wire  [39:0]  kernel_img_mul_52[0:24];
assign kernel_img_mul_52[0] = layer0[52][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_52[1] = layer0[52][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_52[2] = layer0[52][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_52[3] = layer0[52][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_52[4] = layer0[52][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_52[5] = layer1[52][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_52[6] = layer1[52][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_52[7] = layer1[52][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_52[8] = layer1[52][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_52[9] = layer1[52][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_52[10] = layer2[52][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_52[11] = layer2[52][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_52[12] = layer2[52][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_52[13] = layer2[52][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_52[14] = layer2[52][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_52[15] = layer3[52][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_52[16] = layer3[52][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_52[17] = layer3[52][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_52[18] = layer3[52][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_52[19] = layer3[52][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_52[20] = layer4[52][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_52[21] = layer4[52][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_52[22] = layer4[52][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_52[23] = layer4[52][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_52[24] = layer4[52][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_52 = kernel_img_mul_52[0] + kernel_img_mul_52[1] + kernel_img_mul_52[2] + 
                kernel_img_mul_52[3] + kernel_img_mul_52[4] + kernel_img_mul_52[5] + 
                kernel_img_mul_52[6] + kernel_img_mul_52[7] + kernel_img_mul_52[8] + 
                kernel_img_mul_52[9] + kernel_img_mul_52[10] + kernel_img_mul_52[11] + 
                kernel_img_mul_52[12] + kernel_img_mul_52[13] + kernel_img_mul_52[14] + 
                kernel_img_mul_52[15] + kernel_img_mul_52[16] + kernel_img_mul_52[17] + 
                kernel_img_mul_52[18] + kernel_img_mul_52[19] + kernel_img_mul_52[20] + 
                kernel_img_mul_52[21] + kernel_img_mul_52[22] + kernel_img_mul_52[23] + 
                kernel_img_mul_52[24];
wire  [39:0]  kernel_img_mul_53[0:24];
assign kernel_img_mul_53[0] = layer0[53][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_53[1] = layer0[53][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_53[2] = layer0[53][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_53[3] = layer0[53][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_53[4] = layer0[53][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_53[5] = layer1[53][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_53[6] = layer1[53][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_53[7] = layer1[53][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_53[8] = layer1[53][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_53[9] = layer1[53][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_53[10] = layer2[53][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_53[11] = layer2[53][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_53[12] = layer2[53][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_53[13] = layer2[53][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_53[14] = layer2[53][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_53[15] = layer3[53][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_53[16] = layer3[53][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_53[17] = layer3[53][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_53[18] = layer3[53][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_53[19] = layer3[53][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_53[20] = layer4[53][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_53[21] = layer4[53][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_53[22] = layer4[53][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_53[23] = layer4[53][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_53[24] = layer4[53][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_53 = kernel_img_mul_53[0] + kernel_img_mul_53[1] + kernel_img_mul_53[2] + 
                kernel_img_mul_53[3] + kernel_img_mul_53[4] + kernel_img_mul_53[5] + 
                kernel_img_mul_53[6] + kernel_img_mul_53[7] + kernel_img_mul_53[8] + 
                kernel_img_mul_53[9] + kernel_img_mul_53[10] + kernel_img_mul_53[11] + 
                kernel_img_mul_53[12] + kernel_img_mul_53[13] + kernel_img_mul_53[14] + 
                kernel_img_mul_53[15] + kernel_img_mul_53[16] + kernel_img_mul_53[17] + 
                kernel_img_mul_53[18] + kernel_img_mul_53[19] + kernel_img_mul_53[20] + 
                kernel_img_mul_53[21] + kernel_img_mul_53[22] + kernel_img_mul_53[23] + 
                kernel_img_mul_53[24];
wire  [39:0]  kernel_img_mul_54[0:24];
assign kernel_img_mul_54[0] = layer0[54][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_54[1] = layer0[54][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_54[2] = layer0[54][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_54[3] = layer0[54][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_54[4] = layer0[54][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_54[5] = layer1[54][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_54[6] = layer1[54][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_54[7] = layer1[54][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_54[8] = layer1[54][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_54[9] = layer1[54][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_54[10] = layer2[54][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_54[11] = layer2[54][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_54[12] = layer2[54][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_54[13] = layer2[54][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_54[14] = layer2[54][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_54[15] = layer3[54][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_54[16] = layer3[54][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_54[17] = layer3[54][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_54[18] = layer3[54][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_54[19] = layer3[54][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_54[20] = layer4[54][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_54[21] = layer4[54][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_54[22] = layer4[54][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_54[23] = layer4[54][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_54[24] = layer4[54][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_54 = kernel_img_mul_54[0] + kernel_img_mul_54[1] + kernel_img_mul_54[2] + 
                kernel_img_mul_54[3] + kernel_img_mul_54[4] + kernel_img_mul_54[5] + 
                kernel_img_mul_54[6] + kernel_img_mul_54[7] + kernel_img_mul_54[8] + 
                kernel_img_mul_54[9] + kernel_img_mul_54[10] + kernel_img_mul_54[11] + 
                kernel_img_mul_54[12] + kernel_img_mul_54[13] + kernel_img_mul_54[14] + 
                kernel_img_mul_54[15] + kernel_img_mul_54[16] + kernel_img_mul_54[17] + 
                kernel_img_mul_54[18] + kernel_img_mul_54[19] + kernel_img_mul_54[20] + 
                kernel_img_mul_54[21] + kernel_img_mul_54[22] + kernel_img_mul_54[23] + 
                kernel_img_mul_54[24];
wire  [39:0]  kernel_img_mul_55[0:24];
assign kernel_img_mul_55[0] = layer0[55][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_55[1] = layer0[55][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_55[2] = layer0[55][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_55[3] = layer0[55][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_55[4] = layer0[55][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_55[5] = layer1[55][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_55[6] = layer1[55][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_55[7] = layer1[55][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_55[8] = layer1[55][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_55[9] = layer1[55][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_55[10] = layer2[55][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_55[11] = layer2[55][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_55[12] = layer2[55][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_55[13] = layer2[55][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_55[14] = layer2[55][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_55[15] = layer3[55][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_55[16] = layer3[55][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_55[17] = layer3[55][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_55[18] = layer3[55][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_55[19] = layer3[55][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_55[20] = layer4[55][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_55[21] = layer4[55][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_55[22] = layer4[55][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_55[23] = layer4[55][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_55[24] = layer4[55][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_55 = kernel_img_mul_55[0] + kernel_img_mul_55[1] + kernel_img_mul_55[2] + 
                kernel_img_mul_55[3] + kernel_img_mul_55[4] + kernel_img_mul_55[5] + 
                kernel_img_mul_55[6] + kernel_img_mul_55[7] + kernel_img_mul_55[8] + 
                kernel_img_mul_55[9] + kernel_img_mul_55[10] + kernel_img_mul_55[11] + 
                kernel_img_mul_55[12] + kernel_img_mul_55[13] + kernel_img_mul_55[14] + 
                kernel_img_mul_55[15] + kernel_img_mul_55[16] + kernel_img_mul_55[17] + 
                kernel_img_mul_55[18] + kernel_img_mul_55[19] + kernel_img_mul_55[20] + 
                kernel_img_mul_55[21] + kernel_img_mul_55[22] + kernel_img_mul_55[23] + 
                kernel_img_mul_55[24];
wire  [39:0]  kernel_img_mul_56[0:24];
assign kernel_img_mul_56[0] = layer0[56][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_56[1] = layer0[56][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_56[2] = layer0[56][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_56[3] = layer0[56][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_56[4] = layer0[56][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_56[5] = layer1[56][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_56[6] = layer1[56][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_56[7] = layer1[56][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_56[8] = layer1[56][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_56[9] = layer1[56][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_56[10] = layer2[56][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_56[11] = layer2[56][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_56[12] = layer2[56][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_56[13] = layer2[56][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_56[14] = layer2[56][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_56[15] = layer3[56][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_56[16] = layer3[56][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_56[17] = layer3[56][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_56[18] = layer3[56][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_56[19] = layer3[56][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_56[20] = layer4[56][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_56[21] = layer4[56][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_56[22] = layer4[56][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_56[23] = layer4[56][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_56[24] = layer4[56][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_56 = kernel_img_mul_56[0] + kernel_img_mul_56[1] + kernel_img_mul_56[2] + 
                kernel_img_mul_56[3] + kernel_img_mul_56[4] + kernel_img_mul_56[5] + 
                kernel_img_mul_56[6] + kernel_img_mul_56[7] + kernel_img_mul_56[8] + 
                kernel_img_mul_56[9] + kernel_img_mul_56[10] + kernel_img_mul_56[11] + 
                kernel_img_mul_56[12] + kernel_img_mul_56[13] + kernel_img_mul_56[14] + 
                kernel_img_mul_56[15] + kernel_img_mul_56[16] + kernel_img_mul_56[17] + 
                kernel_img_mul_56[18] + kernel_img_mul_56[19] + kernel_img_mul_56[20] + 
                kernel_img_mul_56[21] + kernel_img_mul_56[22] + kernel_img_mul_56[23] + 
                kernel_img_mul_56[24];
wire  [39:0]  kernel_img_mul_57[0:24];
assign kernel_img_mul_57[0] = layer0[57][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_57[1] = layer0[57][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_57[2] = layer0[57][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_57[3] = layer0[57][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_57[4] = layer0[57][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_57[5] = layer1[57][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_57[6] = layer1[57][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_57[7] = layer1[57][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_57[8] = layer1[57][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_57[9] = layer1[57][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_57[10] = layer2[57][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_57[11] = layer2[57][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_57[12] = layer2[57][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_57[13] = layer2[57][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_57[14] = layer2[57][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_57[15] = layer3[57][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_57[16] = layer3[57][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_57[17] = layer3[57][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_57[18] = layer3[57][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_57[19] = layer3[57][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_57[20] = layer4[57][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_57[21] = layer4[57][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_57[22] = layer4[57][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_57[23] = layer4[57][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_57[24] = layer4[57][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_57 = kernel_img_mul_57[0] + kernel_img_mul_57[1] + kernel_img_mul_57[2] + 
                kernel_img_mul_57[3] + kernel_img_mul_57[4] + kernel_img_mul_57[5] + 
                kernel_img_mul_57[6] + kernel_img_mul_57[7] + kernel_img_mul_57[8] + 
                kernel_img_mul_57[9] + kernel_img_mul_57[10] + kernel_img_mul_57[11] + 
                kernel_img_mul_57[12] + kernel_img_mul_57[13] + kernel_img_mul_57[14] + 
                kernel_img_mul_57[15] + kernel_img_mul_57[16] + kernel_img_mul_57[17] + 
                kernel_img_mul_57[18] + kernel_img_mul_57[19] + kernel_img_mul_57[20] + 
                kernel_img_mul_57[21] + kernel_img_mul_57[22] + kernel_img_mul_57[23] + 
                kernel_img_mul_57[24];
wire  [39:0]  kernel_img_mul_58[0:24];
assign kernel_img_mul_58[0] = layer0[58][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_58[1] = layer0[58][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_58[2] = layer0[58][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_58[3] = layer0[58][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_58[4] = layer0[58][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_58[5] = layer1[58][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_58[6] = layer1[58][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_58[7] = layer1[58][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_58[8] = layer1[58][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_58[9] = layer1[58][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_58[10] = layer2[58][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_58[11] = layer2[58][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_58[12] = layer2[58][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_58[13] = layer2[58][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_58[14] = layer2[58][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_58[15] = layer3[58][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_58[16] = layer3[58][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_58[17] = layer3[58][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_58[18] = layer3[58][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_58[19] = layer3[58][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_58[20] = layer4[58][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_58[21] = layer4[58][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_58[22] = layer4[58][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_58[23] = layer4[58][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_58[24] = layer4[58][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_58 = kernel_img_mul_58[0] + kernel_img_mul_58[1] + kernel_img_mul_58[2] + 
                kernel_img_mul_58[3] + kernel_img_mul_58[4] + kernel_img_mul_58[5] + 
                kernel_img_mul_58[6] + kernel_img_mul_58[7] + kernel_img_mul_58[8] + 
                kernel_img_mul_58[9] + kernel_img_mul_58[10] + kernel_img_mul_58[11] + 
                kernel_img_mul_58[12] + kernel_img_mul_58[13] + kernel_img_mul_58[14] + 
                kernel_img_mul_58[15] + kernel_img_mul_58[16] + kernel_img_mul_58[17] + 
                kernel_img_mul_58[18] + kernel_img_mul_58[19] + kernel_img_mul_58[20] + 
                kernel_img_mul_58[21] + kernel_img_mul_58[22] + kernel_img_mul_58[23] + 
                kernel_img_mul_58[24];
wire  [39:0]  kernel_img_mul_59[0:24];
assign kernel_img_mul_59[0] = layer0[59][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_59[1] = layer0[59][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_59[2] = layer0[59][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_59[3] = layer0[59][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_59[4] = layer0[59][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_59[5] = layer1[59][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_59[6] = layer1[59][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_59[7] = layer1[59][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_59[8] = layer1[59][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_59[9] = layer1[59][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_59[10] = layer2[59][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_59[11] = layer2[59][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_59[12] = layer2[59][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_59[13] = layer2[59][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_59[14] = layer2[59][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_59[15] = layer3[59][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_59[16] = layer3[59][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_59[17] = layer3[59][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_59[18] = layer3[59][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_59[19] = layer3[59][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_59[20] = layer4[59][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_59[21] = layer4[59][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_59[22] = layer4[59][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_59[23] = layer4[59][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_59[24] = layer4[59][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_59 = kernel_img_mul_59[0] + kernel_img_mul_59[1] + kernel_img_mul_59[2] + 
                kernel_img_mul_59[3] + kernel_img_mul_59[4] + kernel_img_mul_59[5] + 
                kernel_img_mul_59[6] + kernel_img_mul_59[7] + kernel_img_mul_59[8] + 
                kernel_img_mul_59[9] + kernel_img_mul_59[10] + kernel_img_mul_59[11] + 
                kernel_img_mul_59[12] + kernel_img_mul_59[13] + kernel_img_mul_59[14] + 
                kernel_img_mul_59[15] + kernel_img_mul_59[16] + kernel_img_mul_59[17] + 
                kernel_img_mul_59[18] + kernel_img_mul_59[19] + kernel_img_mul_59[20] + 
                kernel_img_mul_59[21] + kernel_img_mul_59[22] + kernel_img_mul_59[23] + 
                kernel_img_mul_59[24];
wire  [39:0]  kernel_img_mul_60[0:24];
assign kernel_img_mul_60[0] = layer0[60][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_60[1] = layer0[60][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_60[2] = layer0[60][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_60[3] = layer0[60][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_60[4] = layer0[60][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_60[5] = layer1[60][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_60[6] = layer1[60][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_60[7] = layer1[60][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_60[8] = layer1[60][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_60[9] = layer1[60][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_60[10] = layer2[60][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_60[11] = layer2[60][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_60[12] = layer2[60][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_60[13] = layer2[60][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_60[14] = layer2[60][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_60[15] = layer3[60][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_60[16] = layer3[60][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_60[17] = layer3[60][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_60[18] = layer3[60][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_60[19] = layer3[60][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_60[20] = layer4[60][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_60[21] = layer4[60][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_60[22] = layer4[60][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_60[23] = layer4[60][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_60[24] = layer4[60][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_60 = kernel_img_mul_60[0] + kernel_img_mul_60[1] + kernel_img_mul_60[2] + 
                kernel_img_mul_60[3] + kernel_img_mul_60[4] + kernel_img_mul_60[5] + 
                kernel_img_mul_60[6] + kernel_img_mul_60[7] + kernel_img_mul_60[8] + 
                kernel_img_mul_60[9] + kernel_img_mul_60[10] + kernel_img_mul_60[11] + 
                kernel_img_mul_60[12] + kernel_img_mul_60[13] + kernel_img_mul_60[14] + 
                kernel_img_mul_60[15] + kernel_img_mul_60[16] + kernel_img_mul_60[17] + 
                kernel_img_mul_60[18] + kernel_img_mul_60[19] + kernel_img_mul_60[20] + 
                kernel_img_mul_60[21] + kernel_img_mul_60[22] + kernel_img_mul_60[23] + 
                kernel_img_mul_60[24];
wire  [39:0]  kernel_img_mul_61[0:24];
assign kernel_img_mul_61[0] = layer0[61][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_61[1] = layer0[61][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_61[2] = layer0[61][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_61[3] = layer0[61][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_61[4] = layer0[61][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_61[5] = layer1[61][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_61[6] = layer1[61][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_61[7] = layer1[61][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_61[8] = layer1[61][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_61[9] = layer1[61][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_61[10] = layer2[61][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_61[11] = layer2[61][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_61[12] = layer2[61][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_61[13] = layer2[61][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_61[14] = layer2[61][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_61[15] = layer3[61][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_61[16] = layer3[61][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_61[17] = layer3[61][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_61[18] = layer3[61][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_61[19] = layer3[61][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_61[20] = layer4[61][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_61[21] = layer4[61][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_61[22] = layer4[61][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_61[23] = layer4[61][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_61[24] = layer4[61][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_61 = kernel_img_mul_61[0] + kernel_img_mul_61[1] + kernel_img_mul_61[2] + 
                kernel_img_mul_61[3] + kernel_img_mul_61[4] + kernel_img_mul_61[5] + 
                kernel_img_mul_61[6] + kernel_img_mul_61[7] + kernel_img_mul_61[8] + 
                kernel_img_mul_61[9] + kernel_img_mul_61[10] + kernel_img_mul_61[11] + 
                kernel_img_mul_61[12] + kernel_img_mul_61[13] + kernel_img_mul_61[14] + 
                kernel_img_mul_61[15] + kernel_img_mul_61[16] + kernel_img_mul_61[17] + 
                kernel_img_mul_61[18] + kernel_img_mul_61[19] + kernel_img_mul_61[20] + 
                kernel_img_mul_61[21] + kernel_img_mul_61[22] + kernel_img_mul_61[23] + 
                kernel_img_mul_61[24];
wire  [39:0]  kernel_img_mul_62[0:24];
assign kernel_img_mul_62[0] = layer0[62][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_62[1] = layer0[62][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_62[2] = layer0[62][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_62[3] = layer0[62][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_62[4] = layer0[62][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_62[5] = layer1[62][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_62[6] = layer1[62][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_62[7] = layer1[62][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_62[8] = layer1[62][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_62[9] = layer1[62][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_62[10] = layer2[62][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_62[11] = layer2[62][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_62[12] = layer2[62][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_62[13] = layer2[62][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_62[14] = layer2[62][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_62[15] = layer3[62][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_62[16] = layer3[62][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_62[17] = layer3[62][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_62[18] = layer3[62][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_62[19] = layer3[62][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_62[20] = layer4[62][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_62[21] = layer4[62][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_62[22] = layer4[62][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_62[23] = layer4[62][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_62[24] = layer4[62][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_62 = kernel_img_mul_62[0] + kernel_img_mul_62[1] + kernel_img_mul_62[2] + 
                kernel_img_mul_62[3] + kernel_img_mul_62[4] + kernel_img_mul_62[5] + 
                kernel_img_mul_62[6] + kernel_img_mul_62[7] + kernel_img_mul_62[8] + 
                kernel_img_mul_62[9] + kernel_img_mul_62[10] + kernel_img_mul_62[11] + 
                kernel_img_mul_62[12] + kernel_img_mul_62[13] + kernel_img_mul_62[14] + 
                kernel_img_mul_62[15] + kernel_img_mul_62[16] + kernel_img_mul_62[17] + 
                kernel_img_mul_62[18] + kernel_img_mul_62[19] + kernel_img_mul_62[20] + 
                kernel_img_mul_62[21] + kernel_img_mul_62[22] + kernel_img_mul_62[23] + 
                kernel_img_mul_62[24];
wire  [39:0]  kernel_img_mul_63[0:24];
assign kernel_img_mul_63[0] = layer0[63][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_63[1] = layer0[63][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_63[2] = layer0[63][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_63[3] = layer0[63][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_63[4] = layer0[63][39:32] *  G_Kernel_5x5[0][159:128];
assign kernel_img_mul_63[5] = layer1[63][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_63[6] = layer1[63][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_63[7] = layer1[63][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_63[8] = layer1[63][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_63[9] = layer1[63][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_63[10] = layer2[63][7:0] *  G_Kernel_5x5[2][31:0];
assign kernel_img_mul_63[11] = layer2[63][15:8] *  G_Kernel_5x5[2][63:32];
assign kernel_img_mul_63[12] = layer2[63][23:16] *  G_Kernel_5x5[2][95:64];
assign kernel_img_mul_63[13] = layer2[63][31:24] *  G_Kernel_5x5[2][127:96];
assign kernel_img_mul_63[14] = layer2[63][39:32] *  G_Kernel_5x5[2][159:128];
assign kernel_img_mul_63[15] = layer3[63][7:0] *  G_Kernel_5x5[1][31:0];
assign kernel_img_mul_63[16] = layer3[63][15:8] *  G_Kernel_5x5[1][63:32];
assign kernel_img_mul_63[17] = layer3[63][23:16] *  G_Kernel_5x5[1][95:64];
assign kernel_img_mul_63[18] = layer3[63][31:24] *  G_Kernel_5x5[1][127:96];
assign kernel_img_mul_63[19] = layer3[63][39:32] *  G_Kernel_5x5[1][159:128];
assign kernel_img_mul_63[20] = layer4[63][7:0] *  G_Kernel_5x5[0][31:0];
assign kernel_img_mul_63[21] = layer4[63][15:8] *  G_Kernel_5x5[0][63:32];
assign kernel_img_mul_63[22] = layer4[63][23:16] *  G_Kernel_5x5[0][95:64];
assign kernel_img_mul_63[23] = layer4[63][31:24] *  G_Kernel_5x5[0][127:96];
assign kernel_img_mul_63[24] = layer4[63][39:32] *  G_Kernel_5x5[0][159:128];
wire  [39:0]  kernel_img_sum_63 = kernel_img_mul_63[0] + kernel_img_mul_63[1] + kernel_img_mul_63[2] + 
                kernel_img_mul_63[3] + kernel_img_mul_63[4] + kernel_img_mul_63[5] + 
                kernel_img_mul_63[6] + kernel_img_mul_63[7] + kernel_img_mul_63[8] + 
                kernel_img_mul_63[9] + kernel_img_mul_63[10] + kernel_img_mul_63[11] + 
                kernel_img_mul_63[12] + kernel_img_mul_63[13] + kernel_img_mul_63[14] + 
                kernel_img_mul_63[15] + kernel_img_mul_63[16] + kernel_img_mul_63[17] + 
                kernel_img_mul_63[18] + kernel_img_mul_63[19] + kernel_img_mul_63[20] + 
                kernel_img_mul_63[21] + kernel_img_mul_63[22] + kernel_img_mul_63[23] + 
                kernel_img_mul_63[24];
always @(posedge clk) begin
  if (!rst_n)
    blur_din[7:0] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[7:0] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[7:0] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[15:8] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[15:8] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[15:8] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[23:16] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[23:16] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[23:16] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[31:24] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[31:24] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[31:24] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[39:32] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[39:32] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[39:32] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[47:40] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[47:40] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[47:40] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[55:48] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[55:48] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[55:48] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[63:56] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[63:56] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[63:56] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[71:64] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[71:64] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[71:64] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[79:72] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[79:72] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[79:72] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[87:80] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[87:80] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[87:80] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[95:88] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[95:88] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[95:88] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[103:96] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[103:96] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[103:96] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[111:104] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[111:104] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[111:104] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[119:112] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[119:112] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[119:112] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[127:120] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[127:120] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[127:120] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[135:128] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[135:128] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[135:128] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[143:136] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[143:136] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[143:136] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[151:144] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[151:144] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[151:144] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[159:152] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[159:152] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[159:152] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[167:160] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[167:160] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[167:160] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[175:168] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[175:168] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[175:168] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[183:176] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[183:176] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[183:176] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[191:184] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[191:184] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[191:184] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[199:192] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[199:192] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[199:192] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[207:200] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[207:200] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[207:200] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[215:208] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[215:208] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[215:208] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[223:216] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[223:216] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[223:216] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[231:224] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[231:224] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[231:224] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[239:232] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[239:232] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[239:232] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[247:240] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[247:240] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[247:240] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[255:248] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[255:248] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[255:248] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[263:256] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[263:256] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[263:256] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[271:264] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[271:264] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[271:264] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[279:272] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[279:272] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[279:272] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[287:280] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[287:280] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[287:280] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[295:288] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[295:288] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[295:288] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[303:296] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[303:296] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[303:296] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[311:304] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[311:304] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[311:304] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[319:312] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[319:312] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[319:312] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[327:320] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[327:320] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[327:320] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[335:328] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[335:328] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[335:328] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[343:336] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[343:336] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[343:336] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[351:344] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[351:344] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[351:344] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[359:352] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[359:352] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[359:352] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[367:360] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[367:360] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[367:360] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[375:368] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[375:368] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[375:368] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[383:376] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[383:376] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[383:376] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[391:384] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[391:384] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[391:384] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[399:392] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[399:392] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[399:392] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[407:400] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[407:400] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[407:400] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[415:408] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[415:408] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[415:408] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[423:416] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[423:416] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[423:416] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[431:424] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[431:424] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[431:424] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[439:432] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[439:432] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[439:432] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[447:440] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[447:440] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[447:440] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[455:448] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[455:448] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[455:448] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[463:456] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[463:456] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[463:456] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[471:464] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[471:464] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[471:464] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[479:472] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[479:472] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[479:472] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[487:480] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[487:480] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[487:480] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[495:488] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[495:488] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[495:488] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[503:496] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[503:496] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[503:496] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[511:504] <= 'd0;
  else if (current_state==ST_GAUSSIAN_0)
    blur_din[511:504] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[511:504] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[519:512] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[519:512] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[519:512] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[527:520] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[527:520] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[527:520] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[535:528] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[535:528] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[535:528] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[543:536] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[543:536] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[543:536] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[551:544] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[551:544] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[551:544] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[559:552] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[559:552] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[559:552] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[567:560] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[567:560] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[567:560] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[575:568] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[575:568] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[575:568] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[583:576] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[583:576] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[583:576] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[591:584] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[591:584] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[591:584] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[599:592] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[599:592] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[599:592] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[607:600] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[607:600] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[607:600] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[615:608] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[615:608] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[615:608] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[623:616] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[623:616] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[623:616] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[631:624] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[631:624] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[631:624] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[639:632] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[639:632] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[639:632] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[647:640] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[647:640] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[647:640] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[655:648] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[655:648] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[655:648] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[663:656] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[663:656] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[663:656] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[671:664] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[671:664] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[671:664] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[679:672] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[679:672] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[679:672] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[687:680] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[687:680] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[687:680] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[695:688] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[695:688] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[695:688] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[703:696] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[703:696] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[703:696] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[711:704] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[711:704] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[711:704] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[719:712] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[719:712] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[719:712] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[727:720] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[727:720] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[727:720] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[735:728] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[735:728] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[735:728] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[743:736] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[743:736] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[743:736] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[751:744] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[751:744] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[751:744] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[759:752] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[759:752] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[759:752] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[767:760] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[767:760] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[767:760] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[775:768] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[775:768] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[775:768] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[783:776] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[783:776] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[783:776] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[791:784] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[791:784] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[791:784] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[799:792] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[799:792] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[799:792] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[807:800] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[807:800] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[807:800] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[815:808] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[815:808] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[815:808] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[823:816] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[823:816] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[823:816] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[831:824] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[831:824] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[831:824] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[839:832] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[839:832] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[839:832] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[847:840] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[847:840] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[847:840] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[855:848] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[855:848] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[855:848] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[863:856] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[863:856] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[863:856] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[871:864] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[871:864] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[871:864] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[879:872] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[879:872] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[879:872] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[887:880] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[887:880] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[887:880] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[895:888] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[895:888] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[895:888] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[903:896] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[903:896] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[903:896] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[911:904] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[911:904] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[911:904] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[919:912] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[919:912] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[919:912] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[927:920] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[927:920] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[927:920] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[935:928] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[935:928] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[935:928] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[943:936] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[943:936] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[943:936] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[951:944] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[951:944] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[951:944] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[959:952] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[959:952] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[959:952] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[967:960] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[967:960] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[967:960] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[975:968] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[975:968] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[975:968] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[983:976] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[983:976] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[983:976] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[991:984] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[991:984] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[991:984] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[999:992] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[999:992] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[999:992] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1007:1000] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[1007:1000] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1007:1000] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1015:1008] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[1015:1008] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1015:1008] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1023:1016] <= 'd0;
  else if (current_state==ST_GAUSSIAN_1)
    blur_din[1023:1016] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1023:1016] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1031:1024] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1031:1024] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1031:1024] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1039:1032] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1039:1032] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1039:1032] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1047:1040] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1047:1040] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1047:1040] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1055:1048] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1055:1048] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1055:1048] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1063:1056] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1063:1056] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1063:1056] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1071:1064] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1071:1064] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1071:1064] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1079:1072] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1079:1072] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1079:1072] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1087:1080] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1087:1080] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1087:1080] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1095:1088] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1095:1088] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1095:1088] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1103:1096] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1103:1096] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1103:1096] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1111:1104] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1111:1104] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1111:1104] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1119:1112] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1119:1112] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1119:1112] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1127:1120] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1127:1120] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1127:1120] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1135:1128] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1135:1128] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1135:1128] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1143:1136] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1143:1136] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1143:1136] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1151:1144] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1151:1144] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1151:1144] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1159:1152] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1159:1152] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1159:1152] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1167:1160] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1167:1160] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1167:1160] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1175:1168] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1175:1168] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1175:1168] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1183:1176] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1183:1176] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1183:1176] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1191:1184] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1191:1184] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1191:1184] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1199:1192] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1199:1192] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1199:1192] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1207:1200] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1207:1200] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1207:1200] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1215:1208] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1215:1208] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1215:1208] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1223:1216] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1223:1216] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1223:1216] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1231:1224] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1231:1224] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1231:1224] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1239:1232] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1239:1232] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1239:1232] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1247:1240] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1247:1240] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1247:1240] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1255:1248] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1255:1248] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1255:1248] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1263:1256] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1263:1256] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1263:1256] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1271:1264] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1271:1264] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1271:1264] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1279:1272] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1279:1272] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1279:1272] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1287:1280] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1287:1280] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1287:1280] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1295:1288] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1295:1288] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1295:1288] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1303:1296] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1303:1296] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1303:1296] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1311:1304] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1311:1304] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1311:1304] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1319:1312] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1319:1312] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1319:1312] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1327:1320] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1327:1320] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1327:1320] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1335:1328] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1335:1328] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1335:1328] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1343:1336] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1343:1336] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1343:1336] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1351:1344] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1351:1344] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1351:1344] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1359:1352] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1359:1352] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1359:1352] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1367:1360] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1367:1360] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1367:1360] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1375:1368] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1375:1368] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1375:1368] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1383:1376] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1383:1376] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1383:1376] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1391:1384] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1391:1384] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1391:1384] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1399:1392] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1399:1392] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1399:1392] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1407:1400] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1407:1400] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1407:1400] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1415:1408] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1415:1408] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1415:1408] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1423:1416] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1423:1416] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1423:1416] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1431:1424] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1431:1424] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1431:1424] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1439:1432] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1439:1432] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1439:1432] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1447:1440] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1447:1440] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1447:1440] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1455:1448] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1455:1448] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1455:1448] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1463:1456] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1463:1456] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1463:1456] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1471:1464] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1471:1464] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1471:1464] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1479:1472] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1479:1472] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1479:1472] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1487:1480] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1487:1480] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1487:1480] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1495:1488] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1495:1488] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1495:1488] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1503:1496] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1503:1496] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1503:1496] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1511:1504] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1511:1504] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1511:1504] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1519:1512] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1519:1512] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1519:1512] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1527:1520] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1527:1520] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1527:1520] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1535:1528] <= 'd0;
  else if (current_state==ST_GAUSSIAN_2)
    blur_din[1535:1528] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1535:1528] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1543:1536] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1543:1536] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1543:1536] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1551:1544] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1551:1544] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1551:1544] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1559:1552] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1559:1552] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1559:1552] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1567:1560] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1567:1560] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1567:1560] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1575:1568] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1575:1568] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1575:1568] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1583:1576] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1583:1576] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1583:1576] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1591:1584] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1591:1584] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1591:1584] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1599:1592] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1599:1592] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1599:1592] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1607:1600] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1607:1600] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1607:1600] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1615:1608] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1615:1608] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1615:1608] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1623:1616] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1623:1616] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1623:1616] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1631:1624] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1631:1624] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1631:1624] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1639:1632] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1639:1632] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1639:1632] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1647:1640] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1647:1640] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1647:1640] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1655:1648] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1655:1648] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1655:1648] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1663:1656] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1663:1656] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1663:1656] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1671:1664] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1671:1664] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1671:1664] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1679:1672] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1679:1672] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1679:1672] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1687:1680] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1687:1680] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1687:1680] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1695:1688] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1695:1688] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1695:1688] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1703:1696] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1703:1696] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1703:1696] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1711:1704] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1711:1704] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1711:1704] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1719:1712] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1719:1712] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1719:1712] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1727:1720] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1727:1720] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1727:1720] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1735:1728] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1735:1728] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1735:1728] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1743:1736] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1743:1736] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1743:1736] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1751:1744] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1751:1744] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1751:1744] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1759:1752] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1759:1752] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1759:1752] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1767:1760] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1767:1760] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1767:1760] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1775:1768] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1775:1768] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1775:1768] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1783:1776] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1783:1776] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1783:1776] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1791:1784] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1791:1784] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1791:1784] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1799:1792] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1799:1792] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1799:1792] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1807:1800] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1807:1800] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1807:1800] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1815:1808] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1815:1808] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1815:1808] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1823:1816] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1823:1816] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1823:1816] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1831:1824] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1831:1824] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1831:1824] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1839:1832] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1839:1832] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1839:1832] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1847:1840] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1847:1840] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1847:1840] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1855:1848] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1855:1848] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1855:1848] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1863:1856] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1863:1856] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1863:1856] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1871:1864] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1871:1864] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1871:1864] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1879:1872] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1879:1872] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1879:1872] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1887:1880] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1887:1880] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1887:1880] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1895:1888] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1895:1888] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1895:1888] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1903:1896] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1903:1896] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1903:1896] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1911:1904] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1911:1904] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1911:1904] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1919:1912] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1919:1912] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1919:1912] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1927:1920] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1927:1920] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1927:1920] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1935:1928] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1935:1928] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1935:1928] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1943:1936] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1943:1936] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1943:1936] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1951:1944] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1951:1944] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1951:1944] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1959:1952] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1959:1952] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1959:1952] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1967:1960] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1967:1960] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1967:1960] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1975:1968] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1975:1968] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1975:1968] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1983:1976] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1983:1976] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1983:1976] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1991:1984] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1991:1984] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1991:1984] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[1999:1992] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[1999:1992] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[1999:1992] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2007:2000] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[2007:2000] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2007:2000] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2015:2008] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[2015:2008] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2015:2008] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2023:2016] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[2023:2016] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2023:2016] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2031:2024] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[2031:2024] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2031:2024] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2039:2032] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[2039:2032] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2039:2032] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2047:2040] <= 'd0;
  else if (current_state==ST_GAUSSIAN_3)
    blur_din[2047:2040] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2047:2040] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2055:2048] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2055:2048] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2055:2048] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2063:2056] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2063:2056] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2063:2056] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2071:2064] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2071:2064] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2071:2064] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2079:2072] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2079:2072] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2079:2072] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2087:2080] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2087:2080] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2087:2080] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2095:2088] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2095:2088] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2095:2088] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2103:2096] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2103:2096] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2103:2096] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2111:2104] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2111:2104] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2111:2104] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2119:2112] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2119:2112] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2119:2112] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2127:2120] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2127:2120] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2127:2120] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2135:2128] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2135:2128] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2135:2128] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2143:2136] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2143:2136] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2143:2136] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2151:2144] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2151:2144] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2151:2144] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2159:2152] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2159:2152] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2159:2152] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2167:2160] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2167:2160] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2167:2160] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2175:2168] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2175:2168] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2175:2168] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2183:2176] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2183:2176] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2183:2176] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2191:2184] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2191:2184] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2191:2184] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2199:2192] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2199:2192] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2199:2192] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2207:2200] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2207:2200] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2207:2200] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2215:2208] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2215:2208] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2215:2208] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2223:2216] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2223:2216] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2223:2216] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2231:2224] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2231:2224] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2231:2224] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2239:2232] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2239:2232] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2239:2232] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2247:2240] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2247:2240] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2247:2240] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2255:2248] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2255:2248] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2255:2248] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2263:2256] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2263:2256] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2263:2256] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2271:2264] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2271:2264] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2271:2264] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2279:2272] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2279:2272] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2279:2272] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2287:2280] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2287:2280] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2287:2280] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2295:2288] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2295:2288] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2295:2288] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2303:2296] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2303:2296] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2303:2296] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2311:2304] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2311:2304] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2311:2304] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2319:2312] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2319:2312] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2319:2312] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2327:2320] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2327:2320] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2327:2320] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2335:2328] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2335:2328] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2335:2328] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2343:2336] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2343:2336] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2343:2336] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2351:2344] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2351:2344] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2351:2344] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2359:2352] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2359:2352] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2359:2352] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2367:2360] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2367:2360] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2367:2360] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2375:2368] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2375:2368] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2375:2368] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2383:2376] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2383:2376] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2383:2376] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2391:2384] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2391:2384] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2391:2384] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2399:2392] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2399:2392] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2399:2392] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2407:2400] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2407:2400] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2407:2400] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2415:2408] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2415:2408] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2415:2408] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2423:2416] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2423:2416] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2423:2416] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2431:2424] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2431:2424] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2431:2424] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2439:2432] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2439:2432] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2439:2432] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2447:2440] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2447:2440] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2447:2440] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2455:2448] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2455:2448] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2455:2448] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2463:2456] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2463:2456] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2463:2456] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2471:2464] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2471:2464] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2471:2464] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2479:2472] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2479:2472] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2479:2472] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2487:2480] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2487:2480] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2487:2480] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2495:2488] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2495:2488] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2495:2488] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2503:2496] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2503:2496] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2503:2496] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2511:2504] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2511:2504] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2511:2504] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2519:2512] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2519:2512] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2519:2512] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2527:2520] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2527:2520] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2527:2520] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2535:2528] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2535:2528] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2535:2528] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2543:2536] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2543:2536] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2543:2536] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2551:2544] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2551:2544] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2551:2544] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2559:2552] <= 'd0;
  else if (current_state==ST_GAUSSIAN_4)
    blur_din[2559:2552] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2559:2552] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2567:2560] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2567:2560] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2567:2560] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2575:2568] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2575:2568] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2575:2568] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2583:2576] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2583:2576] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2583:2576] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2591:2584] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2591:2584] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2591:2584] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2599:2592] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2599:2592] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2599:2592] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2607:2600] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2607:2600] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2607:2600] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2615:2608] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2615:2608] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2615:2608] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2623:2616] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2623:2616] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2623:2616] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2631:2624] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2631:2624] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2631:2624] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2639:2632] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2639:2632] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2639:2632] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2647:2640] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2647:2640] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2647:2640] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2655:2648] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2655:2648] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2655:2648] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2663:2656] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2663:2656] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2663:2656] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2671:2664] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2671:2664] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2671:2664] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2679:2672] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2679:2672] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2679:2672] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2687:2680] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2687:2680] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2687:2680] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2695:2688] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2695:2688] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2695:2688] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2703:2696] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2703:2696] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2703:2696] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2711:2704] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2711:2704] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2711:2704] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2719:2712] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2719:2712] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2719:2712] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2727:2720] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2727:2720] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2727:2720] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2735:2728] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2735:2728] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2735:2728] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2743:2736] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2743:2736] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2743:2736] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2751:2744] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2751:2744] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2751:2744] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2759:2752] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2759:2752] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2759:2752] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2767:2760] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2767:2760] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2767:2760] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2775:2768] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2775:2768] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2775:2768] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2783:2776] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2783:2776] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2783:2776] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2791:2784] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2791:2784] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2791:2784] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2799:2792] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2799:2792] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2799:2792] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2807:2800] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2807:2800] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2807:2800] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2815:2808] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2815:2808] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2815:2808] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2823:2816] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2823:2816] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2823:2816] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2831:2824] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2831:2824] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2831:2824] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2839:2832] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2839:2832] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2839:2832] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2847:2840] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2847:2840] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2847:2840] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2855:2848] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2855:2848] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2855:2848] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2863:2856] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2863:2856] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2863:2856] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2871:2864] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2871:2864] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2871:2864] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2879:2872] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2879:2872] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2879:2872] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2887:2880] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2887:2880] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2887:2880] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2895:2888] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2895:2888] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2895:2888] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2903:2896] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2903:2896] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2903:2896] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2911:2904] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2911:2904] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2911:2904] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2919:2912] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2919:2912] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2919:2912] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2927:2920] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2927:2920] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2927:2920] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2935:2928] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2935:2928] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2935:2928] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2943:2936] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2943:2936] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2943:2936] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2951:2944] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2951:2944] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2951:2944] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2959:2952] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2959:2952] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2959:2952] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2967:2960] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2967:2960] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2967:2960] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2975:2968] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2975:2968] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2975:2968] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2983:2976] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2983:2976] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2983:2976] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2991:2984] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2991:2984] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2991:2984] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[2999:2992] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[2999:2992] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[2999:2992] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3007:3000] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3007:3000] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3007:3000] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3015:3008] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3015:3008] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3015:3008] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3023:3016] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3023:3016] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3023:3016] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3031:3024] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3031:3024] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3031:3024] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3039:3032] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3039:3032] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3039:3032] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3047:3040] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3047:3040] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3047:3040] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3055:3048] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3055:3048] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3055:3048] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3063:3056] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3063:3056] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3063:3056] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3071:3064] <= 'd0;
  else if (current_state==ST_GAUSSIAN_5)
    blur_din[3071:3064] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3071:3064] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3079:3072] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3079:3072] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3079:3072] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3087:3080] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3087:3080] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3087:3080] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3095:3088] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3095:3088] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3095:3088] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3103:3096] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3103:3096] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3103:3096] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3111:3104] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3111:3104] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3111:3104] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3119:3112] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3119:3112] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3119:3112] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3127:3120] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3127:3120] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3127:3120] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3135:3128] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3135:3128] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3135:3128] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3143:3136] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3143:3136] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3143:3136] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3151:3144] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3151:3144] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3151:3144] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3159:3152] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3159:3152] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3159:3152] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3167:3160] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3167:3160] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3167:3160] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3175:3168] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3175:3168] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3175:3168] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3183:3176] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3183:3176] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3183:3176] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3191:3184] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3191:3184] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3191:3184] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3199:3192] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3199:3192] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3199:3192] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3207:3200] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3207:3200] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3207:3200] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3215:3208] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3215:3208] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3215:3208] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3223:3216] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3223:3216] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3223:3216] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3231:3224] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3231:3224] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3231:3224] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3239:3232] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3239:3232] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3239:3232] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3247:3240] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3247:3240] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3247:3240] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3255:3248] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3255:3248] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3255:3248] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3263:3256] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3263:3256] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3263:3256] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3271:3264] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3271:3264] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3271:3264] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3279:3272] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3279:3272] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3279:3272] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3287:3280] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3287:3280] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3287:3280] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3295:3288] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3295:3288] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3295:3288] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3303:3296] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3303:3296] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3303:3296] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3311:3304] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3311:3304] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3311:3304] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3319:3312] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3319:3312] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3319:3312] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3327:3320] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3327:3320] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3327:3320] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3335:3328] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3335:3328] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3335:3328] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3343:3336] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3343:3336] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3343:3336] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3351:3344] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3351:3344] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3351:3344] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3359:3352] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3359:3352] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3359:3352] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3367:3360] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3367:3360] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3367:3360] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3375:3368] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3375:3368] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3375:3368] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3383:3376] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3383:3376] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3383:3376] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3391:3384] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3391:3384] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3391:3384] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3399:3392] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3399:3392] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3399:3392] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3407:3400] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3407:3400] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3407:3400] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3415:3408] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3415:3408] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3415:3408] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3423:3416] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3423:3416] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3423:3416] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3431:3424] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3431:3424] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3431:3424] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3439:3432] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3439:3432] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3439:3432] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3447:3440] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3447:3440] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3447:3440] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3455:3448] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3455:3448] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3455:3448] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3463:3456] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3463:3456] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3463:3456] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3471:3464] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3471:3464] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3471:3464] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3479:3472] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3479:3472] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3479:3472] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3487:3480] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3487:3480] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3487:3480] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3495:3488] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3495:3488] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3495:3488] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3503:3496] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3503:3496] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3503:3496] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3511:3504] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3511:3504] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3511:3504] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3519:3512] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3519:3512] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3519:3512] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3527:3520] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3527:3520] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3527:3520] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3535:3528] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3535:3528] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3535:3528] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3543:3536] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3543:3536] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3543:3536] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3551:3544] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3551:3544] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3551:3544] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3559:3552] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3559:3552] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3559:3552] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3567:3560] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3567:3560] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3567:3560] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3575:3568] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3575:3568] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3575:3568] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3583:3576] <= 'd0;
  else if (current_state==ST_GAUSSIAN_6)
    blur_din[3583:3576] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3583:3576] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3591:3584] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3591:3584] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3591:3584] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3599:3592] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3599:3592] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3599:3592] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3607:3600] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3607:3600] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3607:3600] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3615:3608] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3615:3608] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3615:3608] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3623:3616] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3623:3616] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3623:3616] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3631:3624] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3631:3624] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3631:3624] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3639:3632] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3639:3632] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3639:3632] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3647:3640] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3647:3640] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3647:3640] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3655:3648] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3655:3648] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3655:3648] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3663:3656] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3663:3656] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3663:3656] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3671:3664] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3671:3664] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3671:3664] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3679:3672] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3679:3672] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3679:3672] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3687:3680] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3687:3680] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3687:3680] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3695:3688] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3695:3688] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3695:3688] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3703:3696] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3703:3696] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3703:3696] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3711:3704] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3711:3704] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3711:3704] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3719:3712] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3719:3712] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3719:3712] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3727:3720] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3727:3720] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3727:3720] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3735:3728] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3735:3728] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3735:3728] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3743:3736] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3743:3736] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3743:3736] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3751:3744] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3751:3744] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3751:3744] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3759:3752] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3759:3752] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3759:3752] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3767:3760] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3767:3760] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3767:3760] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3775:3768] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3775:3768] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3775:3768] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3783:3776] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3783:3776] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3783:3776] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3791:3784] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3791:3784] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3791:3784] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3799:3792] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3799:3792] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3799:3792] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3807:3800] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3807:3800] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3807:3800] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3815:3808] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3815:3808] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3815:3808] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3823:3816] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3823:3816] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3823:3816] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3831:3824] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3831:3824] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3831:3824] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3839:3832] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3839:3832] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3839:3832] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3847:3840] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3847:3840] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3847:3840] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3855:3848] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3855:3848] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3855:3848] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3863:3856] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3863:3856] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3863:3856] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3871:3864] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3871:3864] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3871:3864] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3879:3872] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3879:3872] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3879:3872] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3887:3880] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3887:3880] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3887:3880] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3895:3888] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3895:3888] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3895:3888] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3903:3896] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3903:3896] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3903:3896] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3911:3904] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3911:3904] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3911:3904] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3919:3912] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3919:3912] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3919:3912] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3927:3920] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3927:3920] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3927:3920] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3935:3928] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3935:3928] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3935:3928] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3943:3936] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3943:3936] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3943:3936] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3951:3944] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3951:3944] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3951:3944] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3959:3952] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3959:3952] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3959:3952] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3967:3960] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3967:3960] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3967:3960] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3975:3968] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3975:3968] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3975:3968] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3983:3976] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3983:3976] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3983:3976] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3991:3984] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3991:3984] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3991:3984] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[3999:3992] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[3999:3992] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[3999:3992] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4007:4000] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4007:4000] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4007:4000] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4015:4008] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4015:4008] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4015:4008] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4023:4016] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4023:4016] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4023:4016] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4031:4024] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4031:4024] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4031:4024] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4039:4032] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4039:4032] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4039:4032] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4047:4040] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4047:4040] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4047:4040] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4055:4048] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4055:4048] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4055:4048] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4063:4056] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4063:4056] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4063:4056] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4071:4064] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4071:4064] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4071:4064] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4079:4072] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4079:4072] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4079:4072] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4087:4080] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4087:4080] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4087:4080] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4095:4088] <= 'd0;
  else if (current_state==ST_GAUSSIAN_7)
    blur_din[4095:4088] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4095:4088] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4103:4096] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4103:4096] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4103:4096] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4111:4104] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4111:4104] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4111:4104] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4119:4112] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4119:4112] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4119:4112] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4127:4120] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4127:4120] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4127:4120] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4135:4128] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4135:4128] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4135:4128] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4143:4136] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4143:4136] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4143:4136] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4151:4144] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4151:4144] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4151:4144] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4159:4152] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4159:4152] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4159:4152] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4167:4160] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4167:4160] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4167:4160] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4175:4168] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4175:4168] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4175:4168] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4183:4176] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4183:4176] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4183:4176] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4191:4184] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4191:4184] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4191:4184] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4199:4192] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4199:4192] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4199:4192] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4207:4200] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4207:4200] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4207:4200] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4215:4208] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4215:4208] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4215:4208] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4223:4216] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4223:4216] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4223:4216] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4231:4224] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4231:4224] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4231:4224] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4239:4232] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4239:4232] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4239:4232] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4247:4240] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4247:4240] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4247:4240] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4255:4248] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4255:4248] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4255:4248] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4263:4256] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4263:4256] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4263:4256] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4271:4264] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4271:4264] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4271:4264] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4279:4272] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4279:4272] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4279:4272] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4287:4280] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4287:4280] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4287:4280] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4295:4288] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4295:4288] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4295:4288] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4303:4296] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4303:4296] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4303:4296] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4311:4304] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4311:4304] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4311:4304] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4319:4312] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4319:4312] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4319:4312] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4327:4320] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4327:4320] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4327:4320] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4335:4328] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4335:4328] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4335:4328] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4343:4336] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4343:4336] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4343:4336] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4351:4344] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4351:4344] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4351:4344] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4359:4352] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4359:4352] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4359:4352] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4367:4360] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4367:4360] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4367:4360] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4375:4368] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4375:4368] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4375:4368] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4383:4376] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4383:4376] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4383:4376] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4391:4384] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4391:4384] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4391:4384] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4399:4392] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4399:4392] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4399:4392] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4407:4400] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4407:4400] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4407:4400] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4415:4408] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4415:4408] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4415:4408] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4423:4416] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4423:4416] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4423:4416] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4431:4424] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4431:4424] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4431:4424] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4439:4432] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4439:4432] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4439:4432] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4447:4440] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4447:4440] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4447:4440] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4455:4448] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4455:4448] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4455:4448] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4463:4456] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4463:4456] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4463:4456] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4471:4464] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4471:4464] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4471:4464] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4479:4472] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4479:4472] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4479:4472] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4487:4480] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4487:4480] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4487:4480] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4495:4488] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4495:4488] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4495:4488] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4503:4496] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4503:4496] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4503:4496] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4511:4504] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4511:4504] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4511:4504] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4519:4512] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4519:4512] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4519:4512] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4527:4520] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4527:4520] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4527:4520] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4535:4528] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4535:4528] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4535:4528] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4543:4536] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4543:4536] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4543:4536] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4551:4544] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4551:4544] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4551:4544] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4559:4552] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4559:4552] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4559:4552] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4567:4560] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4567:4560] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4567:4560] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4575:4568] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4575:4568] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4575:4568] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4583:4576] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4583:4576] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4583:4576] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4591:4584] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4591:4584] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4591:4584] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4599:4592] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4599:4592] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4599:4592] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4607:4600] <= 'd0;
  else if (current_state==ST_GAUSSIAN_8)
    blur_din[4607:4600] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4607:4600] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4615:4608] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4615:4608] <= kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4615:4608] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4623:4616] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4623:4616] <= kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4623:4616] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4631:4624] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4631:4624] <= kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4631:4624] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4639:4632] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4639:4632] <= kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4639:4632] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4647:4640] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4647:4640] <= kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4647:4640] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4655:4648] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4655:4648] <= kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4655:4648] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4663:4656] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4663:4656] <= kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4663:4656] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4671:4664] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4671:4664] <= kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4671:4664] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4679:4672] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4679:4672] <= kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4679:4672] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4687:4680] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4687:4680] <= kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4687:4680] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4695:4688] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4695:4688] <= kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4695:4688] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4703:4696] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4703:4696] <= kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4703:4696] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4711:4704] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4711:4704] <= kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4711:4704] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4719:4712] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4719:4712] <= kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4719:4712] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4727:4720] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4727:4720] <= kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4727:4720] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4735:4728] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4735:4728] <= kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4735:4728] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4743:4736] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4743:4736] <= kernel_img_sum_16[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4743:4736] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4751:4744] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4751:4744] <= kernel_img_sum_17[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4751:4744] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4759:4752] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4759:4752] <= kernel_img_sum_18[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4759:4752] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4767:4760] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4767:4760] <= kernel_img_sum_19[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4767:4760] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4775:4768] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4775:4768] <= kernel_img_sum_20[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4775:4768] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4783:4776] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4783:4776] <= kernel_img_sum_21[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4783:4776] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4791:4784] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4791:4784] <= kernel_img_sum_22[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4791:4784] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4799:4792] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4799:4792] <= kernel_img_sum_23[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4799:4792] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4807:4800] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4807:4800] <= kernel_img_sum_24[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4807:4800] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4815:4808] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4815:4808] <= kernel_img_sum_25[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4815:4808] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4823:4816] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4823:4816] <= kernel_img_sum_26[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4823:4816] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4831:4824] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4831:4824] <= kernel_img_sum_27[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4831:4824] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4839:4832] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4839:4832] <= kernel_img_sum_28[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4839:4832] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4847:4840] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4847:4840] <= kernel_img_sum_29[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4847:4840] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4855:4848] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4855:4848] <= kernel_img_sum_30[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4855:4848] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4863:4856] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4863:4856] <= kernel_img_sum_31[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4863:4856] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4871:4864] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4871:4864] <= kernel_img_sum_32[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4871:4864] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4879:4872] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4879:4872] <= kernel_img_sum_33[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4879:4872] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4887:4880] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4887:4880] <= kernel_img_sum_34[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4887:4880] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4895:4888] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4895:4888] <= kernel_img_sum_35[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4895:4888] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4903:4896] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4903:4896] <= kernel_img_sum_36[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4903:4896] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4911:4904] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4911:4904] <= kernel_img_sum_37[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4911:4904] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4919:4912] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4919:4912] <= kernel_img_sum_38[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4919:4912] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4927:4920] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4927:4920] <= kernel_img_sum_39[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4927:4920] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4935:4928] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4935:4928] <= kernel_img_sum_40[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4935:4928] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4943:4936] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4943:4936] <= kernel_img_sum_41[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4943:4936] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4951:4944] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4951:4944] <= kernel_img_sum_42[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4951:4944] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4959:4952] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4959:4952] <= kernel_img_sum_43[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4959:4952] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4967:4960] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4967:4960] <= kernel_img_sum_44[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4967:4960] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4975:4968] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4975:4968] <= kernel_img_sum_45[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4975:4968] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4983:4976] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4983:4976] <= kernel_img_sum_46[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4983:4976] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4991:4984] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4991:4984] <= kernel_img_sum_47[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4991:4984] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[4999:4992] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[4999:4992] <= kernel_img_sum_48[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[4999:4992] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5007:5000] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5007:5000] <= kernel_img_sum_49[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5007:5000] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5015:5008] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5015:5008] <= kernel_img_sum_50[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5015:5008] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5023:5016] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5023:5016] <= kernel_img_sum_51[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5023:5016] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5031:5024] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5031:5024] <= kernel_img_sum_52[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5031:5024] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5039:5032] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5039:5032] <= kernel_img_sum_53[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5039:5032] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5047:5040] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5047:5040] <= kernel_img_sum_54[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5047:5040] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5055:5048] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5055:5048] <= kernel_img_sum_55[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5055:5048] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5063:5056] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5063:5056] <= kernel_img_sum_56[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5063:5056] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5071:5064] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5071:5064] <= kernel_img_sum_57[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5071:5064] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5079:5072] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5079:5072] <= kernel_img_sum_58[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5079:5072] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5087:5080] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5087:5080] <= kernel_img_sum_59[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5087:5080] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5095:5088] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5095:5088] <= kernel_img_sum_60[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5095:5088] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5103:5096] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5103:5096] <= kernel_img_sum_61[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5103:5096] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5111:5104] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5111:5104] <= kernel_img_sum_62[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5111:5104] <= 'd0;
end

always @(posedge clk) begin
  if (!rst_n)
    blur_din[5119:5112] <= 'd0;
  else if (current_state==ST_GAUSSIAN_9)
    blur_din[5119:5112] <= kernel_img_sum_63[39:32];/*Q8.32 -> Q8.0*/
  else if (current_state==ST_IDLE)
    blur_din[5119:5112] <= 'd0;
end


endmodule