module Gaussian_Blur_7x7(
  clk,
  rst_n,
  buffer_data_0,
  buffer_data_1,
  buffer_data_2,
  buffer_data_3,
  buffer_data_4,
  buffer_data_5,
  buffer_data_6,
  current_col,
  blur_out
);

input                 clk;
input                 rst_n;
input         [5:0]   current_col;
input       [175:0]   buffer_data_0;
input       [175:0]   buffer_data_1;
input       [175:0]   buffer_data_2;
input       [175:0]   buffer_data_3;
input       [175:0]   buffer_data_4;
input       [175:0]   buffer_data_5;
input       [175:0]   buffer_data_6;
output reg  [127:0]   blur_out; // wire

reg       [223:0] G_Kernel_7x7  [0:3];
always @(*) begin
  if (!rst_n) begin
    G_Kernel_7x7[0][31:0]    = 32'h03C6EBCB; //18'b000000111100011011;//'d014754;
    G_Kernel_7x7[0][63:32]   = 32'h046AA8A8; //18'b000001000110101010;//'d017252;
    G_Kernel_7x7[0][95:64]   = 32'h04D9ED31; //18'b000001001101100111;//'d018950;
    G_Kernel_7x7[0][127:96]  = 32'h050165DE; //18'b000001010000000101;//'d019552;
    G_Kernel_7x7[0][159:128] = 32'h04D9ED31; //18'b000001001101100111;//'d018950;
    G_Kernel_7x7[0][191:160] = 32'h046AA8A8; //18'b000001000110101010;//'d017252;
    G_Kernel_7x7[0][223:192] = 32'h03C6EBCB; //18'b000000111100011011;//'d014754;
    G_Kernel_7x7[1][31:0]    = 32'h046AA8A8; //18'b000001000110101010;//'d017252;
    G_Kernel_7x7[1][63:32]   = 32'h052A1FB1; //18'b000001010010101000;//'d020174;
    G_Kernel_7x7[1][95:64]   = 32'h05AC3BC7; //18'b000001011010110000;//'d022159;
    G_Kernel_7x7[1][127:96]  = 32'h05DA6392; //18'b000001011101101001;//'d022863;
    G_Kernel_7x7[1][159:128] = 32'h05AC3BC7; //18'b000001011010110000;//'d022159;
    G_Kernel_7x7[1][191:160] = 32'h052A1FB1; //18'b000001010010101000;//'d020174;
    G_Kernel_7x7[1][223:192] = 32'h046AA8A8; //18'b000001000110101010;//'d017252;
    G_Kernel_7x7[2][31:0]    = 32'h04D9ED31; //18'b000001001101100111;//'d018950;
    G_Kernel_7x7[2][63:32]   = 32'h05AC3BC7; //18'b000001011010110000;//'d022159;
    G_Kernel_7x7[2][95:64]   = 32'h063B25B2; //18'b000001100011101100;//'d024340;
    G_Kernel_7x7[2][127:96]  = 32'h066DD847; //18'b000001100110110111;//'d025113;
    G_Kernel_7x7[2][159:128] = 32'h063B25B2; //18'b000001100011101100;//'d024340;
    G_Kernel_7x7[2][191:160] = 32'h05AC3BC7; //18'b000001011010110000;//'d022159;
    G_Kernel_7x7[2][223:192] = 32'h04D9ED31; //18'b000001001101100111;//'d018950;
    G_Kernel_7x7[3][31:0]    = 32'h050165DE; //18'b000001010000000101;//'d019552;
    G_Kernel_7x7[3][63:32]   = 32'h05DA6392; //18'b000001011101101001;//'d022863;
    G_Kernel_7x7[3][95:64]   = 32'h066DD847; //18'b000001100110110111;//'d025113;
    G_Kernel_7x7[3][127:96]  = 32'h06A2275A; //18'b000001101010001000;//'d025911;
    G_Kernel_7x7[3][159:128] = 32'h066DD847; //18'b000001100110110111;//'d025113;
    G_Kernel_7x7[3][191:160] = 32'h05DA6392; //18'b000001011101101001;//'d022863;
    G_Kernel_7x7[3][223:192] = 32'h050165DE; //18'b000001010000000101;//'d019552;
  end
end

reg    [55:0]    layer0[0:15]; //wire
reg    [55:0]    layer1[0:15]; //wire
reg    [55:0]    layer2[0:15]; //wire
reg    [55:0]    layer3[0:15]; //wire
reg    [55:0]    layer4[0:15]; //wire
reg    [55:0]    layer5[0:15]; //wire
reg    [55:0]    layer6[0:15]; //wire
always @(*) begin
  case(current_col)
    'd0: begin
        layer0[0][7:0] = 0;
        layer0[0][15:8] = 0;
        layer0[0][23:16] = 0;
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = 0;
        layer1[0][15:8] = 0;
        layer1[0][23:16] = 0;
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = 0;
        layer2[0][15:8] = 0;
        layer2[0][23:16] = 0;
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = 0;
        layer3[0][15:8] = 0;
        layer3[0][23:16] = 0;
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = 0;
        layer4[0][15:8] = 0;
        layer4[0][23:16] = 0;
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = 0;
        layer5[0][15:8] = 0;
        layer5[0][23:16] = 0;
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = 0;
        layer6[0][15:8] = 0;
        layer6[0][23:16] = 0;
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = 0;
        layer0[1][15:8] = 0;
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = 0;
        layer1[1][15:8] = 0;
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = 0;
        layer2[1][15:8] = 0;
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = 0;
        layer3[1][15:8] = 0;
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = 0;
        layer4[1][15:8] = 0;
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = 0;
        layer5[1][15:8] = 0;
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = 0;
        layer6[1][15:8] = 0;
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = 0;
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = 0;
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = 0;
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = 0;
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = 0;
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = 0;
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = 0;
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd1: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd2: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd3: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd4: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd5: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd6: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd7: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd8: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd9: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd10: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd11: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd12: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd13: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd14: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd15: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd16: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd17: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd18: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd19: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd20: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd21: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd22: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd23: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd24: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd25: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd26: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd27: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd28: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd29: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd30: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd31: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd32: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd33: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd34: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd35: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd36: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd37: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd38: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = buffer_data_6[159:152];
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = buffer_data_5[159:152];
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = buffer_data_4[159:152];
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = buffer_data_3[159:152];
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = buffer_data_2[159:152];
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = buffer_data_1[159:152];
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = buffer_data_0[159:152];
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = buffer_data_6[159:152];
        layer0[14][55:48] = buffer_data_6[167:160];
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = buffer_data_5[159:152];
        layer1[14][55:48] = buffer_data_5[167:160];
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = buffer_data_4[159:152];
        layer2[14][55:48] = buffer_data_4[167:160];
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = buffer_data_3[159:152];
        layer3[14][55:48] = buffer_data_3[167:160];
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = buffer_data_2[159:152];
        layer4[14][55:48] = buffer_data_2[167:160];
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = buffer_data_1[159:152];
        layer5[14][55:48] = buffer_data_1[167:160];
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = buffer_data_0[159:152];
        layer6[14][55:48] = buffer_data_0[167:160];
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = buffer_data_6[159:152];
        layer0[15][47:40] = buffer_data_6[167:160];
        layer0[15][55:48] = buffer_data_6[175:168];
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = buffer_data_5[159:152];
        layer1[15][47:40] = buffer_data_5[167:160];
        layer1[15][55:48] = buffer_data_5[175:168];
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = buffer_data_4[159:152];
        layer2[15][47:40] = buffer_data_4[167:160];
        layer2[15][55:48] = buffer_data_4[175:168];
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = buffer_data_3[159:152];
        layer3[15][47:40] = buffer_data_3[167:160];
        layer3[15][55:48] = buffer_data_3[175:168];
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = buffer_data_2[159:152];
        layer4[15][47:40] = buffer_data_2[167:160];
        layer4[15][55:48] = buffer_data_2[175:168];
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = buffer_data_1[159:152];
        layer5[15][47:40] = buffer_data_1[167:160];
        layer5[15][55:48] = buffer_data_1[175:168];
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = buffer_data_0[159:152];
        layer6[15][47:40] = buffer_data_0[167:160];
        layer6[15][55:48] = buffer_data_0[175:168];
    'd39: begin
        layer0[0][7:0] = buffer_data_6[7:0];
        layer0[0][15:8] = buffer_data_6[15:8];
        layer0[0][23:16] = buffer_data_6[23:16];
        layer0[0][31:24] = buffer_data_6[31:24];
        layer0[0][39:32] = buffer_data_6[39:32];
        layer0[0][47:40] = buffer_data_6[47:40];
        layer0[0][55:48] = buffer_data_6[55:48];
        layer1[0][7:0] = buffer_data_5[7:0];
        layer1[0][15:8] = buffer_data_5[15:8];
        layer1[0][23:16] = buffer_data_5[23:16];
        layer1[0][31:24] = buffer_data_5[31:24];
        layer1[0][39:32] = buffer_data_5[39:32];
        layer1[0][47:40] = buffer_data_5[47:40];
        layer1[0][55:48] = buffer_data_5[55:48];
        layer2[0][7:0] = buffer_data_4[7:0];
        layer2[0][15:8] = buffer_data_4[15:8];
        layer2[0][23:16] = buffer_data_4[23:16];
        layer2[0][31:24] = buffer_data_4[31:24];
        layer2[0][39:32] = buffer_data_4[39:32];
        layer2[0][47:40] = buffer_data_4[47:40];
        layer2[0][55:48] = buffer_data_4[55:48];
        layer3[0][7:0] = buffer_data_3[7:0];
        layer3[0][15:8] = buffer_data_3[15:8];
        layer3[0][23:16] = buffer_data_3[23:16];
        layer3[0][31:24] = buffer_data_3[31:24];
        layer3[0][39:32] = buffer_data_3[39:32];
        layer3[0][47:40] = buffer_data_3[47:40];
        layer3[0][55:48] = buffer_data_3[55:48];
        layer4[0][7:0] = buffer_data_2[7:0];
        layer4[0][15:8] = buffer_data_2[15:8];
        layer4[0][23:16] = buffer_data_2[23:16];
        layer4[0][31:24] = buffer_data_2[31:24];
        layer4[0][39:32] = buffer_data_2[39:32];
        layer4[0][47:40] = buffer_data_2[47:40];
        layer4[0][55:48] = buffer_data_2[55:48];
        layer5[0][7:0] = buffer_data_1[7:0];
        layer5[0][15:8] = buffer_data_1[15:8];
        layer5[0][23:16] = buffer_data_1[23:16];
        layer5[0][31:24] = buffer_data_1[31:24];
        layer5[0][39:32] = buffer_data_1[39:32];
        layer5[0][47:40] = buffer_data_1[47:40];
        layer5[0][55:48] = buffer_data_1[55:48];
        layer6[0][7:0] = buffer_data_0[7:0];
        layer6[0][15:8] = buffer_data_0[15:8];
        layer6[0][23:16] = buffer_data_0[23:16];
        layer6[0][31:24] = buffer_data_0[31:24];
        layer6[0][39:32] = buffer_data_0[39:32];
        layer6[0][47:40] = buffer_data_0[47:40];
        layer6[0][55:48] = buffer_data_0[55:48];
        layer0[1][7:0] = buffer_data_6[15:8];
        layer0[1][15:8] = buffer_data_6[23:16];
        layer0[1][23:16] = buffer_data_6[31:24];
        layer0[1][31:24] = buffer_data_6[39:32];
        layer0[1][39:32] = buffer_data_6[47:40];
        layer0[1][47:40] = buffer_data_6[55:48];
        layer0[1][55:48] = buffer_data_6[63:56];
        layer1[1][7:0] = buffer_data_5[15:8];
        layer1[1][15:8] = buffer_data_5[23:16];
        layer1[1][23:16] = buffer_data_5[31:24];
        layer1[1][31:24] = buffer_data_5[39:32];
        layer1[1][39:32] = buffer_data_5[47:40];
        layer1[1][47:40] = buffer_data_5[55:48];
        layer1[1][55:48] = buffer_data_5[63:56];
        layer2[1][7:0] = buffer_data_4[15:8];
        layer2[1][15:8] = buffer_data_4[23:16];
        layer2[1][23:16] = buffer_data_4[31:24];
        layer2[1][31:24] = buffer_data_4[39:32];
        layer2[1][39:32] = buffer_data_4[47:40];
        layer2[1][47:40] = buffer_data_4[55:48];
        layer2[1][55:48] = buffer_data_4[63:56];
        layer3[1][7:0] = buffer_data_3[15:8];
        layer3[1][15:8] = buffer_data_3[23:16];
        layer3[1][23:16] = buffer_data_3[31:24];
        layer3[1][31:24] = buffer_data_3[39:32];
        layer3[1][39:32] = buffer_data_3[47:40];
        layer3[1][47:40] = buffer_data_3[55:48];
        layer3[1][55:48] = buffer_data_3[63:56];
        layer4[1][7:0] = buffer_data_2[15:8];
        layer4[1][15:8] = buffer_data_2[23:16];
        layer4[1][23:16] = buffer_data_2[31:24];
        layer4[1][31:24] = buffer_data_2[39:32];
        layer4[1][39:32] = buffer_data_2[47:40];
        layer4[1][47:40] = buffer_data_2[55:48];
        layer4[1][55:48] = buffer_data_2[63:56];
        layer5[1][7:0] = buffer_data_1[15:8];
        layer5[1][15:8] = buffer_data_1[23:16];
        layer5[1][23:16] = buffer_data_1[31:24];
        layer5[1][31:24] = buffer_data_1[39:32];
        layer5[1][39:32] = buffer_data_1[47:40];
        layer5[1][47:40] = buffer_data_1[55:48];
        layer5[1][55:48] = buffer_data_1[63:56];
        layer6[1][7:0] = buffer_data_0[15:8];
        layer6[1][15:8] = buffer_data_0[23:16];
        layer6[1][23:16] = buffer_data_0[31:24];
        layer6[1][31:24] = buffer_data_0[39:32];
        layer6[1][39:32] = buffer_data_0[47:40];
        layer6[1][47:40] = buffer_data_0[55:48];
        layer6[1][55:48] = buffer_data_0[63:56];
        layer0[2][7:0] = buffer_data_6[23:16];
        layer0[2][15:8] = buffer_data_6[31:24];
        layer0[2][23:16] = buffer_data_6[39:32];
        layer0[2][31:24] = buffer_data_6[47:40];
        layer0[2][39:32] = buffer_data_6[55:48];
        layer0[2][47:40] = buffer_data_6[63:56];
        layer0[2][55:48] = buffer_data_6[71:64];
        layer1[2][7:0] = buffer_data_5[23:16];
        layer1[2][15:8] = buffer_data_5[31:24];
        layer1[2][23:16] = buffer_data_5[39:32];
        layer1[2][31:24] = buffer_data_5[47:40];
        layer1[2][39:32] = buffer_data_5[55:48];
        layer1[2][47:40] = buffer_data_5[63:56];
        layer1[2][55:48] = buffer_data_5[71:64];
        layer2[2][7:0] = buffer_data_4[23:16];
        layer2[2][15:8] = buffer_data_4[31:24];
        layer2[2][23:16] = buffer_data_4[39:32];
        layer2[2][31:24] = buffer_data_4[47:40];
        layer2[2][39:32] = buffer_data_4[55:48];
        layer2[2][47:40] = buffer_data_4[63:56];
        layer2[2][55:48] = buffer_data_4[71:64];
        layer3[2][7:0] = buffer_data_3[23:16];
        layer3[2][15:8] = buffer_data_3[31:24];
        layer3[2][23:16] = buffer_data_3[39:32];
        layer3[2][31:24] = buffer_data_3[47:40];
        layer3[2][39:32] = buffer_data_3[55:48];
        layer3[2][47:40] = buffer_data_3[63:56];
        layer3[2][55:48] = buffer_data_3[71:64];
        layer4[2][7:0] = buffer_data_2[23:16];
        layer4[2][15:8] = buffer_data_2[31:24];
        layer4[2][23:16] = buffer_data_2[39:32];
        layer4[2][31:24] = buffer_data_2[47:40];
        layer4[2][39:32] = buffer_data_2[55:48];
        layer4[2][47:40] = buffer_data_2[63:56];
        layer4[2][55:48] = buffer_data_2[71:64];
        layer5[2][7:0] = buffer_data_1[23:16];
        layer5[2][15:8] = buffer_data_1[31:24];
        layer5[2][23:16] = buffer_data_1[39:32];
        layer5[2][31:24] = buffer_data_1[47:40];
        layer5[2][39:32] = buffer_data_1[55:48];
        layer5[2][47:40] = buffer_data_1[63:56];
        layer5[2][55:48] = buffer_data_1[71:64];
        layer6[2][7:0] = buffer_data_0[23:16];
        layer6[2][15:8] = buffer_data_0[31:24];
        layer6[2][23:16] = buffer_data_0[39:32];
        layer6[2][31:24] = buffer_data_0[47:40];
        layer6[2][39:32] = buffer_data_0[55:48];
        layer6[2][47:40] = buffer_data_0[63:56];
        layer6[2][55:48] = buffer_data_0[71:64];
        layer0[3][7:0] = buffer_data_6[31:24];
        layer0[3][15:8] = buffer_data_6[39:32];
        layer0[3][23:16] = buffer_data_6[47:40];
        layer0[3][31:24] = buffer_data_6[55:48];
        layer0[3][39:32] = buffer_data_6[63:56];
        layer0[3][47:40] = buffer_data_6[71:64];
        layer0[3][55:48] = buffer_data_6[79:72];
        layer1[3][7:0] = buffer_data_5[31:24];
        layer1[3][15:8] = buffer_data_5[39:32];
        layer1[3][23:16] = buffer_data_5[47:40];
        layer1[3][31:24] = buffer_data_5[55:48];
        layer1[3][39:32] = buffer_data_5[63:56];
        layer1[3][47:40] = buffer_data_5[71:64];
        layer1[3][55:48] = buffer_data_5[79:72];
        layer2[3][7:0] = buffer_data_4[31:24];
        layer2[3][15:8] = buffer_data_4[39:32];
        layer2[3][23:16] = buffer_data_4[47:40];
        layer2[3][31:24] = buffer_data_4[55:48];
        layer2[3][39:32] = buffer_data_4[63:56];
        layer2[3][47:40] = buffer_data_4[71:64];
        layer2[3][55:48] = buffer_data_4[79:72];
        layer3[3][7:0] = buffer_data_3[31:24];
        layer3[3][15:8] = buffer_data_3[39:32];
        layer3[3][23:16] = buffer_data_3[47:40];
        layer3[3][31:24] = buffer_data_3[55:48];
        layer3[3][39:32] = buffer_data_3[63:56];
        layer3[3][47:40] = buffer_data_3[71:64];
        layer3[3][55:48] = buffer_data_3[79:72];
        layer4[3][7:0] = buffer_data_2[31:24];
        layer4[3][15:8] = buffer_data_2[39:32];
        layer4[3][23:16] = buffer_data_2[47:40];
        layer4[3][31:24] = buffer_data_2[55:48];
        layer4[3][39:32] = buffer_data_2[63:56];
        layer4[3][47:40] = buffer_data_2[71:64];
        layer4[3][55:48] = buffer_data_2[79:72];
        layer5[3][7:0] = buffer_data_1[31:24];
        layer5[3][15:8] = buffer_data_1[39:32];
        layer5[3][23:16] = buffer_data_1[47:40];
        layer5[3][31:24] = buffer_data_1[55:48];
        layer5[3][39:32] = buffer_data_1[63:56];
        layer5[3][47:40] = buffer_data_1[71:64];
        layer5[3][55:48] = buffer_data_1[79:72];
        layer6[3][7:0] = buffer_data_0[31:24];
        layer6[3][15:8] = buffer_data_0[39:32];
        layer6[3][23:16] = buffer_data_0[47:40];
        layer6[3][31:24] = buffer_data_0[55:48];
        layer6[3][39:32] = buffer_data_0[63:56];
        layer6[3][47:40] = buffer_data_0[71:64];
        layer6[3][55:48] = buffer_data_0[79:72];
        layer0[4][7:0] = buffer_data_6[39:32];
        layer0[4][15:8] = buffer_data_6[47:40];
        layer0[4][23:16] = buffer_data_6[55:48];
        layer0[4][31:24] = buffer_data_6[63:56];
        layer0[4][39:32] = buffer_data_6[71:64];
        layer0[4][47:40] = buffer_data_6[79:72];
        layer0[4][55:48] = buffer_data_6[87:80];
        layer1[4][7:0] = buffer_data_5[39:32];
        layer1[4][15:8] = buffer_data_5[47:40];
        layer1[4][23:16] = buffer_data_5[55:48];
        layer1[4][31:24] = buffer_data_5[63:56];
        layer1[4][39:32] = buffer_data_5[71:64];
        layer1[4][47:40] = buffer_data_5[79:72];
        layer1[4][55:48] = buffer_data_5[87:80];
        layer2[4][7:0] = buffer_data_4[39:32];
        layer2[4][15:8] = buffer_data_4[47:40];
        layer2[4][23:16] = buffer_data_4[55:48];
        layer2[4][31:24] = buffer_data_4[63:56];
        layer2[4][39:32] = buffer_data_4[71:64];
        layer2[4][47:40] = buffer_data_4[79:72];
        layer2[4][55:48] = buffer_data_4[87:80];
        layer3[4][7:0] = buffer_data_3[39:32];
        layer3[4][15:8] = buffer_data_3[47:40];
        layer3[4][23:16] = buffer_data_3[55:48];
        layer3[4][31:24] = buffer_data_3[63:56];
        layer3[4][39:32] = buffer_data_3[71:64];
        layer3[4][47:40] = buffer_data_3[79:72];
        layer3[4][55:48] = buffer_data_3[87:80];
        layer4[4][7:0] = buffer_data_2[39:32];
        layer4[4][15:8] = buffer_data_2[47:40];
        layer4[4][23:16] = buffer_data_2[55:48];
        layer4[4][31:24] = buffer_data_2[63:56];
        layer4[4][39:32] = buffer_data_2[71:64];
        layer4[4][47:40] = buffer_data_2[79:72];
        layer4[4][55:48] = buffer_data_2[87:80];
        layer5[4][7:0] = buffer_data_1[39:32];
        layer5[4][15:8] = buffer_data_1[47:40];
        layer5[4][23:16] = buffer_data_1[55:48];
        layer5[4][31:24] = buffer_data_1[63:56];
        layer5[4][39:32] = buffer_data_1[71:64];
        layer5[4][47:40] = buffer_data_1[79:72];
        layer5[4][55:48] = buffer_data_1[87:80];
        layer6[4][7:0] = buffer_data_0[39:32];
        layer6[4][15:8] = buffer_data_0[47:40];
        layer6[4][23:16] = buffer_data_0[55:48];
        layer6[4][31:24] = buffer_data_0[63:56];
        layer6[4][39:32] = buffer_data_0[71:64];
        layer6[4][47:40] = buffer_data_0[79:72];
        layer6[4][55:48] = buffer_data_0[87:80];
        layer0[5][7:0] = buffer_data_6[47:40];
        layer0[5][15:8] = buffer_data_6[55:48];
        layer0[5][23:16] = buffer_data_6[63:56];
        layer0[5][31:24] = buffer_data_6[71:64];
        layer0[5][39:32] = buffer_data_6[79:72];
        layer0[5][47:40] = buffer_data_6[87:80];
        layer0[5][55:48] = buffer_data_6[95:88];
        layer1[5][7:0] = buffer_data_5[47:40];
        layer1[5][15:8] = buffer_data_5[55:48];
        layer1[5][23:16] = buffer_data_5[63:56];
        layer1[5][31:24] = buffer_data_5[71:64];
        layer1[5][39:32] = buffer_data_5[79:72];
        layer1[5][47:40] = buffer_data_5[87:80];
        layer1[5][55:48] = buffer_data_5[95:88];
        layer2[5][7:0] = buffer_data_4[47:40];
        layer2[5][15:8] = buffer_data_4[55:48];
        layer2[5][23:16] = buffer_data_4[63:56];
        layer2[5][31:24] = buffer_data_4[71:64];
        layer2[5][39:32] = buffer_data_4[79:72];
        layer2[5][47:40] = buffer_data_4[87:80];
        layer2[5][55:48] = buffer_data_4[95:88];
        layer3[5][7:0] = buffer_data_3[47:40];
        layer3[5][15:8] = buffer_data_3[55:48];
        layer3[5][23:16] = buffer_data_3[63:56];
        layer3[5][31:24] = buffer_data_3[71:64];
        layer3[5][39:32] = buffer_data_3[79:72];
        layer3[5][47:40] = buffer_data_3[87:80];
        layer3[5][55:48] = buffer_data_3[95:88];
        layer4[5][7:0] = buffer_data_2[47:40];
        layer4[5][15:8] = buffer_data_2[55:48];
        layer4[5][23:16] = buffer_data_2[63:56];
        layer4[5][31:24] = buffer_data_2[71:64];
        layer4[5][39:32] = buffer_data_2[79:72];
        layer4[5][47:40] = buffer_data_2[87:80];
        layer4[5][55:48] = buffer_data_2[95:88];
        layer5[5][7:0] = buffer_data_1[47:40];
        layer5[5][15:8] = buffer_data_1[55:48];
        layer5[5][23:16] = buffer_data_1[63:56];
        layer5[5][31:24] = buffer_data_1[71:64];
        layer5[5][39:32] = buffer_data_1[79:72];
        layer5[5][47:40] = buffer_data_1[87:80];
        layer5[5][55:48] = buffer_data_1[95:88];
        layer6[5][7:0] = buffer_data_0[47:40];
        layer6[5][15:8] = buffer_data_0[55:48];
        layer6[5][23:16] = buffer_data_0[63:56];
        layer6[5][31:24] = buffer_data_0[71:64];
        layer6[5][39:32] = buffer_data_0[79:72];
        layer6[5][47:40] = buffer_data_0[87:80];
        layer6[5][55:48] = buffer_data_0[95:88];
        layer0[6][7:0] = buffer_data_6[55:48];
        layer0[6][15:8] = buffer_data_6[63:56];
        layer0[6][23:16] = buffer_data_6[71:64];
        layer0[6][31:24] = buffer_data_6[79:72];
        layer0[6][39:32] = buffer_data_6[87:80];
        layer0[6][47:40] = buffer_data_6[95:88];
        layer0[6][55:48] = buffer_data_6[103:96];
        layer1[6][7:0] = buffer_data_5[55:48];
        layer1[6][15:8] = buffer_data_5[63:56];
        layer1[6][23:16] = buffer_data_5[71:64];
        layer1[6][31:24] = buffer_data_5[79:72];
        layer1[6][39:32] = buffer_data_5[87:80];
        layer1[6][47:40] = buffer_data_5[95:88];
        layer1[6][55:48] = buffer_data_5[103:96];
        layer2[6][7:0] = buffer_data_4[55:48];
        layer2[6][15:8] = buffer_data_4[63:56];
        layer2[6][23:16] = buffer_data_4[71:64];
        layer2[6][31:24] = buffer_data_4[79:72];
        layer2[6][39:32] = buffer_data_4[87:80];
        layer2[6][47:40] = buffer_data_4[95:88];
        layer2[6][55:48] = buffer_data_4[103:96];
        layer3[6][7:0] = buffer_data_3[55:48];
        layer3[6][15:8] = buffer_data_3[63:56];
        layer3[6][23:16] = buffer_data_3[71:64];
        layer3[6][31:24] = buffer_data_3[79:72];
        layer3[6][39:32] = buffer_data_3[87:80];
        layer3[6][47:40] = buffer_data_3[95:88];
        layer3[6][55:48] = buffer_data_3[103:96];
        layer4[6][7:0] = buffer_data_2[55:48];
        layer4[6][15:8] = buffer_data_2[63:56];
        layer4[6][23:16] = buffer_data_2[71:64];
        layer4[6][31:24] = buffer_data_2[79:72];
        layer4[6][39:32] = buffer_data_2[87:80];
        layer4[6][47:40] = buffer_data_2[95:88];
        layer4[6][55:48] = buffer_data_2[103:96];
        layer5[6][7:0] = buffer_data_1[55:48];
        layer5[6][15:8] = buffer_data_1[63:56];
        layer5[6][23:16] = buffer_data_1[71:64];
        layer5[6][31:24] = buffer_data_1[79:72];
        layer5[6][39:32] = buffer_data_1[87:80];
        layer5[6][47:40] = buffer_data_1[95:88];
        layer5[6][55:48] = buffer_data_1[103:96];
        layer6[6][7:0] = buffer_data_0[55:48];
        layer6[6][15:8] = buffer_data_0[63:56];
        layer6[6][23:16] = buffer_data_0[71:64];
        layer6[6][31:24] = buffer_data_0[79:72];
        layer6[6][39:32] = buffer_data_0[87:80];
        layer6[6][47:40] = buffer_data_0[95:88];
        layer6[6][55:48] = buffer_data_0[103:96];
        layer0[7][7:0] = buffer_data_6[63:56];
        layer0[7][15:8] = buffer_data_6[71:64];
        layer0[7][23:16] = buffer_data_6[79:72];
        layer0[7][31:24] = buffer_data_6[87:80];
        layer0[7][39:32] = buffer_data_6[95:88];
        layer0[7][47:40] = buffer_data_6[103:96];
        layer0[7][55:48] = buffer_data_6[111:104];
        layer1[7][7:0] = buffer_data_5[63:56];
        layer1[7][15:8] = buffer_data_5[71:64];
        layer1[7][23:16] = buffer_data_5[79:72];
        layer1[7][31:24] = buffer_data_5[87:80];
        layer1[7][39:32] = buffer_data_5[95:88];
        layer1[7][47:40] = buffer_data_5[103:96];
        layer1[7][55:48] = buffer_data_5[111:104];
        layer2[7][7:0] = buffer_data_4[63:56];
        layer2[7][15:8] = buffer_data_4[71:64];
        layer2[7][23:16] = buffer_data_4[79:72];
        layer2[7][31:24] = buffer_data_4[87:80];
        layer2[7][39:32] = buffer_data_4[95:88];
        layer2[7][47:40] = buffer_data_4[103:96];
        layer2[7][55:48] = buffer_data_4[111:104];
        layer3[7][7:0] = buffer_data_3[63:56];
        layer3[7][15:8] = buffer_data_3[71:64];
        layer3[7][23:16] = buffer_data_3[79:72];
        layer3[7][31:24] = buffer_data_3[87:80];
        layer3[7][39:32] = buffer_data_3[95:88];
        layer3[7][47:40] = buffer_data_3[103:96];
        layer3[7][55:48] = buffer_data_3[111:104];
        layer4[7][7:0] = buffer_data_2[63:56];
        layer4[7][15:8] = buffer_data_2[71:64];
        layer4[7][23:16] = buffer_data_2[79:72];
        layer4[7][31:24] = buffer_data_2[87:80];
        layer4[7][39:32] = buffer_data_2[95:88];
        layer4[7][47:40] = buffer_data_2[103:96];
        layer4[7][55:48] = buffer_data_2[111:104];
        layer5[7][7:0] = buffer_data_1[63:56];
        layer5[7][15:8] = buffer_data_1[71:64];
        layer5[7][23:16] = buffer_data_1[79:72];
        layer5[7][31:24] = buffer_data_1[87:80];
        layer5[7][39:32] = buffer_data_1[95:88];
        layer5[7][47:40] = buffer_data_1[103:96];
        layer5[7][55:48] = buffer_data_1[111:104];
        layer6[7][7:0] = buffer_data_0[63:56];
        layer6[7][15:8] = buffer_data_0[71:64];
        layer6[7][23:16] = buffer_data_0[79:72];
        layer6[7][31:24] = buffer_data_0[87:80];
        layer6[7][39:32] = buffer_data_0[95:88];
        layer6[7][47:40] = buffer_data_0[103:96];
        layer6[7][55:48] = buffer_data_0[111:104];
        layer0[8][7:0] = buffer_data_6[71:64];
        layer0[8][15:8] = buffer_data_6[79:72];
        layer0[8][23:16] = buffer_data_6[87:80];
        layer0[8][31:24] = buffer_data_6[95:88];
        layer0[8][39:32] = buffer_data_6[103:96];
        layer0[8][47:40] = buffer_data_6[111:104];
        layer0[8][55:48] = buffer_data_6[119:112];
        layer1[8][7:0] = buffer_data_5[71:64];
        layer1[8][15:8] = buffer_data_5[79:72];
        layer1[8][23:16] = buffer_data_5[87:80];
        layer1[8][31:24] = buffer_data_5[95:88];
        layer1[8][39:32] = buffer_data_5[103:96];
        layer1[8][47:40] = buffer_data_5[111:104];
        layer1[8][55:48] = buffer_data_5[119:112];
        layer2[8][7:0] = buffer_data_4[71:64];
        layer2[8][15:8] = buffer_data_4[79:72];
        layer2[8][23:16] = buffer_data_4[87:80];
        layer2[8][31:24] = buffer_data_4[95:88];
        layer2[8][39:32] = buffer_data_4[103:96];
        layer2[8][47:40] = buffer_data_4[111:104];
        layer2[8][55:48] = buffer_data_4[119:112];
        layer3[8][7:0] = buffer_data_3[71:64];
        layer3[8][15:8] = buffer_data_3[79:72];
        layer3[8][23:16] = buffer_data_3[87:80];
        layer3[8][31:24] = buffer_data_3[95:88];
        layer3[8][39:32] = buffer_data_3[103:96];
        layer3[8][47:40] = buffer_data_3[111:104];
        layer3[8][55:48] = buffer_data_3[119:112];
        layer4[8][7:0] = buffer_data_2[71:64];
        layer4[8][15:8] = buffer_data_2[79:72];
        layer4[8][23:16] = buffer_data_2[87:80];
        layer4[8][31:24] = buffer_data_2[95:88];
        layer4[8][39:32] = buffer_data_2[103:96];
        layer4[8][47:40] = buffer_data_2[111:104];
        layer4[8][55:48] = buffer_data_2[119:112];
        layer5[8][7:0] = buffer_data_1[71:64];
        layer5[8][15:8] = buffer_data_1[79:72];
        layer5[8][23:16] = buffer_data_1[87:80];
        layer5[8][31:24] = buffer_data_1[95:88];
        layer5[8][39:32] = buffer_data_1[103:96];
        layer5[8][47:40] = buffer_data_1[111:104];
        layer5[8][55:48] = buffer_data_1[119:112];
        layer6[8][7:0] = buffer_data_0[71:64];
        layer6[8][15:8] = buffer_data_0[79:72];
        layer6[8][23:16] = buffer_data_0[87:80];
        layer6[8][31:24] = buffer_data_0[95:88];
        layer6[8][39:32] = buffer_data_0[103:96];
        layer6[8][47:40] = buffer_data_0[111:104];
        layer6[8][55:48] = buffer_data_0[119:112];
        layer0[9][7:0] = buffer_data_6[79:72];
        layer0[9][15:8] = buffer_data_6[87:80];
        layer0[9][23:16] = buffer_data_6[95:88];
        layer0[9][31:24] = buffer_data_6[103:96];
        layer0[9][39:32] = buffer_data_6[111:104];
        layer0[9][47:40] = buffer_data_6[119:112];
        layer0[9][55:48] = buffer_data_6[127:120];
        layer1[9][7:0] = buffer_data_5[79:72];
        layer1[9][15:8] = buffer_data_5[87:80];
        layer1[9][23:16] = buffer_data_5[95:88];
        layer1[9][31:24] = buffer_data_5[103:96];
        layer1[9][39:32] = buffer_data_5[111:104];
        layer1[9][47:40] = buffer_data_5[119:112];
        layer1[9][55:48] = buffer_data_5[127:120];
        layer2[9][7:0] = buffer_data_4[79:72];
        layer2[9][15:8] = buffer_data_4[87:80];
        layer2[9][23:16] = buffer_data_4[95:88];
        layer2[9][31:24] = buffer_data_4[103:96];
        layer2[9][39:32] = buffer_data_4[111:104];
        layer2[9][47:40] = buffer_data_4[119:112];
        layer2[9][55:48] = buffer_data_4[127:120];
        layer3[9][7:0] = buffer_data_3[79:72];
        layer3[9][15:8] = buffer_data_3[87:80];
        layer3[9][23:16] = buffer_data_3[95:88];
        layer3[9][31:24] = buffer_data_3[103:96];
        layer3[9][39:32] = buffer_data_3[111:104];
        layer3[9][47:40] = buffer_data_3[119:112];
        layer3[9][55:48] = buffer_data_3[127:120];
        layer4[9][7:0] = buffer_data_2[79:72];
        layer4[9][15:8] = buffer_data_2[87:80];
        layer4[9][23:16] = buffer_data_2[95:88];
        layer4[9][31:24] = buffer_data_2[103:96];
        layer4[9][39:32] = buffer_data_2[111:104];
        layer4[9][47:40] = buffer_data_2[119:112];
        layer4[9][55:48] = buffer_data_2[127:120];
        layer5[9][7:0] = buffer_data_1[79:72];
        layer5[9][15:8] = buffer_data_1[87:80];
        layer5[9][23:16] = buffer_data_1[95:88];
        layer5[9][31:24] = buffer_data_1[103:96];
        layer5[9][39:32] = buffer_data_1[111:104];
        layer5[9][47:40] = buffer_data_1[119:112];
        layer5[9][55:48] = buffer_data_1[127:120];
        layer6[9][7:0] = buffer_data_0[79:72];
        layer6[9][15:8] = buffer_data_0[87:80];
        layer6[9][23:16] = buffer_data_0[95:88];
        layer6[9][31:24] = buffer_data_0[103:96];
        layer6[9][39:32] = buffer_data_0[111:104];
        layer6[9][47:40] = buffer_data_0[119:112];
        layer6[9][55:48] = buffer_data_0[127:120];
        layer0[10][7:0] = buffer_data_6[87:80];
        layer0[10][15:8] = buffer_data_6[95:88];
        layer0[10][23:16] = buffer_data_6[103:96];
        layer0[10][31:24] = buffer_data_6[111:104];
        layer0[10][39:32] = buffer_data_6[119:112];
        layer0[10][47:40] = buffer_data_6[127:120];
        layer0[10][55:48] = buffer_data_6[135:128];
        layer1[10][7:0] = buffer_data_5[87:80];
        layer1[10][15:8] = buffer_data_5[95:88];
        layer1[10][23:16] = buffer_data_5[103:96];
        layer1[10][31:24] = buffer_data_5[111:104];
        layer1[10][39:32] = buffer_data_5[119:112];
        layer1[10][47:40] = buffer_data_5[127:120];
        layer1[10][55:48] = buffer_data_5[135:128];
        layer2[10][7:0] = buffer_data_4[87:80];
        layer2[10][15:8] = buffer_data_4[95:88];
        layer2[10][23:16] = buffer_data_4[103:96];
        layer2[10][31:24] = buffer_data_4[111:104];
        layer2[10][39:32] = buffer_data_4[119:112];
        layer2[10][47:40] = buffer_data_4[127:120];
        layer2[10][55:48] = buffer_data_4[135:128];
        layer3[10][7:0] = buffer_data_3[87:80];
        layer3[10][15:8] = buffer_data_3[95:88];
        layer3[10][23:16] = buffer_data_3[103:96];
        layer3[10][31:24] = buffer_data_3[111:104];
        layer3[10][39:32] = buffer_data_3[119:112];
        layer3[10][47:40] = buffer_data_3[127:120];
        layer3[10][55:48] = buffer_data_3[135:128];
        layer4[10][7:0] = buffer_data_2[87:80];
        layer4[10][15:8] = buffer_data_2[95:88];
        layer4[10][23:16] = buffer_data_2[103:96];
        layer4[10][31:24] = buffer_data_2[111:104];
        layer4[10][39:32] = buffer_data_2[119:112];
        layer4[10][47:40] = buffer_data_2[127:120];
        layer4[10][55:48] = buffer_data_2[135:128];
        layer5[10][7:0] = buffer_data_1[87:80];
        layer5[10][15:8] = buffer_data_1[95:88];
        layer5[10][23:16] = buffer_data_1[103:96];
        layer5[10][31:24] = buffer_data_1[111:104];
        layer5[10][39:32] = buffer_data_1[119:112];
        layer5[10][47:40] = buffer_data_1[127:120];
        layer5[10][55:48] = buffer_data_1[135:128];
        layer6[10][7:0] = buffer_data_0[87:80];
        layer6[10][15:8] = buffer_data_0[95:88];
        layer6[10][23:16] = buffer_data_0[103:96];
        layer6[10][31:24] = buffer_data_0[111:104];
        layer6[10][39:32] = buffer_data_0[119:112];
        layer6[10][47:40] = buffer_data_0[127:120];
        layer6[10][55:48] = buffer_data_0[135:128];
        layer0[11][7:0] = buffer_data_6[95:88];
        layer0[11][15:8] = buffer_data_6[103:96];
        layer0[11][23:16] = buffer_data_6[111:104];
        layer0[11][31:24] = buffer_data_6[119:112];
        layer0[11][39:32] = buffer_data_6[127:120];
        layer0[11][47:40] = buffer_data_6[135:128];
        layer0[11][55:48] = buffer_data_6[143:136];
        layer1[11][7:0] = buffer_data_5[95:88];
        layer1[11][15:8] = buffer_data_5[103:96];
        layer1[11][23:16] = buffer_data_5[111:104];
        layer1[11][31:24] = buffer_data_5[119:112];
        layer1[11][39:32] = buffer_data_5[127:120];
        layer1[11][47:40] = buffer_data_5[135:128];
        layer1[11][55:48] = buffer_data_5[143:136];
        layer2[11][7:0] = buffer_data_4[95:88];
        layer2[11][15:8] = buffer_data_4[103:96];
        layer2[11][23:16] = buffer_data_4[111:104];
        layer2[11][31:24] = buffer_data_4[119:112];
        layer2[11][39:32] = buffer_data_4[127:120];
        layer2[11][47:40] = buffer_data_4[135:128];
        layer2[11][55:48] = buffer_data_4[143:136];
        layer3[11][7:0] = buffer_data_3[95:88];
        layer3[11][15:8] = buffer_data_3[103:96];
        layer3[11][23:16] = buffer_data_3[111:104];
        layer3[11][31:24] = buffer_data_3[119:112];
        layer3[11][39:32] = buffer_data_3[127:120];
        layer3[11][47:40] = buffer_data_3[135:128];
        layer3[11][55:48] = buffer_data_3[143:136];
        layer4[11][7:0] = buffer_data_2[95:88];
        layer4[11][15:8] = buffer_data_2[103:96];
        layer4[11][23:16] = buffer_data_2[111:104];
        layer4[11][31:24] = buffer_data_2[119:112];
        layer4[11][39:32] = buffer_data_2[127:120];
        layer4[11][47:40] = buffer_data_2[135:128];
        layer4[11][55:48] = buffer_data_2[143:136];
        layer5[11][7:0] = buffer_data_1[95:88];
        layer5[11][15:8] = buffer_data_1[103:96];
        layer5[11][23:16] = buffer_data_1[111:104];
        layer5[11][31:24] = buffer_data_1[119:112];
        layer5[11][39:32] = buffer_data_1[127:120];
        layer5[11][47:40] = buffer_data_1[135:128];
        layer5[11][55:48] = buffer_data_1[143:136];
        layer6[11][7:0] = buffer_data_0[95:88];
        layer6[11][15:8] = buffer_data_0[103:96];
        layer6[11][23:16] = buffer_data_0[111:104];
        layer6[11][31:24] = buffer_data_0[119:112];
        layer6[11][39:32] = buffer_data_0[127:120];
        layer6[11][47:40] = buffer_data_0[135:128];
        layer6[11][55:48] = buffer_data_0[143:136];
        layer0[12][7:0] = buffer_data_6[103:96];
        layer0[12][15:8] = buffer_data_6[111:104];
        layer0[12][23:16] = buffer_data_6[119:112];
        layer0[12][31:24] = buffer_data_6[127:120];
        layer0[12][39:32] = buffer_data_6[135:128];
        layer0[12][47:40] = buffer_data_6[143:136];
        layer0[12][55:48] = buffer_data_6[151:144];
        layer1[12][7:0] = buffer_data_5[103:96];
        layer1[12][15:8] = buffer_data_5[111:104];
        layer1[12][23:16] = buffer_data_5[119:112];
        layer1[12][31:24] = buffer_data_5[127:120];
        layer1[12][39:32] = buffer_data_5[135:128];
        layer1[12][47:40] = buffer_data_5[143:136];
        layer1[12][55:48] = buffer_data_5[151:144];
        layer2[12][7:0] = buffer_data_4[103:96];
        layer2[12][15:8] = buffer_data_4[111:104];
        layer2[12][23:16] = buffer_data_4[119:112];
        layer2[12][31:24] = buffer_data_4[127:120];
        layer2[12][39:32] = buffer_data_4[135:128];
        layer2[12][47:40] = buffer_data_4[143:136];
        layer2[12][55:48] = buffer_data_4[151:144];
        layer3[12][7:0] = buffer_data_3[103:96];
        layer3[12][15:8] = buffer_data_3[111:104];
        layer3[12][23:16] = buffer_data_3[119:112];
        layer3[12][31:24] = buffer_data_3[127:120];
        layer3[12][39:32] = buffer_data_3[135:128];
        layer3[12][47:40] = buffer_data_3[143:136];
        layer3[12][55:48] = buffer_data_3[151:144];
        layer4[12][7:0] = buffer_data_2[103:96];
        layer4[12][15:8] = buffer_data_2[111:104];
        layer4[12][23:16] = buffer_data_2[119:112];
        layer4[12][31:24] = buffer_data_2[127:120];
        layer4[12][39:32] = buffer_data_2[135:128];
        layer4[12][47:40] = buffer_data_2[143:136];
        layer4[12][55:48] = buffer_data_2[151:144];
        layer5[12][7:0] = buffer_data_1[103:96];
        layer5[12][15:8] = buffer_data_1[111:104];
        layer5[12][23:16] = buffer_data_1[119:112];
        layer5[12][31:24] = buffer_data_1[127:120];
        layer5[12][39:32] = buffer_data_1[135:128];
        layer5[12][47:40] = buffer_data_1[143:136];
        layer5[12][55:48] = buffer_data_1[151:144];
        layer6[12][7:0] = buffer_data_0[103:96];
        layer6[12][15:8] = buffer_data_0[111:104];
        layer6[12][23:16] = buffer_data_0[119:112];
        layer6[12][31:24] = buffer_data_0[127:120];
        layer6[12][39:32] = buffer_data_0[135:128];
        layer6[12][47:40] = buffer_data_0[143:136];
        layer6[12][55:48] = buffer_data_0[151:144];
        layer0[13][7:0] = buffer_data_6[111:104];
        layer0[13][15:8] = buffer_data_6[119:112];
        layer0[13][23:16] = buffer_data_6[127:120];
        layer0[13][31:24] = buffer_data_6[135:128];
        layer0[13][39:32] = buffer_data_6[143:136];
        layer0[13][47:40] = buffer_data_6[151:144];
        layer0[13][55:48] = 0;
        layer1[13][7:0] = buffer_data_5[111:104];
        layer1[13][15:8] = buffer_data_5[119:112];
        layer1[13][23:16] = buffer_data_5[127:120];
        layer1[13][31:24] = buffer_data_5[135:128];
        layer1[13][39:32] = buffer_data_5[143:136];
        layer1[13][47:40] = buffer_data_5[151:144];
        layer1[13][55:48] = 0;
        layer2[13][7:0] = buffer_data_4[111:104];
        layer2[13][15:8] = buffer_data_4[119:112];
        layer2[13][23:16] = buffer_data_4[127:120];
        layer2[13][31:24] = buffer_data_4[135:128];
        layer2[13][39:32] = buffer_data_4[143:136];
        layer2[13][47:40] = buffer_data_4[151:144];
        layer2[13][55:48] = 0;
        layer3[13][7:0] = buffer_data_3[111:104];
        layer3[13][15:8] = buffer_data_3[119:112];
        layer3[13][23:16] = buffer_data_3[127:120];
        layer3[13][31:24] = buffer_data_3[135:128];
        layer3[13][39:32] = buffer_data_3[143:136];
        layer3[13][47:40] = buffer_data_3[151:144];
        layer3[13][55:48] = 0;
        layer4[13][7:0] = buffer_data_2[111:104];
        layer4[13][15:8] = buffer_data_2[119:112];
        layer4[13][23:16] = buffer_data_2[127:120];
        layer4[13][31:24] = buffer_data_2[135:128];
        layer4[13][39:32] = buffer_data_2[143:136];
        layer4[13][47:40] = buffer_data_2[151:144];
        layer4[13][55:48] = 0;
        layer5[13][7:0] = buffer_data_1[111:104];
        layer5[13][15:8] = buffer_data_1[119:112];
        layer5[13][23:16] = buffer_data_1[127:120];
        layer5[13][31:24] = buffer_data_1[135:128];
        layer5[13][39:32] = buffer_data_1[143:136];
        layer5[13][47:40] = buffer_data_1[151:144];
        layer5[13][55:48] = 0;
        layer6[13][7:0] = buffer_data_0[111:104];
        layer6[13][15:8] = buffer_data_0[119:112];
        layer6[13][23:16] = buffer_data_0[127:120];
        layer6[13][31:24] = buffer_data_0[135:128];
        layer6[13][39:32] = buffer_data_0[143:136];
        layer6[13][47:40] = buffer_data_0[151:144];
        layer6[13][55:48] = 0;
        layer0[14][7:0] = buffer_data_6[119:112];
        layer0[14][15:8] = buffer_data_6[127:120];
        layer0[14][23:16] = buffer_data_6[135:128];
        layer0[14][31:24] = buffer_data_6[143:136];
        layer0[14][39:32] = buffer_data_6[151:144];
        layer0[14][47:40] = 0;
        layer0[14][55:48] = 0;
        layer1[14][7:0] = buffer_data_5[119:112];
        layer1[14][15:8] = buffer_data_5[127:120];
        layer1[14][23:16] = buffer_data_5[135:128];
        layer1[14][31:24] = buffer_data_5[143:136];
        layer1[14][39:32] = buffer_data_5[151:144];
        layer1[14][47:40] = 0;
        layer1[14][55:48] = 0;
        layer2[14][7:0] = buffer_data_4[119:112];
        layer2[14][15:8] = buffer_data_4[127:120];
        layer2[14][23:16] = buffer_data_4[135:128];
        layer2[14][31:24] = buffer_data_4[143:136];
        layer2[14][39:32] = buffer_data_4[151:144];
        layer2[14][47:40] = 0;
        layer2[14][55:48] = 0;
        layer3[14][7:0] = buffer_data_3[119:112];
        layer3[14][15:8] = buffer_data_3[127:120];
        layer3[14][23:16] = buffer_data_3[135:128];
        layer3[14][31:24] = buffer_data_3[143:136];
        layer3[14][39:32] = buffer_data_3[151:144];
        layer3[14][47:40] = 0;
        layer3[14][55:48] = 0;
        layer4[14][7:0] = buffer_data_2[119:112];
        layer4[14][15:8] = buffer_data_2[127:120];
        layer4[14][23:16] = buffer_data_2[135:128];
        layer4[14][31:24] = buffer_data_2[143:136];
        layer4[14][39:32] = buffer_data_2[151:144];
        layer4[14][47:40] = 0;
        layer4[14][55:48] = 0;
        layer5[14][7:0] = buffer_data_1[119:112];
        layer5[14][15:8] = buffer_data_1[127:120];
        layer5[14][23:16] = buffer_data_1[135:128];
        layer5[14][31:24] = buffer_data_1[143:136];
        layer5[14][39:32] = buffer_data_1[151:144];
        layer5[14][47:40] = 0;
        layer5[14][55:48] = 0;
        layer6[14][7:0] = buffer_data_0[119:112];
        layer6[14][15:8] = buffer_data_0[127:120];
        layer6[14][23:16] = buffer_data_0[135:128];
        layer6[14][31:24] = buffer_data_0[143:136];
        layer6[14][39:32] = buffer_data_0[151:144];
        layer6[14][47:40] = 0;
        layer6[14][55:48] = 0;
        layer0[15][7:0] = buffer_data_6[127:120];
        layer0[15][15:8] = buffer_data_6[135:128];
        layer0[15][23:16] = buffer_data_6[143:136];
        layer0[15][31:24] = buffer_data_6[151:144];
        layer0[15][39:32] = 0;
        layer0[15][47:40] = 0;
        layer0[15][55:48] = 0;
        layer1[15][7:0] = buffer_data_5[127:120];
        layer1[15][15:8] = buffer_data_5[135:128];
        layer1[15][23:16] = buffer_data_5[143:136];
        layer1[15][31:24] = buffer_data_5[151:144];
        layer1[15][39:32] = 0;
        layer1[15][47:40] = 0;
        layer1[15][55:48] = 0;
        layer2[15][7:0] = buffer_data_4[127:120];
        layer2[15][15:8] = buffer_data_4[135:128];
        layer2[15][23:16] = buffer_data_4[143:136];
        layer2[15][31:24] = buffer_data_4[151:144];
        layer2[15][39:32] = 0;
        layer2[15][47:40] = 0;
        layer2[15][55:48] = 0;
        layer3[15][7:0] = buffer_data_3[127:120];
        layer3[15][15:8] = buffer_data_3[135:128];
        layer3[15][23:16] = buffer_data_3[143:136];
        layer3[15][31:24] = buffer_data_3[151:144];
        layer3[15][39:32] = 0;
        layer3[15][47:40] = 0;
        layer3[15][55:48] = 0;
        layer4[15][7:0] = buffer_data_2[127:120];
        layer4[15][15:8] = buffer_data_2[135:128];
        layer4[15][23:16] = buffer_data_2[143:136];
        layer4[15][31:24] = buffer_data_2[151:144];
        layer4[15][39:32] = 0;
        layer4[15][47:40] = 0;
        layer4[15][55:48] = 0;
        layer5[15][7:0] = buffer_data_1[127:120];
        layer5[15][15:8] = buffer_data_1[135:128];
        layer5[15][23:16] = buffer_data_1[143:136];
        layer5[15][31:24] = buffer_data_1[151:144];
        layer5[15][39:32] = 0;
        layer5[15][47:40] = 0;
        layer5[15][55:48] = 0;
        layer6[15][7:0] = buffer_data_0[127:120];
        layer6[15][15:8] = buffer_data_0[135:128];
        layer6[15][23:16] = buffer_data_0[143:136];
        layer6[15][31:24] = buffer_data_0[151:144];
        layer6[15][39:32] = 0;
        layer6[15][47:40] = 0;
        layer6[15][55:48] = 0;
    default: begin
        layer0[0][7:0] = 'd0;
        layer0[0][15:8] = 'd0;
        layer0[0][23:16] = 'd0;
        layer0[0][31:24] = 'd0;
        layer0[0][39:32] = 'd0;
        layer0[0][47:40] = 'd0;
        layer0[0][55:48] = 'd0;
        layer1[0][7:0] = 'd0;
        layer1[0][15:8] = 'd0;
        layer1[0][23:16] = 'd0;
        layer1[0][31:24] = 'd0;
        layer1[0][39:32] = 'd0;
        layer1[0][47:40] = 'd0;
        layer1[0][55:48] = 'd0;
        layer2[0][7:0] = 'd0;
        layer2[0][15:8] = 'd0;
        layer2[0][23:16] = 'd0;
        layer2[0][31:24] = 'd0;
        layer2[0][39:32] = 'd0;
        layer2[0][47:40] = 'd0;
        layer2[0][55:48] = 'd0;
        layer3[0][7:0] = 'd0;
        layer3[0][15:8] = 'd0;
        layer3[0][23:16] = 'd0;
        layer3[0][31:24] = 'd0;
        layer3[0][39:32] = 'd0;
        layer3[0][47:40] = 'd0;
        layer3[0][55:48] = 'd0;
        layer4[0][7:0] = 'd0;
        layer4[0][15:8] = 'd0;
        layer4[0][23:16] = 'd0;
        layer4[0][31:24] = 'd0;
        layer4[0][39:32] = 'd0;
        layer4[0][47:40] = 'd0;
        layer4[0][55:48] = 'd0;
        layer5[0][7:0] = 'd0;
        layer5[0][15:8] = 'd0;
        layer5[0][23:16] = 'd0;
        layer5[0][31:24] = 'd0;
        layer5[0][39:32] = 'd0;
        layer5[0][47:40] = 'd0;
        layer5[0][55:48] = 'd0;
        layer6[0][7:0] = 'd0;
        layer6[0][15:8] = 'd0;
        layer6[0][23:16] = 'd0;
        layer6[0][31:24] = 'd0;
        layer6[0][39:32] = 'd0;
        layer6[0][47:40] = 'd0;
        layer6[0][55:48] = 'd0;
        layer0[1][7:0] = 'd0;
        layer0[1][15:8] = 'd0;
        layer0[1][23:16] = 'd0;
        layer0[1][31:24] = 'd0;
        layer0[1][39:32] = 'd0;
        layer0[1][47:40] = 'd0;
        layer0[1][55:48] = 'd0;
        layer1[1][7:0] = 'd0;
        layer1[1][15:8] = 'd0;
        layer1[1][23:16] = 'd0;
        layer1[1][31:24] = 'd0;
        layer1[1][39:32] = 'd0;
        layer1[1][47:40] = 'd0;
        layer1[1][55:48] = 'd0;
        layer2[1][7:0] = 'd0;
        layer2[1][15:8] = 'd0;
        layer2[1][23:16] = 'd0;
        layer2[1][31:24] = 'd0;
        layer2[1][39:32] = 'd0;
        layer2[1][47:40] = 'd0;
        layer2[1][55:48] = 'd0;
        layer3[1][7:0] = 'd0;
        layer3[1][15:8] = 'd0;
        layer3[1][23:16] = 'd0;
        layer3[1][31:24] = 'd0;
        layer3[1][39:32] = 'd0;
        layer3[1][47:40] = 'd0;
        layer3[1][55:48] = 'd0;
        layer4[1][7:0] = 'd0;
        layer4[1][15:8] = 'd0;
        layer4[1][23:16] = 'd0;
        layer4[1][31:24] = 'd0;
        layer4[1][39:32] = 'd0;
        layer4[1][47:40] = 'd0;
        layer4[1][55:48] = 'd0;
        layer5[1][7:0] = 'd0;
        layer5[1][15:8] = 'd0;
        layer5[1][23:16] = 'd0;
        layer5[1][31:24] = 'd0;
        layer5[1][39:32] = 'd0;
        layer5[1][47:40] = 'd0;
        layer5[1][55:48] = 'd0;
        layer6[1][7:0] = 'd0;
        layer6[1][15:8] = 'd0;
        layer6[1][23:16] = 'd0;
        layer6[1][31:24] = 'd0;
        layer6[1][39:32] = 'd0;
        layer6[1][47:40] = 'd0;
        layer6[1][55:48] = 'd0;
        layer0[2][7:0] = 'd0;
        layer0[2][15:8] = 'd0;
        layer0[2][23:16] = 'd0;
        layer0[2][31:24] = 'd0;
        layer0[2][39:32] = 'd0;
        layer0[2][47:40] = 'd0;
        layer0[2][55:48] = 'd0;
        layer1[2][7:0] = 'd0;
        layer1[2][15:8] = 'd0;
        layer1[2][23:16] = 'd0;
        layer1[2][31:24] = 'd0;
        layer1[2][39:32] = 'd0;
        layer1[2][47:40] = 'd0;
        layer1[2][55:48] = 'd0;
        layer2[2][7:0] = 'd0;
        layer2[2][15:8] = 'd0;
        layer2[2][23:16] = 'd0;
        layer2[2][31:24] = 'd0;
        layer2[2][39:32] = 'd0;
        layer2[2][47:40] = 'd0;
        layer2[2][55:48] = 'd0;
        layer3[2][7:0] = 'd0;
        layer3[2][15:8] = 'd0;
        layer3[2][23:16] = 'd0;
        layer3[2][31:24] = 'd0;
        layer3[2][39:32] = 'd0;
        layer3[2][47:40] = 'd0;
        layer3[2][55:48] = 'd0;
        layer4[2][7:0] = 'd0;
        layer4[2][15:8] = 'd0;
        layer4[2][23:16] = 'd0;
        layer4[2][31:24] = 'd0;
        layer4[2][39:32] = 'd0;
        layer4[2][47:40] = 'd0;
        layer4[2][55:48] = 'd0;
        layer5[2][7:0] = 'd0;
        layer5[2][15:8] = 'd0;
        layer5[2][23:16] = 'd0;
        layer5[2][31:24] = 'd0;
        layer5[2][39:32] = 'd0;
        layer5[2][47:40] = 'd0;
        layer5[2][55:48] = 'd0;
        layer6[2][7:0] = 'd0;
        layer6[2][15:8] = 'd0;
        layer6[2][23:16] = 'd0;
        layer6[2][31:24] = 'd0;
        layer6[2][39:32] = 'd0;
        layer6[2][47:40] = 'd0;
        layer6[2][55:48] = 'd0;
        layer0[3][7:0] = 'd0;
        layer0[3][15:8] = 'd0;
        layer0[3][23:16] = 'd0;
        layer0[3][31:24] = 'd0;
        layer0[3][39:32] = 'd0;
        layer0[3][47:40] = 'd0;
        layer0[3][55:48] = 'd0;
        layer1[3][7:0] = 'd0;
        layer1[3][15:8] = 'd0;
        layer1[3][23:16] = 'd0;
        layer1[3][31:24] = 'd0;
        layer1[3][39:32] = 'd0;
        layer1[3][47:40] = 'd0;
        layer1[3][55:48] = 'd0;
        layer2[3][7:0] = 'd0;
        layer2[3][15:8] = 'd0;
        layer2[3][23:16] = 'd0;
        layer2[3][31:24] = 'd0;
        layer2[3][39:32] = 'd0;
        layer2[3][47:40] = 'd0;
        layer2[3][55:48] = 'd0;
        layer3[3][7:0] = 'd0;
        layer3[3][15:8] = 'd0;
        layer3[3][23:16] = 'd0;
        layer3[3][31:24] = 'd0;
        layer3[3][39:32] = 'd0;
        layer3[3][47:40] = 'd0;
        layer3[3][55:48] = 'd0;
        layer4[3][7:0] = 'd0;
        layer4[3][15:8] = 'd0;
        layer4[3][23:16] = 'd0;
        layer4[3][31:24] = 'd0;
        layer4[3][39:32] = 'd0;
        layer4[3][47:40] = 'd0;
        layer4[3][55:48] = 'd0;
        layer5[3][7:0] = 'd0;
        layer5[3][15:8] = 'd0;
        layer5[3][23:16] = 'd0;
        layer5[3][31:24] = 'd0;
        layer5[3][39:32] = 'd0;
        layer5[3][47:40] = 'd0;
        layer5[3][55:48] = 'd0;
        layer6[3][7:0] = 'd0;
        layer6[3][15:8] = 'd0;
        layer6[3][23:16] = 'd0;
        layer6[3][31:24] = 'd0;
        layer6[3][39:32] = 'd0;
        layer6[3][47:40] = 'd0;
        layer6[3][55:48] = 'd0;
        layer0[4][7:0] = 'd0;
        layer0[4][15:8] = 'd0;
        layer0[4][23:16] = 'd0;
        layer0[4][31:24] = 'd0;
        layer0[4][39:32] = 'd0;
        layer0[4][47:40] = 'd0;
        layer0[4][55:48] = 'd0;
        layer1[4][7:0] = 'd0;
        layer1[4][15:8] = 'd0;
        layer1[4][23:16] = 'd0;
        layer1[4][31:24] = 'd0;
        layer1[4][39:32] = 'd0;
        layer1[4][47:40] = 'd0;
        layer1[4][55:48] = 'd0;
        layer2[4][7:0] = 'd0;
        layer2[4][15:8] = 'd0;
        layer2[4][23:16] = 'd0;
        layer2[4][31:24] = 'd0;
        layer2[4][39:32] = 'd0;
        layer2[4][47:40] = 'd0;
        layer2[4][55:48] = 'd0;
        layer3[4][7:0] = 'd0;
        layer3[4][15:8] = 'd0;
        layer3[4][23:16] = 'd0;
        layer3[4][31:24] = 'd0;
        layer3[4][39:32] = 'd0;
        layer3[4][47:40] = 'd0;
        layer3[4][55:48] = 'd0;
        layer4[4][7:0] = 'd0;
        layer4[4][15:8] = 'd0;
        layer4[4][23:16] = 'd0;
        layer4[4][31:24] = 'd0;
        layer4[4][39:32] = 'd0;
        layer4[4][47:40] = 'd0;
        layer4[4][55:48] = 'd0;
        layer5[4][7:0] = 'd0;
        layer5[4][15:8] = 'd0;
        layer5[4][23:16] = 'd0;
        layer5[4][31:24] = 'd0;
        layer5[4][39:32] = 'd0;
        layer5[4][47:40] = 'd0;
        layer5[4][55:48] = 'd0;
        layer6[4][7:0] = 'd0;
        layer6[4][15:8] = 'd0;
        layer6[4][23:16] = 'd0;
        layer6[4][31:24] = 'd0;
        layer6[4][39:32] = 'd0;
        layer6[4][47:40] = 'd0;
        layer6[4][55:48] = 'd0;
        layer0[5][7:0] = 'd0;
        layer0[5][15:8] = 'd0;
        layer0[5][23:16] = 'd0;
        layer0[5][31:24] = 'd0;
        layer0[5][39:32] = 'd0;
        layer0[5][47:40] = 'd0;
        layer0[5][55:48] = 'd0;
        layer1[5][7:0] = 'd0;
        layer1[5][15:8] = 'd0;
        layer1[5][23:16] = 'd0;
        layer1[5][31:24] = 'd0;
        layer1[5][39:32] = 'd0;
        layer1[5][47:40] = 'd0;
        layer1[5][55:48] = 'd0;
        layer2[5][7:0] = 'd0;
        layer2[5][15:8] = 'd0;
        layer2[5][23:16] = 'd0;
        layer2[5][31:24] = 'd0;
        layer2[5][39:32] = 'd0;
        layer2[5][47:40] = 'd0;
        layer2[5][55:48] = 'd0;
        layer3[5][7:0] = 'd0;
        layer3[5][15:8] = 'd0;
        layer3[5][23:16] = 'd0;
        layer3[5][31:24] = 'd0;
        layer3[5][39:32] = 'd0;
        layer3[5][47:40] = 'd0;
        layer3[5][55:48] = 'd0;
        layer4[5][7:0] = 'd0;
        layer4[5][15:8] = 'd0;
        layer4[5][23:16] = 'd0;
        layer4[5][31:24] = 'd0;
        layer4[5][39:32] = 'd0;
        layer4[5][47:40] = 'd0;
        layer4[5][55:48] = 'd0;
        layer5[5][7:0] = 'd0;
        layer5[5][15:8] = 'd0;
        layer5[5][23:16] = 'd0;
        layer5[5][31:24] = 'd0;
        layer5[5][39:32] = 'd0;
        layer5[5][47:40] = 'd0;
        layer5[5][55:48] = 'd0;
        layer6[5][7:0] = 'd0;
        layer6[5][15:8] = 'd0;
        layer6[5][23:16] = 'd0;
        layer6[5][31:24] = 'd0;
        layer6[5][39:32] = 'd0;
        layer6[5][47:40] = 'd0;
        layer6[5][55:48] = 'd0;
        layer0[6][7:0] = 'd0;
        layer0[6][15:8] = 'd0;
        layer0[6][23:16] = 'd0;
        layer0[6][31:24] = 'd0;
        layer0[6][39:32] = 'd0;
        layer0[6][47:40] = 'd0;
        layer0[6][55:48] = 'd0;
        layer1[6][7:0] = 'd0;
        layer1[6][15:8] = 'd0;
        layer1[6][23:16] = 'd0;
        layer1[6][31:24] = 'd0;
        layer1[6][39:32] = 'd0;
        layer1[6][47:40] = 'd0;
        layer1[6][55:48] = 'd0;
        layer2[6][7:0] = 'd0;
        layer2[6][15:8] = 'd0;
        layer2[6][23:16] = 'd0;
        layer2[6][31:24] = 'd0;
        layer2[6][39:32] = 'd0;
        layer2[6][47:40] = 'd0;
        layer2[6][55:48] = 'd0;
        layer3[6][7:0] = 'd0;
        layer3[6][15:8] = 'd0;
        layer3[6][23:16] = 'd0;
        layer3[6][31:24] = 'd0;
        layer3[6][39:32] = 'd0;
        layer3[6][47:40] = 'd0;
        layer3[6][55:48] = 'd0;
        layer4[6][7:0] = 'd0;
        layer4[6][15:8] = 'd0;
        layer4[6][23:16] = 'd0;
        layer4[6][31:24] = 'd0;
        layer4[6][39:32] = 'd0;
        layer4[6][47:40] = 'd0;
        layer4[6][55:48] = 'd0;
        layer5[6][7:0] = 'd0;
        layer5[6][15:8] = 'd0;
        layer5[6][23:16] = 'd0;
        layer5[6][31:24] = 'd0;
        layer5[6][39:32] = 'd0;
        layer5[6][47:40] = 'd0;
        layer5[6][55:48] = 'd0;
        layer6[6][7:0] = 'd0;
        layer6[6][15:8] = 'd0;
        layer6[6][23:16] = 'd0;
        layer6[6][31:24] = 'd0;
        layer6[6][39:32] = 'd0;
        layer6[6][47:40] = 'd0;
        layer6[6][55:48] = 'd0;
        layer0[7][7:0] = 'd0;
        layer0[7][15:8] = 'd0;
        layer0[7][23:16] = 'd0;
        layer0[7][31:24] = 'd0;
        layer0[7][39:32] = 'd0;
        layer0[7][47:40] = 'd0;
        layer0[7][55:48] = 'd0;
        layer1[7][7:0] = 'd0;
        layer1[7][15:8] = 'd0;
        layer1[7][23:16] = 'd0;
        layer1[7][31:24] = 'd0;
        layer1[7][39:32] = 'd0;
        layer1[7][47:40] = 'd0;
        layer1[7][55:48] = 'd0;
        layer2[7][7:0] = 'd0;
        layer2[7][15:8] = 'd0;
        layer2[7][23:16] = 'd0;
        layer2[7][31:24] = 'd0;
        layer2[7][39:32] = 'd0;
        layer2[7][47:40] = 'd0;
        layer2[7][55:48] = 'd0;
        layer3[7][7:0] = 'd0;
        layer3[7][15:8] = 'd0;
        layer3[7][23:16] = 'd0;
        layer3[7][31:24] = 'd0;
        layer3[7][39:32] = 'd0;
        layer3[7][47:40] = 'd0;
        layer3[7][55:48] = 'd0;
        layer4[7][7:0] = 'd0;
        layer4[7][15:8] = 'd0;
        layer4[7][23:16] = 'd0;
        layer4[7][31:24] = 'd0;
        layer4[7][39:32] = 'd0;
        layer4[7][47:40] = 'd0;
        layer4[7][55:48] = 'd0;
        layer5[7][7:0] = 'd0;
        layer5[7][15:8] = 'd0;
        layer5[7][23:16] = 'd0;
        layer5[7][31:24] = 'd0;
        layer5[7][39:32] = 'd0;
        layer5[7][47:40] = 'd0;
        layer5[7][55:48] = 'd0;
        layer6[7][7:0] = 'd0;
        layer6[7][15:8] = 'd0;
        layer6[7][23:16] = 'd0;
        layer6[7][31:24] = 'd0;
        layer6[7][39:32] = 'd0;
        layer6[7][47:40] = 'd0;
        layer6[7][55:48] = 'd0;
        layer0[8][7:0] = 'd0;
        layer0[8][15:8] = 'd0;
        layer0[8][23:16] = 'd0;
        layer0[8][31:24] = 'd0;
        layer0[8][39:32] = 'd0;
        layer0[8][47:40] = 'd0;
        layer0[8][55:48] = 'd0;
        layer1[8][7:0] = 'd0;
        layer1[8][15:8] = 'd0;
        layer1[8][23:16] = 'd0;
        layer1[8][31:24] = 'd0;
        layer1[8][39:32] = 'd0;
        layer1[8][47:40] = 'd0;
        layer1[8][55:48] = 'd0;
        layer2[8][7:0] = 'd0;
        layer2[8][15:8] = 'd0;
        layer2[8][23:16] = 'd0;
        layer2[8][31:24] = 'd0;
        layer2[8][39:32] = 'd0;
        layer2[8][47:40] = 'd0;
        layer2[8][55:48] = 'd0;
        layer3[8][7:0] = 'd0;
        layer3[8][15:8] = 'd0;
        layer3[8][23:16] = 'd0;
        layer3[8][31:24] = 'd0;
        layer3[8][39:32] = 'd0;
        layer3[8][47:40] = 'd0;
        layer3[8][55:48] = 'd0;
        layer4[8][7:0] = 'd0;
        layer4[8][15:8] = 'd0;
        layer4[8][23:16] = 'd0;
        layer4[8][31:24] = 'd0;
        layer4[8][39:32] = 'd0;
        layer4[8][47:40] = 'd0;
        layer4[8][55:48] = 'd0;
        layer5[8][7:0] = 'd0;
        layer5[8][15:8] = 'd0;
        layer5[8][23:16] = 'd0;
        layer5[8][31:24] = 'd0;
        layer5[8][39:32] = 'd0;
        layer5[8][47:40] = 'd0;
        layer5[8][55:48] = 'd0;
        layer6[8][7:0] = 'd0;
        layer6[8][15:8] = 'd0;
        layer6[8][23:16] = 'd0;
        layer6[8][31:24] = 'd0;
        layer6[8][39:32] = 'd0;
        layer6[8][47:40] = 'd0;
        layer6[8][55:48] = 'd0;
        layer0[9][7:0] = 'd0;
        layer0[9][15:8] = 'd0;
        layer0[9][23:16] = 'd0;
        layer0[9][31:24] = 'd0;
        layer0[9][39:32] = 'd0;
        layer0[9][47:40] = 'd0;
        layer0[9][55:48] = 'd0;
        layer1[9][7:0] = 'd0;
        layer1[9][15:8] = 'd0;
        layer1[9][23:16] = 'd0;
        layer1[9][31:24] = 'd0;
        layer1[9][39:32] = 'd0;
        layer1[9][47:40] = 'd0;
        layer1[9][55:48] = 'd0;
        layer2[9][7:0] = 'd0;
        layer2[9][15:8] = 'd0;
        layer2[9][23:16] = 'd0;
        layer2[9][31:24] = 'd0;
        layer2[9][39:32] = 'd0;
        layer2[9][47:40] = 'd0;
        layer2[9][55:48] = 'd0;
        layer3[9][7:0] = 'd0;
        layer3[9][15:8] = 'd0;
        layer3[9][23:16] = 'd0;
        layer3[9][31:24] = 'd0;
        layer3[9][39:32] = 'd0;
        layer3[9][47:40] = 'd0;
        layer3[9][55:48] = 'd0;
        layer4[9][7:0] = 'd0;
        layer4[9][15:8] = 'd0;
        layer4[9][23:16] = 'd0;
        layer4[9][31:24] = 'd0;
        layer4[9][39:32] = 'd0;
        layer4[9][47:40] = 'd0;
        layer4[9][55:48] = 'd0;
        layer5[9][7:0] = 'd0;
        layer5[9][15:8] = 'd0;
        layer5[9][23:16] = 'd0;
        layer5[9][31:24] = 'd0;
        layer5[9][39:32] = 'd0;
        layer5[9][47:40] = 'd0;
        layer5[9][55:48] = 'd0;
        layer6[9][7:0] = 'd0;
        layer6[9][15:8] = 'd0;
        layer6[9][23:16] = 'd0;
        layer6[9][31:24] = 'd0;
        layer6[9][39:32] = 'd0;
        layer6[9][47:40] = 'd0;
        layer6[9][55:48] = 'd0;
        layer0[10][7:0] = 'd0;
        layer0[10][15:8] = 'd0;
        layer0[10][23:16] = 'd0;
        layer0[10][31:24] = 'd0;
        layer0[10][39:32] = 'd0;
        layer0[10][47:40] = 'd0;
        layer0[10][55:48] = 'd0;
        layer1[10][7:0] = 'd0;
        layer1[10][15:8] = 'd0;
        layer1[10][23:16] = 'd0;
        layer1[10][31:24] = 'd0;
        layer1[10][39:32] = 'd0;
        layer1[10][47:40] = 'd0;
        layer1[10][55:48] = 'd0;
        layer2[10][7:0] = 'd0;
        layer2[10][15:8] = 'd0;
        layer2[10][23:16] = 'd0;
        layer2[10][31:24] = 'd0;
        layer2[10][39:32] = 'd0;
        layer2[10][47:40] = 'd0;
        layer2[10][55:48] = 'd0;
        layer3[10][7:0] = 'd0;
        layer3[10][15:8] = 'd0;
        layer3[10][23:16] = 'd0;
        layer3[10][31:24] = 'd0;
        layer3[10][39:32] = 'd0;
        layer3[10][47:40] = 'd0;
        layer3[10][55:48] = 'd0;
        layer4[10][7:0] = 'd0;
        layer4[10][15:8] = 'd0;
        layer4[10][23:16] = 'd0;
        layer4[10][31:24] = 'd0;
        layer4[10][39:32] = 'd0;
        layer4[10][47:40] = 'd0;
        layer4[10][55:48] = 'd0;
        layer5[10][7:0] = 'd0;
        layer5[10][15:8] = 'd0;
        layer5[10][23:16] = 'd0;
        layer5[10][31:24] = 'd0;
        layer5[10][39:32] = 'd0;
        layer5[10][47:40] = 'd0;
        layer5[10][55:48] = 'd0;
        layer6[10][7:0] = 'd0;
        layer6[10][15:8] = 'd0;
        layer6[10][23:16] = 'd0;
        layer6[10][31:24] = 'd0;
        layer6[10][39:32] = 'd0;
        layer6[10][47:40] = 'd0;
        layer6[10][55:48] = 'd0;
        layer0[11][7:0] = 'd0;
        layer0[11][15:8] = 'd0;
        layer0[11][23:16] = 'd0;
        layer0[11][31:24] = 'd0;
        layer0[11][39:32] = 'd0;
        layer0[11][47:40] = 'd0;
        layer0[11][55:48] = 'd0;
        layer1[11][7:0] = 'd0;
        layer1[11][15:8] = 'd0;
        layer1[11][23:16] = 'd0;
        layer1[11][31:24] = 'd0;
        layer1[11][39:32] = 'd0;
        layer1[11][47:40] = 'd0;
        layer1[11][55:48] = 'd0;
        layer2[11][7:0] = 'd0;
        layer2[11][15:8] = 'd0;
        layer2[11][23:16] = 'd0;
        layer2[11][31:24] = 'd0;
        layer2[11][39:32] = 'd0;
        layer2[11][47:40] = 'd0;
        layer2[11][55:48] = 'd0;
        layer3[11][7:0] = 'd0;
        layer3[11][15:8] = 'd0;
        layer3[11][23:16] = 'd0;
        layer3[11][31:24] = 'd0;
        layer3[11][39:32] = 'd0;
        layer3[11][47:40] = 'd0;
        layer3[11][55:48] = 'd0;
        layer4[11][7:0] = 'd0;
        layer4[11][15:8] = 'd0;
        layer4[11][23:16] = 'd0;
        layer4[11][31:24] = 'd0;
        layer4[11][39:32] = 'd0;
        layer4[11][47:40] = 'd0;
        layer4[11][55:48] = 'd0;
        layer5[11][7:0] = 'd0;
        layer5[11][15:8] = 'd0;
        layer5[11][23:16] = 'd0;
        layer5[11][31:24] = 'd0;
        layer5[11][39:32] = 'd0;
        layer5[11][47:40] = 'd0;
        layer5[11][55:48] = 'd0;
        layer6[11][7:0] = 'd0;
        layer6[11][15:8] = 'd0;
        layer6[11][23:16] = 'd0;
        layer6[11][31:24] = 'd0;
        layer6[11][39:32] = 'd0;
        layer6[11][47:40] = 'd0;
        layer6[11][55:48] = 'd0;
        layer0[12][7:0] = 'd0;
        layer0[12][15:8] = 'd0;
        layer0[12][23:16] = 'd0;
        layer0[12][31:24] = 'd0;
        layer0[12][39:32] = 'd0;
        layer0[12][47:40] = 'd0;
        layer0[12][55:48] = 'd0;
        layer1[12][7:0] = 'd0;
        layer1[12][15:8] = 'd0;
        layer1[12][23:16] = 'd0;
        layer1[12][31:24] = 'd0;
        layer1[12][39:32] = 'd0;
        layer1[12][47:40] = 'd0;
        layer1[12][55:48] = 'd0;
        layer2[12][7:0] = 'd0;
        layer2[12][15:8] = 'd0;
        layer2[12][23:16] = 'd0;
        layer2[12][31:24] = 'd0;
        layer2[12][39:32] = 'd0;
        layer2[12][47:40] = 'd0;
        layer2[12][55:48] = 'd0;
        layer3[12][7:0] = 'd0;
        layer3[12][15:8] = 'd0;
        layer3[12][23:16] = 'd0;
        layer3[12][31:24] = 'd0;
        layer3[12][39:32] = 'd0;
        layer3[12][47:40] = 'd0;
        layer3[12][55:48] = 'd0;
        layer4[12][7:0] = 'd0;
        layer4[12][15:8] = 'd0;
        layer4[12][23:16] = 'd0;
        layer4[12][31:24] = 'd0;
        layer4[12][39:32] = 'd0;
        layer4[12][47:40] = 'd0;
        layer4[12][55:48] = 'd0;
        layer5[12][7:0] = 'd0;
        layer5[12][15:8] = 'd0;
        layer5[12][23:16] = 'd0;
        layer5[12][31:24] = 'd0;
        layer5[12][39:32] = 'd0;
        layer5[12][47:40] = 'd0;
        layer5[12][55:48] = 'd0;
        layer6[12][7:0] = 'd0;
        layer6[12][15:8] = 'd0;
        layer6[12][23:16] = 'd0;
        layer6[12][31:24] = 'd0;
        layer6[12][39:32] = 'd0;
        layer6[12][47:40] = 'd0;
        layer6[12][55:48] = 'd0;
        layer0[13][7:0] = 'd0;
        layer0[13][15:8] = 'd0;
        layer0[13][23:16] = 'd0;
        layer0[13][31:24] = 'd0;
        layer0[13][39:32] = 'd0;
        layer0[13][47:40] = 'd0;
        layer0[13][55:48] = 'd0;
        layer1[13][7:0] = 'd0;
        layer1[13][15:8] = 'd0;
        layer1[13][23:16] = 'd0;
        layer1[13][31:24] = 'd0;
        layer1[13][39:32] = 'd0;
        layer1[13][47:40] = 'd0;
        layer1[13][55:48] = 'd0;
        layer2[13][7:0] = 'd0;
        layer2[13][15:8] = 'd0;
        layer2[13][23:16] = 'd0;
        layer2[13][31:24] = 'd0;
        layer2[13][39:32] = 'd0;
        layer2[13][47:40] = 'd0;
        layer2[13][55:48] = 'd0;
        layer3[13][7:0] = 'd0;
        layer3[13][15:8] = 'd0;
        layer3[13][23:16] = 'd0;
        layer3[13][31:24] = 'd0;
        layer3[13][39:32] = 'd0;
        layer3[13][47:40] = 'd0;
        layer3[13][55:48] = 'd0;
        layer4[13][7:0] = 'd0;
        layer4[13][15:8] = 'd0;
        layer4[13][23:16] = 'd0;
        layer4[13][31:24] = 'd0;
        layer4[13][39:32] = 'd0;
        layer4[13][47:40] = 'd0;
        layer4[13][55:48] = 'd0;
        layer5[13][7:0] = 'd0;
        layer5[13][15:8] = 'd0;
        layer5[13][23:16] = 'd0;
        layer5[13][31:24] = 'd0;
        layer5[13][39:32] = 'd0;
        layer5[13][47:40] = 'd0;
        layer5[13][55:48] = 'd0;
        layer6[13][7:0] = 'd0;
        layer6[13][15:8] = 'd0;
        layer6[13][23:16] = 'd0;
        layer6[13][31:24] = 'd0;
        layer6[13][39:32] = 'd0;
        layer6[13][47:40] = 'd0;
        layer6[13][55:48] = 'd0;
        layer0[14][7:0] = 'd0;
        layer0[14][15:8] = 'd0;
        layer0[14][23:16] = 'd0;
        layer0[14][31:24] = 'd0;
        layer0[14][39:32] = 'd0;
        layer0[14][47:40] = 'd0;
        layer0[14][55:48] = 'd0;
        layer1[14][7:0] = 'd0;
        layer1[14][15:8] = 'd0;
        layer1[14][23:16] = 'd0;
        layer1[14][31:24] = 'd0;
        layer1[14][39:32] = 'd0;
        layer1[14][47:40] = 'd0;
        layer1[14][55:48] = 'd0;
        layer2[14][7:0] = 'd0;
        layer2[14][15:8] = 'd0;
        layer2[14][23:16] = 'd0;
        layer2[14][31:24] = 'd0;
        layer2[14][39:32] = 'd0;
        layer2[14][47:40] = 'd0;
        layer2[14][55:48] = 'd0;
        layer3[14][7:0] = 'd0;
        layer3[14][15:8] = 'd0;
        layer3[14][23:16] = 'd0;
        layer3[14][31:24] = 'd0;
        layer3[14][39:32] = 'd0;
        layer3[14][47:40] = 'd0;
        layer3[14][55:48] = 'd0;
        layer4[14][7:0] = 'd0;
        layer4[14][15:8] = 'd0;
        layer4[14][23:16] = 'd0;
        layer4[14][31:24] = 'd0;
        layer4[14][39:32] = 'd0;
        layer4[14][47:40] = 'd0;
        layer4[14][55:48] = 'd0;
        layer5[14][7:0] = 'd0;
        layer5[14][15:8] = 'd0;
        layer5[14][23:16] = 'd0;
        layer5[14][31:24] = 'd0;
        layer5[14][39:32] = 'd0;
        layer5[14][47:40] = 'd0;
        layer5[14][55:48] = 'd0;
        layer6[14][7:0] = 'd0;
        layer6[14][15:8] = 'd0;
        layer6[14][23:16] = 'd0;
        layer6[14][31:24] = 'd0;
        layer6[14][39:32] = 'd0;
        layer6[14][47:40] = 'd0;
        layer6[14][55:48] = 'd0;
        layer0[15][7:0] = 'd0;
        layer0[15][15:8] = 'd0;
        layer0[15][23:16] = 'd0;
        layer0[15][31:24] = 'd0;
        layer0[15][39:32] = 'd0;
        layer0[15][47:40] = 'd0;
        layer0[15][55:48] = 'd0;
        layer1[15][7:0] = 'd0;
        layer1[15][15:8] = 'd0;
        layer1[15][23:16] = 'd0;
        layer1[15][31:24] = 'd0;
        layer1[15][39:32] = 'd0;
        layer1[15][47:40] = 'd0;
        layer1[15][55:48] = 'd0;
        layer2[15][7:0] = 'd0;
        layer2[15][15:8] = 'd0;
        layer2[15][23:16] = 'd0;
        layer2[15][31:24] = 'd0;
        layer2[15][39:32] = 'd0;
        layer2[15][47:40] = 'd0;
        layer2[15][55:48] = 'd0;
        layer3[15][7:0] = 'd0;
        layer3[15][15:8] = 'd0;
        layer3[15][23:16] = 'd0;
        layer3[15][31:24] = 'd0;
        layer3[15][39:32] = 'd0;
        layer3[15][47:40] = 'd0;
        layer3[15][55:48] = 'd0;
        layer4[15][7:0] = 'd0;
        layer4[15][15:8] = 'd0;
        layer4[15][23:16] = 'd0;
        layer4[15][31:24] = 'd0;
        layer4[15][39:32] = 'd0;
        layer4[15][47:40] = 'd0;
        layer4[15][55:48] = 'd0;
        layer5[15][7:0] = 'd0;
        layer5[15][15:8] = 'd0;
        layer5[15][23:16] = 'd0;
        layer5[15][31:24] = 'd0;
        layer5[15][39:32] = 'd0;
        layer5[15][47:40] = 'd0;
        layer5[15][55:48] = 'd0;
        layer6[15][7:0] = 'd0;
        layer6[15][15:8] = 'd0;
        layer6[15][23:16] = 'd0;
        layer6[15][31:24] = 'd0;
        layer6[15][39:32] = 'd0;
        layer6[15][47:40] = 'd0;
        layer6[15][55:48] = 'd0;
    end
  endcase
end

wire  [39:0]  kernel_img_mul_0[0:48];
assign kernel_img_mul_0[0] = layer0[0][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_0[1] = layer0[0][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_0[2] = layer0[0][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_0[3] = layer0[0][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_0[4] = layer0[0][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_0[5] = layer0[0][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_0[6] = layer0[0][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_0[7] = layer1[0][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_0[8] = layer1[0][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_0[9] = layer1[0][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_0[10] = layer1[0][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_0[11] = layer1[0][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_0[12] = layer1[0][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_0[13] = layer1[0][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_0[14] = layer2[0][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_0[15] = layer2[0][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_0[16] = layer2[0][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_0[17] = layer2[0][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_0[18] = layer2[0][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_0[19] = layer2[0][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_0[20] = layer2[0][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_0[21] = layer3[0][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_0[22] = layer3[0][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_0[23] = layer3[0][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_0[24] = layer3[0][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_0[25] = layer3[0][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_0[26] = layer3[0][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_0[27] = layer3[0][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_0[28] = layer4[0][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_0[29] = layer4[0][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_0[30] = layer4[0][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_0[31] = layer4[0][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_0[32] = layer4[0][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_0[33] = layer4[0][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_0[34] = layer4[0][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_0[35] = layer5[0][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_0[36] = layer5[0][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_0[37] = layer5[0][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_0[38] = layer5[0][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_0[39] = layer5[0][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_0[40] = layer5[0][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_0[41] = layer5[0][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_0[42] = layer6[0][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_0[43] = layer6[0][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_0[44] = layer6[0][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_0[45] = layer6[0][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_0[46] = layer6[0][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_0[47] = layer6[0][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_0[48] = layer6[0][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_0 = kernel_img_mul_0[0] + kernel_img_mul_0[1] + kernel_img_mul_0[2] + 
                kernel_img_mul_0[3] + kernel_img_mul_0[4] + kernel_img_mul_0[5] + 
                kernel_img_mul_0[6] + kernel_img_mul_0[7] + kernel_img_mul_0[8] + 
                kernel_img_mul_0[9] + kernel_img_mul_0[10] + kernel_img_mul_0[11] + 
                kernel_img_mul_0[12] + kernel_img_mul_0[13] + kernel_img_mul_0[14] + 
                kernel_img_mul_0[15] + kernel_img_mul_0[16] + kernel_img_mul_0[17] + 
                kernel_img_mul_0[18] + kernel_img_mul_0[19] + kernel_img_mul_0[20] + 
                kernel_img_mul_0[21] + kernel_img_mul_0[22] + kernel_img_mul_0[23] + 
                kernel_img_mul_0[24] + kernel_img_mul_0[25] + kernel_img_mul_0[26] + 
                kernel_img_mul_0[27] + kernel_img_mul_0[28] + kernel_img_mul_0[29] + 
                kernel_img_mul_0[30] + kernel_img_mul_0[31] + kernel_img_mul_0[32] + 
                kernel_img_mul_0[33] + kernel_img_mul_0[34] + kernel_img_mul_0[35] + 
                kernel_img_mul_0[36] + kernel_img_mul_0[37] + kernel_img_mul_0[38] + 
                kernel_img_mul_0[39] + kernel_img_mul_0[40] + kernel_img_mul_0[41] + 
                kernel_img_mul_0[42] + kernel_img_mul_0[43] + kernel_img_mul_0[44] + 
                kernel_img_mul_0[45] + kernel_img_mul_0[46] + kernel_img_mul_0[47] + 
                kernel_img_mul_0[48];
wire  [39:0]  kernel_img_mul_1[0:48];
assign kernel_img_mul_1[0] = layer0[1][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_1[1] = layer0[1][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_1[2] = layer0[1][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_1[3] = layer0[1][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_1[4] = layer0[1][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_1[5] = layer0[1][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_1[6] = layer0[1][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_1[7] = layer1[1][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_1[8] = layer1[1][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_1[9] = layer1[1][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_1[10] = layer1[1][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_1[11] = layer1[1][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_1[12] = layer1[1][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_1[13] = layer1[1][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_1[14] = layer2[1][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_1[15] = layer2[1][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_1[16] = layer2[1][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_1[17] = layer2[1][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_1[18] = layer2[1][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_1[19] = layer2[1][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_1[20] = layer2[1][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_1[21] = layer3[1][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_1[22] = layer3[1][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_1[23] = layer3[1][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_1[24] = layer3[1][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_1[25] = layer3[1][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_1[26] = layer3[1][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_1[27] = layer3[1][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_1[28] = layer4[1][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_1[29] = layer4[1][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_1[30] = layer4[1][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_1[31] = layer4[1][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_1[32] = layer4[1][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_1[33] = layer4[1][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_1[34] = layer4[1][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_1[35] = layer5[1][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_1[36] = layer5[1][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_1[37] = layer5[1][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_1[38] = layer5[1][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_1[39] = layer5[1][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_1[40] = layer5[1][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_1[41] = layer5[1][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_1[42] = layer6[1][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_1[43] = layer6[1][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_1[44] = layer6[1][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_1[45] = layer6[1][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_1[46] = layer6[1][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_1[47] = layer6[1][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_1[48] = layer6[1][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_1 = kernel_img_mul_1[0] + kernel_img_mul_1[1] + kernel_img_mul_1[2] + 
                kernel_img_mul_1[3] + kernel_img_mul_1[4] + kernel_img_mul_1[5] + 
                kernel_img_mul_1[6] + kernel_img_mul_1[7] + kernel_img_mul_1[8] + 
                kernel_img_mul_1[9] + kernel_img_mul_1[10] + kernel_img_mul_1[11] + 
                kernel_img_mul_1[12] + kernel_img_mul_1[13] + kernel_img_mul_1[14] + 
                kernel_img_mul_1[15] + kernel_img_mul_1[16] + kernel_img_mul_1[17] + 
                kernel_img_mul_1[18] + kernel_img_mul_1[19] + kernel_img_mul_1[20] + 
                kernel_img_mul_1[21] + kernel_img_mul_1[22] + kernel_img_mul_1[23] + 
                kernel_img_mul_1[24] + kernel_img_mul_1[25] + kernel_img_mul_1[26] + 
                kernel_img_mul_1[27] + kernel_img_mul_1[28] + kernel_img_mul_1[29] + 
                kernel_img_mul_1[30] + kernel_img_mul_1[31] + kernel_img_mul_1[32] + 
                kernel_img_mul_1[33] + kernel_img_mul_1[34] + kernel_img_mul_1[35] + 
                kernel_img_mul_1[36] + kernel_img_mul_1[37] + kernel_img_mul_1[38] + 
                kernel_img_mul_1[39] + kernel_img_mul_1[40] + kernel_img_mul_1[41] + 
                kernel_img_mul_1[42] + kernel_img_mul_1[43] + kernel_img_mul_1[44] + 
                kernel_img_mul_1[45] + kernel_img_mul_1[46] + kernel_img_mul_1[47] + 
                kernel_img_mul_1[48];
wire  [39:0]  kernel_img_mul_2[0:48];
assign kernel_img_mul_2[0] = layer0[2][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_2[1] = layer0[2][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_2[2] = layer0[2][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_2[3] = layer0[2][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_2[4] = layer0[2][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_2[5] = layer0[2][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_2[6] = layer0[2][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_2[7] = layer1[2][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_2[8] = layer1[2][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_2[9] = layer1[2][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_2[10] = layer1[2][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_2[11] = layer1[2][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_2[12] = layer1[2][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_2[13] = layer1[2][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_2[14] = layer2[2][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_2[15] = layer2[2][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_2[16] = layer2[2][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_2[17] = layer2[2][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_2[18] = layer2[2][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_2[19] = layer2[2][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_2[20] = layer2[2][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_2[21] = layer3[2][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_2[22] = layer3[2][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_2[23] = layer3[2][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_2[24] = layer3[2][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_2[25] = layer3[2][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_2[26] = layer3[2][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_2[27] = layer3[2][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_2[28] = layer4[2][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_2[29] = layer4[2][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_2[30] = layer4[2][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_2[31] = layer4[2][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_2[32] = layer4[2][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_2[33] = layer4[2][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_2[34] = layer4[2][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_2[35] = layer5[2][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_2[36] = layer5[2][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_2[37] = layer5[2][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_2[38] = layer5[2][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_2[39] = layer5[2][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_2[40] = layer5[2][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_2[41] = layer5[2][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_2[42] = layer6[2][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_2[43] = layer6[2][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_2[44] = layer6[2][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_2[45] = layer6[2][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_2[46] = layer6[2][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_2[47] = layer6[2][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_2[48] = layer6[2][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_2 = kernel_img_mul_2[0] + kernel_img_mul_2[1] + kernel_img_mul_2[2] + 
                kernel_img_mul_2[3] + kernel_img_mul_2[4] + kernel_img_mul_2[5] + 
                kernel_img_mul_2[6] + kernel_img_mul_2[7] + kernel_img_mul_2[8] + 
                kernel_img_mul_2[9] + kernel_img_mul_2[10] + kernel_img_mul_2[11] + 
                kernel_img_mul_2[12] + kernel_img_mul_2[13] + kernel_img_mul_2[14] + 
                kernel_img_mul_2[15] + kernel_img_mul_2[16] + kernel_img_mul_2[17] + 
                kernel_img_mul_2[18] + kernel_img_mul_2[19] + kernel_img_mul_2[20] + 
                kernel_img_mul_2[21] + kernel_img_mul_2[22] + kernel_img_mul_2[23] + 
                kernel_img_mul_2[24] + kernel_img_mul_2[25] + kernel_img_mul_2[26] + 
                kernel_img_mul_2[27] + kernel_img_mul_2[28] + kernel_img_mul_2[29] + 
                kernel_img_mul_2[30] + kernel_img_mul_2[31] + kernel_img_mul_2[32] + 
                kernel_img_mul_2[33] + kernel_img_mul_2[34] + kernel_img_mul_2[35] + 
                kernel_img_mul_2[36] + kernel_img_mul_2[37] + kernel_img_mul_2[38] + 
                kernel_img_mul_2[39] + kernel_img_mul_2[40] + kernel_img_mul_2[41] + 
                kernel_img_mul_2[42] + kernel_img_mul_2[43] + kernel_img_mul_2[44] + 
                kernel_img_mul_2[45] + kernel_img_mul_2[46] + kernel_img_mul_2[47] + 
                kernel_img_mul_2[48];
wire  [39:0]  kernel_img_mul_3[0:48];
assign kernel_img_mul_3[0] = layer0[3][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_3[1] = layer0[3][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_3[2] = layer0[3][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_3[3] = layer0[3][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_3[4] = layer0[3][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_3[5] = layer0[3][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_3[6] = layer0[3][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_3[7] = layer1[3][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_3[8] = layer1[3][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_3[9] = layer1[3][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_3[10] = layer1[3][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_3[11] = layer1[3][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_3[12] = layer1[3][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_3[13] = layer1[3][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_3[14] = layer2[3][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_3[15] = layer2[3][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_3[16] = layer2[3][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_3[17] = layer2[3][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_3[18] = layer2[3][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_3[19] = layer2[3][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_3[20] = layer2[3][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_3[21] = layer3[3][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_3[22] = layer3[3][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_3[23] = layer3[3][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_3[24] = layer3[3][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_3[25] = layer3[3][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_3[26] = layer3[3][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_3[27] = layer3[3][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_3[28] = layer4[3][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_3[29] = layer4[3][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_3[30] = layer4[3][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_3[31] = layer4[3][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_3[32] = layer4[3][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_3[33] = layer4[3][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_3[34] = layer4[3][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_3[35] = layer5[3][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_3[36] = layer5[3][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_3[37] = layer5[3][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_3[38] = layer5[3][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_3[39] = layer5[3][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_3[40] = layer5[3][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_3[41] = layer5[3][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_3[42] = layer6[3][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_3[43] = layer6[3][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_3[44] = layer6[3][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_3[45] = layer6[3][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_3[46] = layer6[3][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_3[47] = layer6[3][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_3[48] = layer6[3][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_3 = kernel_img_mul_3[0] + kernel_img_mul_3[1] + kernel_img_mul_3[2] + 
                kernel_img_mul_3[3] + kernel_img_mul_3[4] + kernel_img_mul_3[5] + 
                kernel_img_mul_3[6] + kernel_img_mul_3[7] + kernel_img_mul_3[8] + 
                kernel_img_mul_3[9] + kernel_img_mul_3[10] + kernel_img_mul_3[11] + 
                kernel_img_mul_3[12] + kernel_img_mul_3[13] + kernel_img_mul_3[14] + 
                kernel_img_mul_3[15] + kernel_img_mul_3[16] + kernel_img_mul_3[17] + 
                kernel_img_mul_3[18] + kernel_img_mul_3[19] + kernel_img_mul_3[20] + 
                kernel_img_mul_3[21] + kernel_img_mul_3[22] + kernel_img_mul_3[23] + 
                kernel_img_mul_3[24] + kernel_img_mul_3[25] + kernel_img_mul_3[26] + 
                kernel_img_mul_3[27] + kernel_img_mul_3[28] + kernel_img_mul_3[29] + 
                kernel_img_mul_3[30] + kernel_img_mul_3[31] + kernel_img_mul_3[32] + 
                kernel_img_mul_3[33] + kernel_img_mul_3[34] + kernel_img_mul_3[35] + 
                kernel_img_mul_3[36] + kernel_img_mul_3[37] + kernel_img_mul_3[38] + 
                kernel_img_mul_3[39] + kernel_img_mul_3[40] + kernel_img_mul_3[41] + 
                kernel_img_mul_3[42] + kernel_img_mul_3[43] + kernel_img_mul_3[44] + 
                kernel_img_mul_3[45] + kernel_img_mul_3[46] + kernel_img_mul_3[47] + 
                kernel_img_mul_3[48];
wire  [39:0]  kernel_img_mul_4[0:48];
assign kernel_img_mul_4[0] = layer0[4][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_4[1] = layer0[4][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_4[2] = layer0[4][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_4[3] = layer0[4][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_4[4] = layer0[4][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_4[5] = layer0[4][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_4[6] = layer0[4][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_4[7] = layer1[4][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_4[8] = layer1[4][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_4[9] = layer1[4][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_4[10] = layer1[4][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_4[11] = layer1[4][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_4[12] = layer1[4][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_4[13] = layer1[4][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_4[14] = layer2[4][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_4[15] = layer2[4][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_4[16] = layer2[4][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_4[17] = layer2[4][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_4[18] = layer2[4][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_4[19] = layer2[4][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_4[20] = layer2[4][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_4[21] = layer3[4][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_4[22] = layer3[4][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_4[23] = layer3[4][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_4[24] = layer3[4][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_4[25] = layer3[4][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_4[26] = layer3[4][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_4[27] = layer3[4][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_4[28] = layer4[4][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_4[29] = layer4[4][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_4[30] = layer4[4][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_4[31] = layer4[4][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_4[32] = layer4[4][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_4[33] = layer4[4][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_4[34] = layer4[4][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_4[35] = layer5[4][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_4[36] = layer5[4][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_4[37] = layer5[4][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_4[38] = layer5[4][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_4[39] = layer5[4][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_4[40] = layer5[4][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_4[41] = layer5[4][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_4[42] = layer6[4][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_4[43] = layer6[4][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_4[44] = layer6[4][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_4[45] = layer6[4][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_4[46] = layer6[4][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_4[47] = layer6[4][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_4[48] = layer6[4][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_4 = kernel_img_mul_4[0] + kernel_img_mul_4[1] + kernel_img_mul_4[2] + 
                kernel_img_mul_4[3] + kernel_img_mul_4[4] + kernel_img_mul_4[5] + 
                kernel_img_mul_4[6] + kernel_img_mul_4[7] + kernel_img_mul_4[8] + 
                kernel_img_mul_4[9] + kernel_img_mul_4[10] + kernel_img_mul_4[11] + 
                kernel_img_mul_4[12] + kernel_img_mul_4[13] + kernel_img_mul_4[14] + 
                kernel_img_mul_4[15] + kernel_img_mul_4[16] + kernel_img_mul_4[17] + 
                kernel_img_mul_4[18] + kernel_img_mul_4[19] + kernel_img_mul_4[20] + 
                kernel_img_mul_4[21] + kernel_img_mul_4[22] + kernel_img_mul_4[23] + 
                kernel_img_mul_4[24] + kernel_img_mul_4[25] + kernel_img_mul_4[26] + 
                kernel_img_mul_4[27] + kernel_img_mul_4[28] + kernel_img_mul_4[29] + 
                kernel_img_mul_4[30] + kernel_img_mul_4[31] + kernel_img_mul_4[32] + 
                kernel_img_mul_4[33] + kernel_img_mul_4[34] + kernel_img_mul_4[35] + 
                kernel_img_mul_4[36] + kernel_img_mul_4[37] + kernel_img_mul_4[38] + 
                kernel_img_mul_4[39] + kernel_img_mul_4[40] + kernel_img_mul_4[41] + 
                kernel_img_mul_4[42] + kernel_img_mul_4[43] + kernel_img_mul_4[44] + 
                kernel_img_mul_4[45] + kernel_img_mul_4[46] + kernel_img_mul_4[47] + 
                kernel_img_mul_4[48];
wire  [39:0]  kernel_img_mul_5[0:48];
assign kernel_img_mul_5[0] = layer0[5][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_5[1] = layer0[5][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_5[2] = layer0[5][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_5[3] = layer0[5][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_5[4] = layer0[5][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_5[5] = layer0[5][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_5[6] = layer0[5][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_5[7] = layer1[5][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_5[8] = layer1[5][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_5[9] = layer1[5][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_5[10] = layer1[5][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_5[11] = layer1[5][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_5[12] = layer1[5][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_5[13] = layer1[5][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_5[14] = layer2[5][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_5[15] = layer2[5][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_5[16] = layer2[5][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_5[17] = layer2[5][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_5[18] = layer2[5][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_5[19] = layer2[5][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_5[20] = layer2[5][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_5[21] = layer3[5][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_5[22] = layer3[5][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_5[23] = layer3[5][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_5[24] = layer3[5][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_5[25] = layer3[5][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_5[26] = layer3[5][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_5[27] = layer3[5][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_5[28] = layer4[5][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_5[29] = layer4[5][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_5[30] = layer4[5][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_5[31] = layer4[5][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_5[32] = layer4[5][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_5[33] = layer4[5][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_5[34] = layer4[5][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_5[35] = layer5[5][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_5[36] = layer5[5][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_5[37] = layer5[5][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_5[38] = layer5[5][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_5[39] = layer5[5][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_5[40] = layer5[5][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_5[41] = layer5[5][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_5[42] = layer6[5][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_5[43] = layer6[5][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_5[44] = layer6[5][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_5[45] = layer6[5][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_5[46] = layer6[5][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_5[47] = layer6[5][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_5[48] = layer6[5][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_5 = kernel_img_mul_5[0] + kernel_img_mul_5[1] + kernel_img_mul_5[2] + 
                kernel_img_mul_5[3] + kernel_img_mul_5[4] + kernel_img_mul_5[5] + 
                kernel_img_mul_5[6] + kernel_img_mul_5[7] + kernel_img_mul_5[8] + 
                kernel_img_mul_5[9] + kernel_img_mul_5[10] + kernel_img_mul_5[11] + 
                kernel_img_mul_5[12] + kernel_img_mul_5[13] + kernel_img_mul_5[14] + 
                kernel_img_mul_5[15] + kernel_img_mul_5[16] + kernel_img_mul_5[17] + 
                kernel_img_mul_5[18] + kernel_img_mul_5[19] + kernel_img_mul_5[20] + 
                kernel_img_mul_5[21] + kernel_img_mul_5[22] + kernel_img_mul_5[23] + 
                kernel_img_mul_5[24] + kernel_img_mul_5[25] + kernel_img_mul_5[26] + 
                kernel_img_mul_5[27] + kernel_img_mul_5[28] + kernel_img_mul_5[29] + 
                kernel_img_mul_5[30] + kernel_img_mul_5[31] + kernel_img_mul_5[32] + 
                kernel_img_mul_5[33] + kernel_img_mul_5[34] + kernel_img_mul_5[35] + 
                kernel_img_mul_5[36] + kernel_img_mul_5[37] + kernel_img_mul_5[38] + 
                kernel_img_mul_5[39] + kernel_img_mul_5[40] + kernel_img_mul_5[41] + 
                kernel_img_mul_5[42] + kernel_img_mul_5[43] + kernel_img_mul_5[44] + 
                kernel_img_mul_5[45] + kernel_img_mul_5[46] + kernel_img_mul_5[47] + 
                kernel_img_mul_5[48];
wire  [39:0]  kernel_img_mul_6[0:48];
assign kernel_img_mul_6[0] = layer0[6][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_6[1] = layer0[6][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_6[2] = layer0[6][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_6[3] = layer0[6][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_6[4] = layer0[6][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_6[5] = layer0[6][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_6[6] = layer0[6][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_6[7] = layer1[6][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_6[8] = layer1[6][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_6[9] = layer1[6][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_6[10] = layer1[6][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_6[11] = layer1[6][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_6[12] = layer1[6][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_6[13] = layer1[6][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_6[14] = layer2[6][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_6[15] = layer2[6][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_6[16] = layer2[6][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_6[17] = layer2[6][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_6[18] = layer2[6][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_6[19] = layer2[6][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_6[20] = layer2[6][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_6[21] = layer3[6][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_6[22] = layer3[6][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_6[23] = layer3[6][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_6[24] = layer3[6][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_6[25] = layer3[6][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_6[26] = layer3[6][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_6[27] = layer3[6][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_6[28] = layer4[6][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_6[29] = layer4[6][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_6[30] = layer4[6][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_6[31] = layer4[6][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_6[32] = layer4[6][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_6[33] = layer4[6][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_6[34] = layer4[6][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_6[35] = layer5[6][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_6[36] = layer5[6][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_6[37] = layer5[6][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_6[38] = layer5[6][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_6[39] = layer5[6][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_6[40] = layer5[6][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_6[41] = layer5[6][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_6[42] = layer6[6][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_6[43] = layer6[6][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_6[44] = layer6[6][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_6[45] = layer6[6][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_6[46] = layer6[6][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_6[47] = layer6[6][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_6[48] = layer6[6][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_6 = kernel_img_mul_6[0] + kernel_img_mul_6[1] + kernel_img_mul_6[2] + 
                kernel_img_mul_6[3] + kernel_img_mul_6[4] + kernel_img_mul_6[5] + 
                kernel_img_mul_6[6] + kernel_img_mul_6[7] + kernel_img_mul_6[8] + 
                kernel_img_mul_6[9] + kernel_img_mul_6[10] + kernel_img_mul_6[11] + 
                kernel_img_mul_6[12] + kernel_img_mul_6[13] + kernel_img_mul_6[14] + 
                kernel_img_mul_6[15] + kernel_img_mul_6[16] + kernel_img_mul_6[17] + 
                kernel_img_mul_6[18] + kernel_img_mul_6[19] + kernel_img_mul_6[20] + 
                kernel_img_mul_6[21] + kernel_img_mul_6[22] + kernel_img_mul_6[23] + 
                kernel_img_mul_6[24] + kernel_img_mul_6[25] + kernel_img_mul_6[26] + 
                kernel_img_mul_6[27] + kernel_img_mul_6[28] + kernel_img_mul_6[29] + 
                kernel_img_mul_6[30] + kernel_img_mul_6[31] + kernel_img_mul_6[32] + 
                kernel_img_mul_6[33] + kernel_img_mul_6[34] + kernel_img_mul_6[35] + 
                kernel_img_mul_6[36] + kernel_img_mul_6[37] + kernel_img_mul_6[38] + 
                kernel_img_mul_6[39] + kernel_img_mul_6[40] + kernel_img_mul_6[41] + 
                kernel_img_mul_6[42] + kernel_img_mul_6[43] + kernel_img_mul_6[44] + 
                kernel_img_mul_6[45] + kernel_img_mul_6[46] + kernel_img_mul_6[47] + 
                kernel_img_mul_6[48];
wire  [39:0]  kernel_img_mul_7[0:48];
assign kernel_img_mul_7[0] = layer0[7][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_7[1] = layer0[7][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_7[2] = layer0[7][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_7[3] = layer0[7][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_7[4] = layer0[7][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_7[5] = layer0[7][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_7[6] = layer0[7][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_7[7] = layer1[7][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_7[8] = layer1[7][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_7[9] = layer1[7][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_7[10] = layer1[7][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_7[11] = layer1[7][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_7[12] = layer1[7][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_7[13] = layer1[7][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_7[14] = layer2[7][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_7[15] = layer2[7][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_7[16] = layer2[7][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_7[17] = layer2[7][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_7[18] = layer2[7][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_7[19] = layer2[7][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_7[20] = layer2[7][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_7[21] = layer3[7][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_7[22] = layer3[7][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_7[23] = layer3[7][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_7[24] = layer3[7][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_7[25] = layer3[7][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_7[26] = layer3[7][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_7[27] = layer3[7][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_7[28] = layer4[7][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_7[29] = layer4[7][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_7[30] = layer4[7][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_7[31] = layer4[7][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_7[32] = layer4[7][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_7[33] = layer4[7][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_7[34] = layer4[7][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_7[35] = layer5[7][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_7[36] = layer5[7][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_7[37] = layer5[7][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_7[38] = layer5[7][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_7[39] = layer5[7][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_7[40] = layer5[7][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_7[41] = layer5[7][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_7[42] = layer6[7][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_7[43] = layer6[7][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_7[44] = layer6[7][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_7[45] = layer6[7][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_7[46] = layer6[7][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_7[47] = layer6[7][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_7[48] = layer6[7][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_7 = kernel_img_mul_7[0] + kernel_img_mul_7[1] + kernel_img_mul_7[2] + 
                kernel_img_mul_7[3] + kernel_img_mul_7[4] + kernel_img_mul_7[5] + 
                kernel_img_mul_7[6] + kernel_img_mul_7[7] + kernel_img_mul_7[8] + 
                kernel_img_mul_7[9] + kernel_img_mul_7[10] + kernel_img_mul_7[11] + 
                kernel_img_mul_7[12] + kernel_img_mul_7[13] + kernel_img_mul_7[14] + 
                kernel_img_mul_7[15] + kernel_img_mul_7[16] + kernel_img_mul_7[17] + 
                kernel_img_mul_7[18] + kernel_img_mul_7[19] + kernel_img_mul_7[20] + 
                kernel_img_mul_7[21] + kernel_img_mul_7[22] + kernel_img_mul_7[23] + 
                kernel_img_mul_7[24] + kernel_img_mul_7[25] + kernel_img_mul_7[26] + 
                kernel_img_mul_7[27] + kernel_img_mul_7[28] + kernel_img_mul_7[29] + 
                kernel_img_mul_7[30] + kernel_img_mul_7[31] + kernel_img_mul_7[32] + 
                kernel_img_mul_7[33] + kernel_img_mul_7[34] + kernel_img_mul_7[35] + 
                kernel_img_mul_7[36] + kernel_img_mul_7[37] + kernel_img_mul_7[38] + 
                kernel_img_mul_7[39] + kernel_img_mul_7[40] + kernel_img_mul_7[41] + 
                kernel_img_mul_7[42] + kernel_img_mul_7[43] + kernel_img_mul_7[44] + 
                kernel_img_mul_7[45] + kernel_img_mul_7[46] + kernel_img_mul_7[47] + 
                kernel_img_mul_7[48];
wire  [39:0]  kernel_img_mul_8[0:48];
assign kernel_img_mul_8[0] = layer0[8][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_8[1] = layer0[8][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_8[2] = layer0[8][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_8[3] = layer0[8][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_8[4] = layer0[8][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_8[5] = layer0[8][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_8[6] = layer0[8][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_8[7] = layer1[8][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_8[8] = layer1[8][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_8[9] = layer1[8][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_8[10] = layer1[8][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_8[11] = layer1[8][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_8[12] = layer1[8][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_8[13] = layer1[8][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_8[14] = layer2[8][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_8[15] = layer2[8][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_8[16] = layer2[8][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_8[17] = layer2[8][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_8[18] = layer2[8][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_8[19] = layer2[8][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_8[20] = layer2[8][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_8[21] = layer3[8][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_8[22] = layer3[8][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_8[23] = layer3[8][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_8[24] = layer3[8][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_8[25] = layer3[8][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_8[26] = layer3[8][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_8[27] = layer3[8][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_8[28] = layer4[8][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_8[29] = layer4[8][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_8[30] = layer4[8][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_8[31] = layer4[8][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_8[32] = layer4[8][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_8[33] = layer4[8][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_8[34] = layer4[8][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_8[35] = layer5[8][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_8[36] = layer5[8][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_8[37] = layer5[8][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_8[38] = layer5[8][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_8[39] = layer5[8][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_8[40] = layer5[8][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_8[41] = layer5[8][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_8[42] = layer6[8][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_8[43] = layer6[8][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_8[44] = layer6[8][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_8[45] = layer6[8][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_8[46] = layer6[8][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_8[47] = layer6[8][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_8[48] = layer6[8][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_8 = kernel_img_mul_8[0] + kernel_img_mul_8[1] + kernel_img_mul_8[2] + 
                kernel_img_mul_8[3] + kernel_img_mul_8[4] + kernel_img_mul_8[5] + 
                kernel_img_mul_8[6] + kernel_img_mul_8[7] + kernel_img_mul_8[8] + 
                kernel_img_mul_8[9] + kernel_img_mul_8[10] + kernel_img_mul_8[11] + 
                kernel_img_mul_8[12] + kernel_img_mul_8[13] + kernel_img_mul_8[14] + 
                kernel_img_mul_8[15] + kernel_img_mul_8[16] + kernel_img_mul_8[17] + 
                kernel_img_mul_8[18] + kernel_img_mul_8[19] + kernel_img_mul_8[20] + 
                kernel_img_mul_8[21] + kernel_img_mul_8[22] + kernel_img_mul_8[23] + 
                kernel_img_mul_8[24] + kernel_img_mul_8[25] + kernel_img_mul_8[26] + 
                kernel_img_mul_8[27] + kernel_img_mul_8[28] + kernel_img_mul_8[29] + 
                kernel_img_mul_8[30] + kernel_img_mul_8[31] + kernel_img_mul_8[32] + 
                kernel_img_mul_8[33] + kernel_img_mul_8[34] + kernel_img_mul_8[35] + 
                kernel_img_mul_8[36] + kernel_img_mul_8[37] + kernel_img_mul_8[38] + 
                kernel_img_mul_8[39] + kernel_img_mul_8[40] + kernel_img_mul_8[41] + 
                kernel_img_mul_8[42] + kernel_img_mul_8[43] + kernel_img_mul_8[44] + 
                kernel_img_mul_8[45] + kernel_img_mul_8[46] + kernel_img_mul_8[47] + 
                kernel_img_mul_8[48];
wire  [39:0]  kernel_img_mul_9[0:48];
assign kernel_img_mul_9[0] = layer0[9][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_9[1] = layer0[9][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_9[2] = layer0[9][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_9[3] = layer0[9][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_9[4] = layer0[9][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_9[5] = layer0[9][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_9[6] = layer0[9][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_9[7] = layer1[9][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_9[8] = layer1[9][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_9[9] = layer1[9][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_9[10] = layer1[9][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_9[11] = layer1[9][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_9[12] = layer1[9][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_9[13] = layer1[9][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_9[14] = layer2[9][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_9[15] = layer2[9][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_9[16] = layer2[9][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_9[17] = layer2[9][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_9[18] = layer2[9][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_9[19] = layer2[9][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_9[20] = layer2[9][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_9[21] = layer3[9][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_9[22] = layer3[9][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_9[23] = layer3[9][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_9[24] = layer3[9][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_9[25] = layer3[9][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_9[26] = layer3[9][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_9[27] = layer3[9][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_9[28] = layer4[9][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_9[29] = layer4[9][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_9[30] = layer4[9][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_9[31] = layer4[9][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_9[32] = layer4[9][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_9[33] = layer4[9][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_9[34] = layer4[9][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_9[35] = layer5[9][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_9[36] = layer5[9][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_9[37] = layer5[9][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_9[38] = layer5[9][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_9[39] = layer5[9][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_9[40] = layer5[9][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_9[41] = layer5[9][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_9[42] = layer6[9][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_9[43] = layer6[9][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_9[44] = layer6[9][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_9[45] = layer6[9][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_9[46] = layer6[9][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_9[47] = layer6[9][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_9[48] = layer6[9][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_9 = kernel_img_mul_9[0] + kernel_img_mul_9[1] + kernel_img_mul_9[2] + 
                kernel_img_mul_9[3] + kernel_img_mul_9[4] + kernel_img_mul_9[5] + 
                kernel_img_mul_9[6] + kernel_img_mul_9[7] + kernel_img_mul_9[8] + 
                kernel_img_mul_9[9] + kernel_img_mul_9[10] + kernel_img_mul_9[11] + 
                kernel_img_mul_9[12] + kernel_img_mul_9[13] + kernel_img_mul_9[14] + 
                kernel_img_mul_9[15] + kernel_img_mul_9[16] + kernel_img_mul_9[17] + 
                kernel_img_mul_9[18] + kernel_img_mul_9[19] + kernel_img_mul_9[20] + 
                kernel_img_mul_9[21] + kernel_img_mul_9[22] + kernel_img_mul_9[23] + 
                kernel_img_mul_9[24] + kernel_img_mul_9[25] + kernel_img_mul_9[26] + 
                kernel_img_mul_9[27] + kernel_img_mul_9[28] + kernel_img_mul_9[29] + 
                kernel_img_mul_9[30] + kernel_img_mul_9[31] + kernel_img_mul_9[32] + 
                kernel_img_mul_9[33] + kernel_img_mul_9[34] + kernel_img_mul_9[35] + 
                kernel_img_mul_9[36] + kernel_img_mul_9[37] + kernel_img_mul_9[38] + 
                kernel_img_mul_9[39] + kernel_img_mul_9[40] + kernel_img_mul_9[41] + 
                kernel_img_mul_9[42] + kernel_img_mul_9[43] + kernel_img_mul_9[44] + 
                kernel_img_mul_9[45] + kernel_img_mul_9[46] + kernel_img_mul_9[47] + 
                kernel_img_mul_9[48];
wire  [39:0]  kernel_img_mul_10[0:48];
assign kernel_img_mul_10[0] = layer0[10][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_10[1] = layer0[10][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_10[2] = layer0[10][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_10[3] = layer0[10][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_10[4] = layer0[10][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_10[5] = layer0[10][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_10[6] = layer0[10][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_10[7] = layer1[10][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_10[8] = layer1[10][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_10[9] = layer1[10][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_10[10] = layer1[10][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_10[11] = layer1[10][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_10[12] = layer1[10][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_10[13] = layer1[10][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_10[14] = layer2[10][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_10[15] = layer2[10][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_10[16] = layer2[10][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_10[17] = layer2[10][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_10[18] = layer2[10][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_10[19] = layer2[10][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_10[20] = layer2[10][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_10[21] = layer3[10][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_10[22] = layer3[10][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_10[23] = layer3[10][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_10[24] = layer3[10][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_10[25] = layer3[10][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_10[26] = layer3[10][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_10[27] = layer3[10][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_10[28] = layer4[10][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_10[29] = layer4[10][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_10[30] = layer4[10][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_10[31] = layer4[10][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_10[32] = layer4[10][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_10[33] = layer4[10][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_10[34] = layer4[10][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_10[35] = layer5[10][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_10[36] = layer5[10][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_10[37] = layer5[10][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_10[38] = layer5[10][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_10[39] = layer5[10][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_10[40] = layer5[10][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_10[41] = layer5[10][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_10[42] = layer6[10][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_10[43] = layer6[10][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_10[44] = layer6[10][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_10[45] = layer6[10][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_10[46] = layer6[10][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_10[47] = layer6[10][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_10[48] = layer6[10][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_10 = kernel_img_mul_10[0] + kernel_img_mul_10[1] + kernel_img_mul_10[2] + 
                kernel_img_mul_10[3] + kernel_img_mul_10[4] + kernel_img_mul_10[5] + 
                kernel_img_mul_10[6] + kernel_img_mul_10[7] + kernel_img_mul_10[8] + 
                kernel_img_mul_10[9] + kernel_img_mul_10[10] + kernel_img_mul_10[11] + 
                kernel_img_mul_10[12] + kernel_img_mul_10[13] + kernel_img_mul_10[14] + 
                kernel_img_mul_10[15] + kernel_img_mul_10[16] + kernel_img_mul_10[17] + 
                kernel_img_mul_10[18] + kernel_img_mul_10[19] + kernel_img_mul_10[20] + 
                kernel_img_mul_10[21] + kernel_img_mul_10[22] + kernel_img_mul_10[23] + 
                kernel_img_mul_10[24] + kernel_img_mul_10[25] + kernel_img_mul_10[26] + 
                kernel_img_mul_10[27] + kernel_img_mul_10[28] + kernel_img_mul_10[29] + 
                kernel_img_mul_10[30] + kernel_img_mul_10[31] + kernel_img_mul_10[32] + 
                kernel_img_mul_10[33] + kernel_img_mul_10[34] + kernel_img_mul_10[35] + 
                kernel_img_mul_10[36] + kernel_img_mul_10[37] + kernel_img_mul_10[38] + 
                kernel_img_mul_10[39] + kernel_img_mul_10[40] + kernel_img_mul_10[41] + 
                kernel_img_mul_10[42] + kernel_img_mul_10[43] + kernel_img_mul_10[44] + 
                kernel_img_mul_10[45] + kernel_img_mul_10[46] + kernel_img_mul_10[47] + 
                kernel_img_mul_10[48];
wire  [39:0]  kernel_img_mul_11[0:48];
assign kernel_img_mul_11[0] = layer0[11][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_11[1] = layer0[11][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_11[2] = layer0[11][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_11[3] = layer0[11][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_11[4] = layer0[11][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_11[5] = layer0[11][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_11[6] = layer0[11][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_11[7] = layer1[11][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_11[8] = layer1[11][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_11[9] = layer1[11][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_11[10] = layer1[11][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_11[11] = layer1[11][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_11[12] = layer1[11][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_11[13] = layer1[11][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_11[14] = layer2[11][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_11[15] = layer2[11][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_11[16] = layer2[11][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_11[17] = layer2[11][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_11[18] = layer2[11][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_11[19] = layer2[11][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_11[20] = layer2[11][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_11[21] = layer3[11][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_11[22] = layer3[11][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_11[23] = layer3[11][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_11[24] = layer3[11][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_11[25] = layer3[11][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_11[26] = layer3[11][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_11[27] = layer3[11][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_11[28] = layer4[11][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_11[29] = layer4[11][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_11[30] = layer4[11][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_11[31] = layer4[11][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_11[32] = layer4[11][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_11[33] = layer4[11][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_11[34] = layer4[11][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_11[35] = layer5[11][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_11[36] = layer5[11][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_11[37] = layer5[11][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_11[38] = layer5[11][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_11[39] = layer5[11][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_11[40] = layer5[11][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_11[41] = layer5[11][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_11[42] = layer6[11][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_11[43] = layer6[11][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_11[44] = layer6[11][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_11[45] = layer6[11][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_11[46] = layer6[11][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_11[47] = layer6[11][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_11[48] = layer6[11][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_11 = kernel_img_mul_11[0] + kernel_img_mul_11[1] + kernel_img_mul_11[2] + 
                kernel_img_mul_11[3] + kernel_img_mul_11[4] + kernel_img_mul_11[5] + 
                kernel_img_mul_11[6] + kernel_img_mul_11[7] + kernel_img_mul_11[8] + 
                kernel_img_mul_11[9] + kernel_img_mul_11[10] + kernel_img_mul_11[11] + 
                kernel_img_mul_11[12] + kernel_img_mul_11[13] + kernel_img_mul_11[14] + 
                kernel_img_mul_11[15] + kernel_img_mul_11[16] + kernel_img_mul_11[17] + 
                kernel_img_mul_11[18] + kernel_img_mul_11[19] + kernel_img_mul_11[20] + 
                kernel_img_mul_11[21] + kernel_img_mul_11[22] + kernel_img_mul_11[23] + 
                kernel_img_mul_11[24] + kernel_img_mul_11[25] + kernel_img_mul_11[26] + 
                kernel_img_mul_11[27] + kernel_img_mul_11[28] + kernel_img_mul_11[29] + 
                kernel_img_mul_11[30] + kernel_img_mul_11[31] + kernel_img_mul_11[32] + 
                kernel_img_mul_11[33] + kernel_img_mul_11[34] + kernel_img_mul_11[35] + 
                kernel_img_mul_11[36] + kernel_img_mul_11[37] + kernel_img_mul_11[38] + 
                kernel_img_mul_11[39] + kernel_img_mul_11[40] + kernel_img_mul_11[41] + 
                kernel_img_mul_11[42] + kernel_img_mul_11[43] + kernel_img_mul_11[44] + 
                kernel_img_mul_11[45] + kernel_img_mul_11[46] + kernel_img_mul_11[47] + 
                kernel_img_mul_11[48];
wire  [39:0]  kernel_img_mul_12[0:48];
assign kernel_img_mul_12[0] = layer0[12][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_12[1] = layer0[12][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_12[2] = layer0[12][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_12[3] = layer0[12][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_12[4] = layer0[12][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_12[5] = layer0[12][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_12[6] = layer0[12][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_12[7] = layer1[12][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_12[8] = layer1[12][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_12[9] = layer1[12][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_12[10] = layer1[12][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_12[11] = layer1[12][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_12[12] = layer1[12][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_12[13] = layer1[12][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_12[14] = layer2[12][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_12[15] = layer2[12][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_12[16] = layer2[12][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_12[17] = layer2[12][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_12[18] = layer2[12][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_12[19] = layer2[12][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_12[20] = layer2[12][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_12[21] = layer3[12][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_12[22] = layer3[12][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_12[23] = layer3[12][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_12[24] = layer3[12][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_12[25] = layer3[12][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_12[26] = layer3[12][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_12[27] = layer3[12][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_12[28] = layer4[12][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_12[29] = layer4[12][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_12[30] = layer4[12][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_12[31] = layer4[12][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_12[32] = layer4[12][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_12[33] = layer4[12][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_12[34] = layer4[12][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_12[35] = layer5[12][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_12[36] = layer5[12][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_12[37] = layer5[12][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_12[38] = layer5[12][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_12[39] = layer5[12][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_12[40] = layer5[12][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_12[41] = layer5[12][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_12[42] = layer6[12][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_12[43] = layer6[12][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_12[44] = layer6[12][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_12[45] = layer6[12][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_12[46] = layer6[12][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_12[47] = layer6[12][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_12[48] = layer6[12][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_12 = kernel_img_mul_12[0] + kernel_img_mul_12[1] + kernel_img_mul_12[2] + 
                kernel_img_mul_12[3] + kernel_img_mul_12[4] + kernel_img_mul_12[5] + 
                kernel_img_mul_12[6] + kernel_img_mul_12[7] + kernel_img_mul_12[8] + 
                kernel_img_mul_12[9] + kernel_img_mul_12[10] + kernel_img_mul_12[11] + 
                kernel_img_mul_12[12] + kernel_img_mul_12[13] + kernel_img_mul_12[14] + 
                kernel_img_mul_12[15] + kernel_img_mul_12[16] + kernel_img_mul_12[17] + 
                kernel_img_mul_12[18] + kernel_img_mul_12[19] + kernel_img_mul_12[20] + 
                kernel_img_mul_12[21] + kernel_img_mul_12[22] + kernel_img_mul_12[23] + 
                kernel_img_mul_12[24] + kernel_img_mul_12[25] + kernel_img_mul_12[26] + 
                kernel_img_mul_12[27] + kernel_img_mul_12[28] + kernel_img_mul_12[29] + 
                kernel_img_mul_12[30] + kernel_img_mul_12[31] + kernel_img_mul_12[32] + 
                kernel_img_mul_12[33] + kernel_img_mul_12[34] + kernel_img_mul_12[35] + 
                kernel_img_mul_12[36] + kernel_img_mul_12[37] + kernel_img_mul_12[38] + 
                kernel_img_mul_12[39] + kernel_img_mul_12[40] + kernel_img_mul_12[41] + 
                kernel_img_mul_12[42] + kernel_img_mul_12[43] + kernel_img_mul_12[44] + 
                kernel_img_mul_12[45] + kernel_img_mul_12[46] + kernel_img_mul_12[47] + 
                kernel_img_mul_12[48];
wire  [39:0]  kernel_img_mul_13[0:48];
assign kernel_img_mul_13[0] = layer0[13][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_13[1] = layer0[13][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_13[2] = layer0[13][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_13[3] = layer0[13][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_13[4] = layer0[13][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_13[5] = layer0[13][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_13[6] = layer0[13][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_13[7] = layer1[13][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_13[8] = layer1[13][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_13[9] = layer1[13][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_13[10] = layer1[13][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_13[11] = layer1[13][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_13[12] = layer1[13][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_13[13] = layer1[13][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_13[14] = layer2[13][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_13[15] = layer2[13][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_13[16] = layer2[13][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_13[17] = layer2[13][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_13[18] = layer2[13][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_13[19] = layer2[13][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_13[20] = layer2[13][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_13[21] = layer3[13][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_13[22] = layer3[13][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_13[23] = layer3[13][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_13[24] = layer3[13][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_13[25] = layer3[13][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_13[26] = layer3[13][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_13[27] = layer3[13][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_13[28] = layer4[13][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_13[29] = layer4[13][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_13[30] = layer4[13][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_13[31] = layer4[13][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_13[32] = layer4[13][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_13[33] = layer4[13][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_13[34] = layer4[13][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_13[35] = layer5[13][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_13[36] = layer5[13][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_13[37] = layer5[13][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_13[38] = layer5[13][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_13[39] = layer5[13][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_13[40] = layer5[13][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_13[41] = layer5[13][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_13[42] = layer6[13][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_13[43] = layer6[13][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_13[44] = layer6[13][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_13[45] = layer6[13][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_13[46] = layer6[13][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_13[47] = layer6[13][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_13[48] = layer6[13][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_13 = kernel_img_mul_13[0] + kernel_img_mul_13[1] + kernel_img_mul_13[2] + 
                kernel_img_mul_13[3] + kernel_img_mul_13[4] + kernel_img_mul_13[5] + 
                kernel_img_mul_13[6] + kernel_img_mul_13[7] + kernel_img_mul_13[8] + 
                kernel_img_mul_13[9] + kernel_img_mul_13[10] + kernel_img_mul_13[11] + 
                kernel_img_mul_13[12] + kernel_img_mul_13[13] + kernel_img_mul_13[14] + 
                kernel_img_mul_13[15] + kernel_img_mul_13[16] + kernel_img_mul_13[17] + 
                kernel_img_mul_13[18] + kernel_img_mul_13[19] + kernel_img_mul_13[20] + 
                kernel_img_mul_13[21] + kernel_img_mul_13[22] + kernel_img_mul_13[23] + 
                kernel_img_mul_13[24] + kernel_img_mul_13[25] + kernel_img_mul_13[26] + 
                kernel_img_mul_13[27] + kernel_img_mul_13[28] + kernel_img_mul_13[29] + 
                kernel_img_mul_13[30] + kernel_img_mul_13[31] + kernel_img_mul_13[32] + 
                kernel_img_mul_13[33] + kernel_img_mul_13[34] + kernel_img_mul_13[35] + 
                kernel_img_mul_13[36] + kernel_img_mul_13[37] + kernel_img_mul_13[38] + 
                kernel_img_mul_13[39] + kernel_img_mul_13[40] + kernel_img_mul_13[41] + 
                kernel_img_mul_13[42] + kernel_img_mul_13[43] + kernel_img_mul_13[44] + 
                kernel_img_mul_13[45] + kernel_img_mul_13[46] + kernel_img_mul_13[47] + 
                kernel_img_mul_13[48];
wire  [39:0]  kernel_img_mul_14[0:48];
assign kernel_img_mul_14[0] = layer0[14][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_14[1] = layer0[14][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_14[2] = layer0[14][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_14[3] = layer0[14][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_14[4] = layer0[14][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_14[5] = layer0[14][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_14[6] = layer0[14][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_14[7] = layer1[14][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_14[8] = layer1[14][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_14[9] = layer1[14][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_14[10] = layer1[14][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_14[11] = layer1[14][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_14[12] = layer1[14][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_14[13] = layer1[14][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_14[14] = layer2[14][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_14[15] = layer2[14][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_14[16] = layer2[14][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_14[17] = layer2[14][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_14[18] = layer2[14][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_14[19] = layer2[14][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_14[20] = layer2[14][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_14[21] = layer3[14][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_14[22] = layer3[14][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_14[23] = layer3[14][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_14[24] = layer3[14][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_14[25] = layer3[14][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_14[26] = layer3[14][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_14[27] = layer3[14][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_14[28] = layer4[14][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_14[29] = layer4[14][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_14[30] = layer4[14][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_14[31] = layer4[14][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_14[32] = layer4[14][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_14[33] = layer4[14][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_14[34] = layer4[14][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_14[35] = layer5[14][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_14[36] = layer5[14][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_14[37] = layer5[14][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_14[38] = layer5[14][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_14[39] = layer5[14][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_14[40] = layer5[14][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_14[41] = layer5[14][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_14[42] = layer6[14][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_14[43] = layer6[14][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_14[44] = layer6[14][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_14[45] = layer6[14][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_14[46] = layer6[14][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_14[47] = layer6[14][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_14[48] = layer6[14][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_14 = kernel_img_mul_14[0] + kernel_img_mul_14[1] + kernel_img_mul_14[2] + 
                kernel_img_mul_14[3] + kernel_img_mul_14[4] + kernel_img_mul_14[5] + 
                kernel_img_mul_14[6] + kernel_img_mul_14[7] + kernel_img_mul_14[8] + 
                kernel_img_mul_14[9] + kernel_img_mul_14[10] + kernel_img_mul_14[11] + 
                kernel_img_mul_14[12] + kernel_img_mul_14[13] + kernel_img_mul_14[14] + 
                kernel_img_mul_14[15] + kernel_img_mul_14[16] + kernel_img_mul_14[17] + 
                kernel_img_mul_14[18] + kernel_img_mul_14[19] + kernel_img_mul_14[20] + 
                kernel_img_mul_14[21] + kernel_img_mul_14[22] + kernel_img_mul_14[23] + 
                kernel_img_mul_14[24] + kernel_img_mul_14[25] + kernel_img_mul_14[26] + 
                kernel_img_mul_14[27] + kernel_img_mul_14[28] + kernel_img_mul_14[29] + 
                kernel_img_mul_14[30] + kernel_img_mul_14[31] + kernel_img_mul_14[32] + 
                kernel_img_mul_14[33] + kernel_img_mul_14[34] + kernel_img_mul_14[35] + 
                kernel_img_mul_14[36] + kernel_img_mul_14[37] + kernel_img_mul_14[38] + 
                kernel_img_mul_14[39] + kernel_img_mul_14[40] + kernel_img_mul_14[41] + 
                kernel_img_mul_14[42] + kernel_img_mul_14[43] + kernel_img_mul_14[44] + 
                kernel_img_mul_14[45] + kernel_img_mul_14[46] + kernel_img_mul_14[47] + 
                kernel_img_mul_14[48];
wire  [39:0]  kernel_img_mul_15[0:48];
assign kernel_img_mul_15[0] = layer0[15][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_15[1] = layer0[15][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_15[2] = layer0[15][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_15[3] = layer0[15][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_15[4] = layer0[15][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_15[5] = layer0[15][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_15[6] = layer0[15][55:48] *  G_Kernel_7x7[0][223:192];
assign kernel_img_mul_15[7] = layer1[15][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_15[8] = layer1[15][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_15[9] = layer1[15][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_15[10] = layer1[15][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_15[11] = layer1[15][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_15[12] = layer1[15][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_15[13] = layer1[15][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_15[14] = layer2[15][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_15[15] = layer2[15][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_15[16] = layer2[15][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_15[17] = layer2[15][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_15[18] = layer2[15][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_15[19] = layer2[15][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_15[20] = layer2[15][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_15[21] = layer3[15][7:0] *  G_Kernel_7x7[3][31:0];
assign kernel_img_mul_15[22] = layer3[15][15:8] *  G_Kernel_7x7[3][63:32];
assign kernel_img_mul_15[23] = layer3[15][23:16] *  G_Kernel_7x7[3][95:64];
assign kernel_img_mul_15[24] = layer3[15][31:24] *  G_Kernel_7x7[3][127:96];
assign kernel_img_mul_15[25] = layer3[15][39:32] *  G_Kernel_7x7[3][159:128];
assign kernel_img_mul_15[26] = layer3[15][47:40] *  G_Kernel_7x7[3][191:160];
assign kernel_img_mul_15[27] = layer3[15][55:48] *  G_Kernel_7x7[3][223:192];
assign kernel_img_mul_15[28] = layer4[15][7:0] *  G_Kernel_7x7[2][31:0];
assign kernel_img_mul_15[29] = layer4[15][15:8] *  G_Kernel_7x7[2][63:32];
assign kernel_img_mul_15[30] = layer4[15][23:16] *  G_Kernel_7x7[2][95:64];
assign kernel_img_mul_15[31] = layer4[15][31:24] *  G_Kernel_7x7[2][127:96];
assign kernel_img_mul_15[32] = layer4[15][39:32] *  G_Kernel_7x7[2][159:128];
assign kernel_img_mul_15[33] = layer4[15][47:40] *  G_Kernel_7x7[2][191:160];
assign kernel_img_mul_15[34] = layer4[15][55:48] *  G_Kernel_7x7[2][223:192];
assign kernel_img_mul_15[35] = layer5[15][7:0] *  G_Kernel_7x7[1][31:0];
assign kernel_img_mul_15[36] = layer5[15][15:8] *  G_Kernel_7x7[1][63:32];
assign kernel_img_mul_15[37] = layer5[15][23:16] *  G_Kernel_7x7[1][95:64];
assign kernel_img_mul_15[38] = layer5[15][31:24] *  G_Kernel_7x7[1][127:96];
assign kernel_img_mul_15[39] = layer5[15][39:32] *  G_Kernel_7x7[1][159:128];
assign kernel_img_mul_15[40] = layer5[15][47:40] *  G_Kernel_7x7[1][191:160];
assign kernel_img_mul_15[41] = layer5[15][55:48] *  G_Kernel_7x7[1][223:192];
assign kernel_img_mul_15[42] = layer6[15][7:0] *  G_Kernel_7x7[0][31:0];
assign kernel_img_mul_15[43] = layer6[15][15:8] *  G_Kernel_7x7[0][63:32];
assign kernel_img_mul_15[44] = layer6[15][23:16] *  G_Kernel_7x7[0][95:64];
assign kernel_img_mul_15[45] = layer6[15][31:24] *  G_Kernel_7x7[0][127:96];
assign kernel_img_mul_15[46] = layer6[15][39:32] *  G_Kernel_7x7[0][159:128];
assign kernel_img_mul_15[47] = layer6[15][47:40] *  G_Kernel_7x7[0][191:160];
assign kernel_img_mul_15[48] = layer6[15][55:48] *  G_Kernel_7x7[0][223:192];
wire  [39:0]  kernel_img_sum_15 = kernel_img_mul_15[0] + kernel_img_mul_15[1] + kernel_img_mul_15[2] + 
                kernel_img_mul_15[3] + kernel_img_mul_15[4] + kernel_img_mul_15[5] + 
                kernel_img_mul_15[6] + kernel_img_mul_15[7] + kernel_img_mul_15[8] + 
                kernel_img_mul_15[9] + kernel_img_mul_15[10] + kernel_img_mul_15[11] + 
                kernel_img_mul_15[12] + kernel_img_mul_15[13] + kernel_img_mul_15[14] + 
                kernel_img_mul_15[15] + kernel_img_mul_15[16] + kernel_img_mul_15[17] + 
                kernel_img_mul_15[18] + kernel_img_mul_15[19] + kernel_img_mul_15[20] + 
                kernel_img_mul_15[21] + kernel_img_mul_15[22] + kernel_img_mul_15[23] + 
                kernel_img_mul_15[24] + kernel_img_mul_15[25] + kernel_img_mul_15[26] + 
                kernel_img_mul_15[27] + kernel_img_mul_15[28] + kernel_img_mul_15[29] + 
                kernel_img_mul_15[30] + kernel_img_mul_15[31] + kernel_img_mul_15[32] + 
                kernel_img_mul_15[33] + kernel_img_mul_15[34] + kernel_img_mul_15[35] + 
                kernel_img_mul_15[36] + kernel_img_mul_15[37] + kernel_img_mul_15[38] + 
                kernel_img_mul_15[39] + kernel_img_mul_15[40] + kernel_img_mul_15[41] + 
                kernel_img_mul_15[42] + kernel_img_mul_15[43] + kernel_img_mul_15[44] + 
                kernel_img_mul_15[45] + kernel_img_mul_15[46] + kernel_img_mul_15[47] + 
                kernel_img_mul_15[48];
always @(*) begin
    blur_out[7:0] = kernel_img_sum_0[39:32];/*Q8.32 -> Q8.0*/
    blur_out[15:8] = kernel_img_sum_1[39:32];/*Q8.32 -> Q8.0*/
    blur_out[23:16] = kernel_img_sum_2[39:32];/*Q8.32 -> Q8.0*/
    blur_out[31:24] = kernel_img_sum_3[39:32];/*Q8.32 -> Q8.0*/
    blur_out[39:32] = kernel_img_sum_4[39:32];/*Q8.32 -> Q8.0*/
    blur_out[47:40] = kernel_img_sum_5[39:32];/*Q8.32 -> Q8.0*/
    blur_out[55:48] = kernel_img_sum_6[39:32];/*Q8.32 -> Q8.0*/
    blur_out[63:56] = kernel_img_sum_7[39:32];/*Q8.32 -> Q8.0*/
    blur_out[71:64] = kernel_img_sum_8[39:32];/*Q8.32 -> Q8.0*/
    blur_out[79:72] = kernel_img_sum_9[39:32];/*Q8.32 -> Q8.0*/
    blur_out[87:80] = kernel_img_sum_10[39:32];/*Q8.32 -> Q8.0*/
    blur_out[95:88] = kernel_img_sum_11[39:32];/*Q8.32 -> Q8.0*/
    blur_out[103:96] = kernel_img_sum_12[39:32];/*Q8.32 -> Q8.0*/
    blur_out[111:104] = kernel_img_sum_13[39:32];/*Q8.32 -> Q8.0*/
    blur_out[119:112] = kernel_img_sum_14[39:32];/*Q8.32 -> Q8.0*/
    blur_out[127:120] = kernel_img_sum_15[39:32];/*Q8.32 -> Q8.0*/
end


endmodule